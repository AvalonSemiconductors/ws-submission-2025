* NGSPICE file created from flattened.ext - technology: gf180mcuD

.subckt opamp_chonky_spice PLUS MINUS ADJ OUT VDD VSS
X0 OUT.t81 a_31459_5010.t2 VSS.t48 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X1 VDD.t49 ADJ.t2 OUT.t17 VDD.t1 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X2 OUT.t37 ADJ.t3 VDD.t48 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X3 OUT.t39 ADJ.t4 VDD.t47 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X4 OUT.t83 ADJ.t5 VDD.t46 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X5 VDD.t45 ADJ.t6 OUT.t11 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X6 OUT.t80 a_31459_5010.t3 VSS.t47 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X7 a_31459_5010.t1 a_30739_5010.t3 VSS.t1 VSS.t0 nfet_05v0 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=0.6u
X8 VSS.t46 a_31459_5010.t4 OUT.t79 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X9 OUT.t78 a_31459_5010.t5 VSS.t40 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X10 VDD.t44 ADJ.t7 OUT.t5 VDD.t13 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X11 VSS.t43 a_31459_5010.t6 OUT.t77 VSS.t4 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X12 VSS.t45 a_31459_5010.t7 OUT.t76 VSS.t11 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X13 a_30873_8186.t2 MINUS.t0 a_30739_5010.t0 VDD.t0 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X14 OUT.t29 ADJ.t8 VDD.t43 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X15 OUT.t75 a_31459_5010.t8 VSS.t44 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X16 VSS.t42 a_31459_5010.t9 OUT.t74 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X17 VSS.t41 a_31459_5010.t10 OUT.t73 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X18 OUT.t72 a_31459_5010.t11 VSS.t39 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X19 VSS.t38 a_31459_5010.t12 OUT.t71 VSS.t6 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X20 VDD.t42 ADJ.t9 OUT.t23 VDD.t13 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X21 VDD.t41 ADJ.t10 OUT.t10 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X22 OUT.t70 a_31459_5010.t13 VSS.t37 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X23 VSS.t36 a_31459_5010.t14 OUT.t69 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X24 VSS.t35 a_31459_5010.t15 OUT.t68 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X25 VSS.t34 a_31459_5010.t16 OUT.t67 VSS.t11 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X26 OUT.t66 a_31459_5010.t17 VSS.t30 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X27 VDD.t40 ADJ.t11 OUT.t2 VDD.t1 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X28 OUT.t65 a_31459_5010.t18 VSS.t33 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X29 VSS.t32 a_31459_5010.t19 OUT.t64 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X30 VDD.t39 ADJ.t12 OUT.t35 VDD.t7 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X31 VSS.t29 a_31459_5010.t20 OUT.t63 VSS.t6 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X32 VDD.t38 ADJ.t13 OUT.t16 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X33 OUT.t28 ADJ.t14 VDD.t37 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X34 VDD.t36 ADJ.t15 OUT.t22 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X35 OUT.t9 ADJ.t16 VDD.t35 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X36 VSS.t31 a_31459_5010.t21 OUT.t62 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X37 VSS.t28 a_31459_5010.t22 OUT.t61 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X38 VDD.t34 ADJ.t17 OUT.t34 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X39 VDD.t33 ADJ.t18 OUT.t15 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X40 VDD.t32 ADJ.t19 OUT.t36 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X41 a_31459_5010.t0 PLUS.t0 a_30873_8186.t1 VDD.t50 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X42 OUT.t38 ADJ.t20 VDD.t31 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X43 OUT.t82 ADJ.t21 VDD.t30 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X44 VSS.t27 a_31459_5010.t23 OUT.t60 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X45 OUT.t59 a_31459_5010.t24 VSS.t26 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X46 VDD.t29 ADJ.t22 OUT.t8 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X47 VDD.t8 ADJ.t23 OUT.t4 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X48 OUT.t27 ADJ.t24 VDD.t28 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X49 OUT.t21 ADJ.t25 VDD.t27 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X50 OUT.t7 ADJ.t26 VDD.t24 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X51 VSS.t25 a_31459_5010.t25 OUT.t58 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X52 VSS.t24 a_31459_5010.t26 OUT.t57 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X53 OUT.t1 ADJ.t27 VDD.t26 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X54 VSS.t20 a_31459_5010.t27 OUT.t56 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X55 OUT.t55 a_31459_5010.t28 VSS.t23 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X56 VDD.t25 ADJ.t28 OUT.t33 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X57 OUT.t54 a_31459_5010.t29 VSS.t22 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X58 VSS.t21 a_31459_5010.t30 OUT.t53 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X59 OUT.t52 a_31459_5010.t31 VSS.t19 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X60 VDD.t23 ADJ.t29 a_30873_8186.t0 VDD.t22 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X61 OUT.t26 ADJ.t30 VDD.t21 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X62 VDD.t20 ADJ.t31 OUT.t20 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X63 VSS.t18 a_31459_5010.t32 OUT.t51 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X64 VSS.t3 a_30739_5010.t1 a_30739_5010.t2 VSS.t2 nfet_05v0 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=0.6u
X65 VSS.t17 a_31459_5010.t33 OUT.t50 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X66 VDD.t19 ADJ.t32 OUT.t6 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X67 OUT.t49 a_31459_5010.t34 VSS.t16 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X68 OUT.t48 a_31459_5010.t35 VSS.t15 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X69 VSS.t14 a_31459_5010.t36 OUT.t47 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X70 VSS.t13 a_31459_5010.t37 OUT.t46 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X71 OUT.t32 ADJ.t33 VDD.t18 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X72 OUT.t45 a_31459_5010.t38 VSS.t9 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X73 OUT.t14 ADJ.t34 VDD.t17 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X74 VDD.t16 ADJ.t35 OUT.t31 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X75 VDD.t15 ADJ.t36 OUT.t13 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X76 OUT.t3 ADJ.t37 VDD.t14 VDD.t13 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X77 OUT.t44 a_31459_5010.t39 VSS.t12 VSS.t11 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X78 OUT.t25 ADJ.t38 VDD.t12 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X79 VDD.t11 ADJ.t39 OUT.t19 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X80 VDD.t6 ADJ.t40 OUT.t0 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X81 OUT.t43 a_31459_5010.t40 VSS.t10 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X82 VDD.t10 ADJ.t41 OUT.t30 VDD.t7 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X83 VDD.t9 ADJ.t42 OUT.t12 VDD.t7 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X84 VSS.t8 a_31459_5010.t41 OUT.t42 VSS.t4 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X85 OUT.t41 a_31459_5010.t42 VSS.t7 VSS.t6 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X86 VDD.t5 ADJ.t0 ADJ.t1 VDD.t4 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X87 OUT.t24 ADJ.t43 VDD.t3 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X88 VDD.t2 ADJ.t44 OUT.t18 VDD.t1 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X89 VSS.t5 a_31459_5010.t43 OUT.t40 VSS.t4 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
R0 a_31459_5010.n11 a_31459_5010.t6 620.048
R1 a_31459_5010.n13 a_31459_5010.t16 620.048
R2 a_31459_5010.t32 a_31459_5010.n2 620.048
R3 a_31459_5010.t27 a_31459_5010.n67 620.048
R4 a_31459_5010.n55 a_31459_5010.t9 620.048
R5 a_31459_5010.n36 a_31459_5010.t7 620.048
R6 a_31459_5010.t41 a_31459_5010.n33 620.048
R7 a_31459_5010.t43 a_31459_5010.n48 620.048
R8 a_31459_5010.t39 a_31459_5010.n36 619.74
R9 a_31459_5010.n33 a_31459_5010.t35 619.74
R10 a_31459_5010.t33 a_31459_5010.n29 619.74
R11 a_31459_5010.t26 a_31459_5010.n24 619.74
R12 a_31459_5010.n44 a_31459_5010.t28 619.74
R13 a_31459_5010.n62 a_31459_5010.t24 619.74
R14 a_31459_5010.t14 a_31459_5010.n56 619.74
R15 a_31459_5010.t4 a_31459_5010.n25 619.74
R16 a_31459_5010.n67 a_31459_5010.t2 619.74
R17 a_31459_5010.t11 a_31459_5010.n2 619.74
R18 a_31459_5010.n66 a_31459_5010.t10 619.74
R19 a_31459_5010.n77 a_31459_5010.t21 619.74
R20 a_31459_5010.n64 a_31459_5010.t3 619.74
R21 a_31459_5010.n78 a_31459_5010.t13 619.74
R22 a_31459_5010.t34 a_31459_5010.n13 619.74
R23 a_31459_5010.t29 a_31459_5010.n11 619.74
R24 a_31459_5010.t25 a_31459_5010.n1 619.74
R25 a_31459_5010.t23 a_31459_5010.n7 619.74
R26 a_31459_5010.n48 a_31459_5010.t40 619.74
R27 a_31459_5010.n55 a_31459_5010.t5 619.74
R28 a_31459_5010.n37 a_31459_5010.t42 614.254
R29 a_31459_5010.n37 a_31459_5010.t39 614.254
R30 a_31459_5010.n32 a_31459_5010.t42 614.254
R31 a_31459_5010.t35 a_31459_5010.n32 614.254
R32 a_31459_5010.n40 a_31459_5010.t36 614.254
R33 a_31459_5010.n40 a_31459_5010.t33 614.254
R34 a_31459_5010.t36 a_31459_5010.n39 614.254
R35 a_31459_5010.n39 a_31459_5010.t26 614.254
R36 a_31459_5010.n43 a_31459_5010.t31 614.254
R37 a_31459_5010.t28 a_31459_5010.n43 614.254
R38 a_31459_5010.n61 a_31459_5010.t31 614.254
R39 a_31459_5010.t24 a_31459_5010.n61 614.254
R40 a_31459_5010.t19 a_31459_5010.n57 614.254
R41 a_31459_5010.n57 a_31459_5010.t14 614.254
R42 a_31459_5010.n58 a_31459_5010.t19 614.254
R43 a_31459_5010.n58 a_31459_5010.t4 614.254
R44 a_31459_5010.n72 a_31459_5010.t2 614.254
R45 a_31459_5010.t17 a_31459_5010.n72 614.254
R46 a_31459_5010.n73 a_31459_5010.t17 614.254
R47 a_31459_5010.n73 a_31459_5010.t11 614.254
R48 a_31459_5010.t10 a_31459_5010.n65 614.254
R49 a_31459_5010.n65 a_31459_5010.t22 614.254
R50 a_31459_5010.n76 a_31459_5010.t22 614.254
R51 a_31459_5010.t21 a_31459_5010.n76 614.254
R52 a_31459_5010.t3 a_31459_5010.n22 614.254
R53 a_31459_5010.n22 a_31459_5010.t18 614.254
R54 a_31459_5010.t18 a_31459_5010.n21 614.254
R55 a_31459_5010.n21 a_31459_5010.t13 614.254
R56 a_31459_5010.n14 a_31459_5010.t38 614.254
R57 a_31459_5010.n14 a_31459_5010.t34 614.254
R58 a_31459_5010.n12 a_31459_5010.t29 614.254
R59 a_31459_5010.t38 a_31459_5010.n12 614.254
R60 a_31459_5010.t30 a_31459_5010.n17 614.254
R61 a_31459_5010.n17 a_31459_5010.t25 614.254
R62 a_31459_5010.n18 a_31459_5010.t23 614.254
R63 a_31459_5010.n18 a_31459_5010.t30 614.254
R64 a_31459_5010.t6 a_31459_5010.n10 614.254
R65 a_31459_5010.n10 a_31459_5010.t20 614.254
R66 a_31459_5010.t20 a_31459_5010.n9 614.254
R67 a_31459_5010.t16 a_31459_5010.n9 614.254
R68 a_31459_5010.t37 a_31459_5010.n68 614.254
R69 a_31459_5010.n68 a_31459_5010.t32 614.254
R70 a_31459_5010.n69 a_31459_5010.t27 614.254
R71 a_31459_5010.n69 a_31459_5010.t37 614.254
R72 a_31459_5010.t40 a_31459_5010.n47 614.254
R73 a_31459_5010.n47 a_31459_5010.t8 614.254
R74 a_31459_5010.n54 a_31459_5010.t8 614.254
R75 a_31459_5010.t5 a_31459_5010.n54 614.254
R76 a_31459_5010.n51 a_31459_5010.t9 614.254
R77 a_31459_5010.n35 a_31459_5010.t12 614.254
R78 a_31459_5010.t7 a_31459_5010.n35 614.254
R79 a_31459_5010.t12 a_31459_5010.n34 614.254
R80 a_31459_5010.n34 a_31459_5010.t41 614.254
R81 a_31459_5010.n50 a_31459_5010.t43 614.254
R82 a_31459_5010.t15 a_31459_5010.n50 614.254
R83 a_31459_5010.n51 a_31459_5010.t15 614.254
R84 a_31459_5010.n63 a_31459_5010.n23 15.7039
R85 a_31459_5010.n46 a_31459_5010.n45 15.3876
R86 a_31459_5010.n46 a_31459_5010.n23 14.6668
R87 a_31459_5010.n15 a_31459_5010.n9 5.13335
R88 a_31459_5010.n10 a_31459_5010.n8 5.13335
R89 a_31459_5010.n35 a_31459_5010.n30 5.02611
R90 a_31459_5010.n54 a_31459_5010.n53 5.02611
R91 a_31459_5010.n34 a_31459_5010.n6 5.02611
R92 a_31459_5010.n38 a_31459_5010.n37 5.02611
R93 a_31459_5010.n32 a_31459_5010.n31 5.02611
R94 a_31459_5010.n41 a_31459_5010.n40 5.02611
R95 a_31459_5010.n39 a_31459_5010.n26 5.02611
R96 a_31459_5010.n43 a_31459_5010.n42 5.02611
R97 a_31459_5010.n61 a_31459_5010.n60 5.02611
R98 a_31459_5010.n57 a_31459_5010.n28 5.02611
R99 a_31459_5010.n59 a_31459_5010.n58 5.02611
R100 a_31459_5010.n50 a_31459_5010.n49 5.02611
R101 a_31459_5010.n70 a_31459_5010.n69 5.02611
R102 a_31459_5010.n68 a_31459_5010.n4 5.02611
R103 a_31459_5010.n74 a_31459_5010.n73 5.02611
R104 a_31459_5010.n72 a_31459_5010.n71 5.02611
R105 a_31459_5010.n76 a_31459_5010.n75 5.02611
R106 a_31459_5010.n65 a_31459_5010.n5 5.02611
R107 a_31459_5010.n21 a_31459_5010.n3 5.02611
R108 a_31459_5010.n22 a_31459_5010.n20 5.02611
R109 a_31459_5010.n12 a_31459_5010.n8 5.02611
R110 a_31459_5010.n15 a_31459_5010.n14 5.02611
R111 a_31459_5010.n19 a_31459_5010.n18 5.02611
R112 a_31459_5010.n17 a_31459_5010.n16 5.02611
R113 a_31459_5010.n47 a_31459_5010.n27 5.02611
R114 a_31459_5010.n52 a_31459_5010.n51 5.02611
R115 a_31459_5010.n64 a_31459_5010.n63 2.8286
R116 a_31459_5010.n79 a_31459_5010.n0 1.12638
R117 a_31459_5010.n0 a_31459_5010.t1 1.04563
R118 a_31459_5010.t0 a_31459_5010.n79 0.96115
R119 a_31459_5010.n70 a_31459_5010.n6 0.437096
R120 a_31459_5010.n30 a_31459_5010.n4 0.437096
R121 a_31459_5010.n63 a_31459_5010.n62 0.321929
R122 a_31459_5010.n45 a_31459_5010.n44 0.321929
R123 a_31459_5010.n79 a_31459_5010.n78 0.321929
R124 a_31459_5010.n64 a_31459_5010.n7 0.308818
R125 a_31459_5010.n11 a_31459_5010.n7 0.308818
R126 a_31459_5010.n13 a_31459_5010.n1 0.308818
R127 a_31459_5010.n78 a_31459_5010.n1 0.308818
R128 a_31459_5010.n78 a_31459_5010.n77 0.308818
R129 a_31459_5010.n77 a_31459_5010.n2 0.308818
R130 a_31459_5010.n67 a_31459_5010.n66 0.308818
R131 a_31459_5010.n66 a_31459_5010.n64 0.308818
R132 a_31459_5010.n56 a_31459_5010.n55 0.308818
R133 a_31459_5010.n56 a_31459_5010.n44 0.308818
R134 a_31459_5010.n44 a_31459_5010.n29 0.308818
R135 a_31459_5010.n36 a_31459_5010.n29 0.308818
R136 a_31459_5010.n33 a_31459_5010.n24 0.308818
R137 a_31459_5010.n62 a_31459_5010.n24 0.308818
R138 a_31459_5010.n62 a_31459_5010.n25 0.308818
R139 a_31459_5010.n48 a_31459_5010.n25 0.308818
R140 a_31459_5010.n45 a_31459_5010.n0 0.157817
R141 a_31459_5010.n49 a_31459_5010.n23 0.130713
R142 a_31459_5010.n52 a_31459_5010.n46 0.130713
R143 a_31459_5010.n19 a_31459_5010.n8 0.107734
R144 a_31459_5010.n20 a_31459_5010.n19 0.107734
R145 a_31459_5010.n20 a_31459_5010.n5 0.107734
R146 a_31459_5010.n71 a_31459_5010.n5 0.107734
R147 a_31459_5010.n71 a_31459_5010.n70 0.107734
R148 a_31459_5010.n31 a_31459_5010.n6 0.107734
R149 a_31459_5010.n31 a_31459_5010.n26 0.107734
R150 a_31459_5010.n60 a_31459_5010.n26 0.107734
R151 a_31459_5010.n60 a_31459_5010.n59 0.107734
R152 a_31459_5010.n59 a_31459_5010.n27 0.107734
R153 a_31459_5010.n49 a_31459_5010.n27 0.107734
R154 a_31459_5010.n16 a_31459_5010.n15 0.107734
R155 a_31459_5010.n16 a_31459_5010.n3 0.107734
R156 a_31459_5010.n75 a_31459_5010.n3 0.107734
R157 a_31459_5010.n75 a_31459_5010.n74 0.107734
R158 a_31459_5010.n74 a_31459_5010.n4 0.107734
R159 a_31459_5010.n38 a_31459_5010.n30 0.107734
R160 a_31459_5010.n41 a_31459_5010.n38 0.107734
R161 a_31459_5010.n42 a_31459_5010.n41 0.107734
R162 a_31459_5010.n42 a_31459_5010.n28 0.107734
R163 a_31459_5010.n53 a_31459_5010.n28 0.107734
R164 a_31459_5010.n53 a_31459_5010.n52 0.107734
R165 VSS.t6 VSS.t4 14065
R166 VSS.t6 VSS.t11 14065
R167 VSS.n72 VSS.t11 7182.67
R168 VSS.t2 VSS.n73 328.293
R169 VSS.n74 VSS.t0 328.077
R170 VSS.n74 VSS.t2 328.077
R171 VSS.t0 VSS.n72 327.49
R172 VSS.n71 VSS.n4 161.779
R173 VSS.n71 VSS.n5 161.779
R174 VSS.n73 VSS.n4 161.779
R175 VSS.n73 VSS.n5 161.779
R176 VSS.n75 VSS.n4 112.001
R177 VSS.n75 VSS.n5 112.001
R178 VSS.n29 VSS.n27 34.1162
R179 VSS.n43 VSS.n41 34.1096
R180 VSS.n35 VSS.n33 34.1096
R181 VSS.n50 VSS.n48 34.1085
R182 VSS.n65 VSS.n63 34.1074
R183 VSS.n57 VSS.n55 34.1063
R184 VSS.n30 VSS.n25 25.6892
R185 VSS.n51 VSS.n22 25.6794
R186 VSS.n61 VSS.n9 25.6774
R187 VSS.n58 VSS.n53 25.6774
R188 VSS.n39 VSS.n24 25.6755
R189 VSS.n36 VSS.n31 25.6559
R190 VSS.n14 VSS.n13 7.83243
R191 VSS.n14 VSS.n0 6.85872
R192 VSS.n36 VSS.n35 6.58153
R193 VSS.n41 VSS.n39 6.56196
R194 VSS.n63 VSS.n61 6.56001
R195 VSS.n58 VSS.n57 6.56001
R196 VSS.n51 VSS.n50 6.55805
R197 VSS.n30 VSS.n29 6.54827
R198 VSS.n17 VSS.n7 5.95109
R199 VSS.n12 VSS.n10 4.41109
R200 VSS.n78 VSS.n1 4.3205
R201 VSS.n68 VSS.n67 4.01281
R202 VSS.n13 VSS.n12 4.0018
R203 VSS.n3 VSS.n2 3.28159
R204 VSS.n19 VSS.n16 3.08674
R205 VSS.n77 VSS.n2 2.79681
R206 VSS.n20 VSS.n11 2.28848
R207 VSS.n69 VSS.n3 1.62406
R208 VSS.n17 VSS.n10 1.5405
R209 VSS.n13 VSS.n11 1.52562
R210 VSS.n68 VSS.n6 1.52318
R211 VSS.n78 VSS.n77 1.01317
R212 VSS.n20 VSS.n19 0.798754
R213 VSS.n76 VSS.n3 0.596161
R214 VSS.n77 VSS.n76 0.596161
R215 VSS.n76 VSS.t3 0.4643
R216 VSS.n76 VSS.t1 0.4643
R217 VSS.n1 VSS.n0 0.459071
R218 VSS.n70 VSS.n69 0.447421
R219 VSS.n71 VSS.n70 0.218565
R220 VSS.n76 VSS.n75 0.217167
R221 VSS.n75 VSS.n74 0.217167
R222 VSS.n73 VSS.n2 0.217167
R223 VSS.n72 VSS.n71 0.217167
R224 VSS.n27 VSS.n23 0.0597094
R225 VSS.n60 VSS.n10 0.0547889
R226 VSS.n37 VSS.n30 0.0547889
R227 VSS.n37 VSS.n36 0.0505
R228 VSS.n39 VSS.n38 0.0505
R229 VSS.n52 VSS.n51 0.0505
R230 VSS.n59 VSS.n58 0.0505
R231 VSS.n61 VSS.n60 0.0505
R232 VSS.n7 VSS.t34 0.0464575
R233 VSS.n17 VSS.t29 0.0464575
R234 VSS.n12 VSS.t43 0.0464575
R235 VSS.n16 VSS.t45 0.0464575
R236 VSS.n19 VSS.t38 0.0464575
R237 VSS.n11 VSS.t8 0.0464575
R238 VSS.n44 VSS.n43 0.043625
R239 VSS.n33 VSS.n23 0.043625
R240 VSS.n48 VSS.n46 0.0422188
R241 VSS.n66 VSS.n65 0.0408125
R242 VSS.n55 VSS.n8 0.039529
R243 VSS.n63 VSS.n62 0.0300775
R244 VSS.n65 VSS.n64 0.0300775
R245 VSS.n57 VSS.n56 0.0300775
R246 VSS.n55 VSS.n54 0.0300775
R247 VSS.n50 VSS.n49 0.0300775
R248 VSS.n48 VSS.n47 0.0300775
R249 VSS.n41 VSS.n40 0.0300775
R250 VSS.n43 VSS.n42 0.0300775
R251 VSS.n35 VSS.n34 0.0300775
R252 VSS.n33 VSS.n32 0.0300775
R253 VSS.n27 VSS.n26 0.0300775
R254 VSS.n29 VSS.n28 0.0300775
R255 VSS.n67 VSS.n66 0.0259594
R256 VSS.n69 VSS.n68 0.0238731
R257 VSS.n19 VSS.n15 0.017599
R258 VSS.n15 VSS.n14 0.017599
R259 VSS.n18 VSS.n17 0.017099
R260 VSS.n19 VSS.n18 0.017099
R261 VSS.n28 VSS.t44 0.01688
R262 VSS.n28 VSS.t35 0.01688
R263 VSS.n26 VSS.t40 0.01688
R264 VSS.n26 VSS.t42 0.01688
R265 VSS.n64 VSS.t16 0.01688
R266 VSS.n64 VSS.t25 0.01688
R267 VSS.n62 VSS.t9 0.01688
R268 VSS.n62 VSS.t21 0.01688
R269 VSS.n9 VSS.t22 0.01688
R270 VSS.n9 VSS.t27 0.01688
R271 VSS.n54 VSS.t37 0.01688
R272 VSS.n54 VSS.t31 0.01688
R273 VSS.n56 VSS.t33 0.01688
R274 VSS.n56 VSS.t28 0.01688
R275 VSS.n53 VSS.t47 0.01688
R276 VSS.n53 VSS.t41 0.01688
R277 VSS.n47 VSS.t39 0.01688
R278 VSS.n47 VSS.t18 0.01688
R279 VSS.n49 VSS.t30 0.01688
R280 VSS.n49 VSS.t13 0.01688
R281 VSS.n22 VSS.t48 0.01688
R282 VSS.n22 VSS.t20 0.01688
R283 VSS.n42 VSS.t12 0.01688
R284 VSS.n42 VSS.t17 0.01688
R285 VSS.n40 VSS.t7 0.01688
R286 VSS.n40 VSS.t14 0.01688
R287 VSS.n24 VSS.t15 0.01688
R288 VSS.n24 VSS.t24 0.01688
R289 VSS.n32 VSS.t23 0.01688
R290 VSS.n32 VSS.t36 0.01688
R291 VSS.n34 VSS.t19 0.01688
R292 VSS.n34 VSS.t32 0.01688
R293 VSS.n31 VSS.t26 0.01688
R294 VSS.n31 VSS.t46 0.01688
R295 VSS.n25 VSS.t10 0.01688
R296 VSS.n25 VSS.t5 0.01688
R297 VSS VSS.n78 0.016025
R298 VSS.n21 VSS.n20 0.00896236
R299 VSS.n70 VSS.n1 0.0086575
R300 VSS.n38 VSS.n21 0.00751474
R301 VSS.n52 VSS.n21 0.00738071
R302 VSS.n67 VSS.n7 0.00491176
R303 VSS.n60 VSS.n59 0.00478891
R304 VSS.n59 VSS.n52 0.00478891
R305 VSS.n38 VSS.n37 0.00478891
R306 VSS.n45 VSS.n6 0.00440625
R307 VSS VSS.n0 0.003875
R308 VSS.n45 VSS.n44 0.00371783
R309 VSS.n46 VSS.n45 0.00341997
R310 VSS.n16 VSS.n6 0.00294068
R311 VSS.n66 VSS.n8 0.00252186
R312 VSS.n46 VSS.n8 0.00252186
R313 VSS.n44 VSS.n23 0.00252186
R314 VSS.t6 VSS.n15 0.00150002
R315 VSS.n18 VSS.t6 0.00100002
R316 OUT.n87 OUT.n85 34.1284
R317 OUT.n82 OUT.n80 34.1273
R318 OUT.n75 OUT.n73 34.1273
R319 OUT.n27 OUT.n25 34.1267
R320 OUT.n18 OUT.n8 34.1262
R321 OUT.n99 OUT.n97 34.1245
R322 OUT.n67 OUT.n66 34.1245
R323 OUT.n38 OUT.n37 34.1225
R324 OUT.n55 OUT.n53 34.1225
R325 OUT.n94 OUT.n93 34.1206
R326 OUT.n62 OUT.n60 34.1206
R327 OUT.n14 OUT.n13 34.1186
R328 OUT.n51 OUT.n50 34.1167
R329 OUT.n44 OUT.n42 34.1147
R330 OUT.n22 OUT.n2 34.1147
R331 OUT.n106 OUT.n105 34.1089
R332 OUT.n23 OUT.t74 26.7643
R333 OUT.n104 OUT.t31 26.7629
R334 OUT.n35 OUT.n33 26.7616
R335 OUT.n57 OUT.n56 26.7616
R336 OUT.n20 OUT.n19 26.7596
R337 OUT.n64 OUT.n63 26.7596
R338 OUT.n92 OUT.t18 26.757
R339 OUT.n71 OUT.n16 26.7538
R340 OUT.n29 OUT.n28 26.7538
R341 OUT.n48 OUT.n40 26.7447
R342 OUT.n11 OUT.n10 26.7408
R343 OUT.n46 OUT.n45 26.7388
R344 OUT.n78 OUT.n77 26.7388
R345 OUT.n101 OUT.n100 26.7369
R346 OUT.n89 OUT.n88 26.7349
R347 OUT.n68 OUT.t51 26.6707
R348 OUT.n89 OUT.n87 7.71659
R349 OUT.n101 OUT.n99 7.71464
R350 OUT.n46 OUT.n44 7.71268
R351 OUT.n80 OUT.n78 7.71268
R352 OUT.n93 OUT.n92 7.71268
R353 OUT.n13 OUT.n11 7.71072
R354 OUT.n23 OUT.n22 7.70877
R355 OUT.n50 OUT.n48 7.70681
R356 OUT.n105 OUT.n104 7.70681
R357 OUT.n73 OUT.n71 7.7029
R358 OUT.n29 OUT.n27 7.7029
R359 OUT.n20 OUT.n18 7.69703
R360 OUT.n64 OUT.n62 7.69703
R361 OUT.n37 OUT.n35 7.69507
R362 OUT.n57 OUT.n55 7.69507
R363 OUT.n68 OUT.n67 7.59954
R364 OUT OUT.n0 1.92133
R365 OUT OUT.n107 0.109695
R366 OUT.n47 OUT.n46 0.0547894
R367 OUT.n30 OUT.n23 0.0547894
R368 OUT.n106 OUT.t20 0.0543631
R369 OUT.n2 OUT.t40 0.0534887
R370 OUT.n30 OUT.n29 0.0505
R371 OUT.n58 OUT.n57 0.0505
R372 OUT.n65 OUT.n64 0.0505
R373 OUT.n69 OUT.n68 0.0505
R374 OUT.n71 OUT.n70 0.0505
R375 OUT.n21 OUT.n20 0.0505
R376 OUT.n35 OUT.n34 0.0505
R377 OUT.n92 OUT.n91 0.0505
R378 OUT.n90 OUT.n89 0.0505
R379 OUT.n78 OUT.n4 0.0505
R380 OUT.n102 OUT.n101 0.0505
R381 OUT.n104 OUT.n103 0.0505
R382 OUT.n11 OUT.n3 0.0505
R383 OUT.n48 OUT.n47 0.0505
R384 OUT.n22 OUT.t68 0.0464575
R385 OUT.n67 OUT.t46 0.0464575
R386 OUT.n66 OUT.t56 0.0464575
R387 OUT.n94 OUT.t13 0.0459256
R388 OUT.n105 OUT.t19 0.0431131
R389 OUT.n93 OUT.t11 0.0431131
R390 OUT.n85 OUT.n83 0.0339259
R391 OUT.n60 OUT.n59 0.03289
R392 OUT.n42 OUT.n41 0.0319444
R393 OUT.n38 OUT.n32 0.0314837
R394 OUT.n53 OUT.n31 0.0314837
R395 OUT.n83 OUT.n82 0.0310915
R396 OUT.n76 OUT.n75 0.0310915
R397 OUT.n51 OUT.n39 0.0305381
R398 OUT.n37 OUT.n36 0.0300775
R399 OUT.n8 OUT.n7 0.0300775
R400 OUT.n18 OUT.n17 0.0300775
R401 OUT.n75 OUT.n74 0.0300775
R402 OUT.n73 OUT.n72 0.0300775
R403 OUT.n62 OUT.n61 0.0300775
R404 OUT.n55 OUT.n54 0.0300775
R405 OUT.n25 OUT.n24 0.0300775
R406 OUT.n27 OUT.n26 0.0300775
R407 OUT.n25 OUT.n6 0.0296852
R408 OUT.n14 OUT.n9 0.0291319
R409 OUT.n96 OUT.n8 0.028279
R410 OUT.n44 OUT.n43 0.0249131
R411 OUT.n50 OUT.n49 0.0249131
R412 OUT.n13 OUT.n12 0.0249131
R413 OUT.n97 OUT.n5 0.0249131
R414 OUT.n99 OUT.n98 0.0249131
R415 OUT.n82 OUT.n81 0.0249131
R416 OUT.n80 OUT.n79 0.0249131
R417 OUT.n85 OUT.n84 0.0249131
R418 OUT.n87 OUT.n86 0.0249131
R419 OUT.n107 OUT.n2 0.0240602
R420 OUT.n53 OUT.n52 0.0240602
R421 OUT.n60 OUT.n1 0.0240602
R422 OUT.n66 OUT.n15 0.0240602
R423 OUT.n52 OUT.n38 0.0240602
R424 OUT.n95 OUT.n94 0.0240602
R425 OUT.n97 OUT.n96 0.0240602
R426 OUT.n107 OUT.n106 0.0240602
R427 OUT.n15 OUT.n14 0.0240602
R428 OUT.n52 OUT.n51 0.0240602
R429 OUT.n42 OUT.n1 0.0240602
R430 OUT.n45 OUT.t17 0.0187
R431 OUT.n45 OUT.t25 0.0187
R432 OUT.n43 OUT.t30 0.0187
R433 OUT.n43 OUT.t32 0.0187
R434 OUT.n41 OUT.t23 0.0187
R435 OUT.n41 OUT.t37 0.0187
R436 OUT.n40 OUT.t8 0.0187
R437 OUT.n40 OUT.t1 0.0187
R438 OUT.n49 OUT.t15 0.0187
R439 OUT.n49 OUT.t7 0.0187
R440 OUT.n39 OUT.t33 0.0187
R441 OUT.n39 OUT.t26 0.0187
R442 OUT.n10 OUT.t36 0.0187
R443 OUT.n10 OUT.t24 0.0187
R444 OUT.n12 OUT.t4 0.0187
R445 OUT.n12 OUT.t39 0.0187
R446 OUT.n9 OUT.t16 0.0187
R447 OUT.n9 OUT.t14 0.0187
R448 OUT.n100 OUT.t2 0.0187
R449 OUT.n100 OUT.t83 0.0187
R450 OUT.n98 OUT.t35 0.0187
R451 OUT.n98 OUT.t29 0.0187
R452 OUT.n5 OUT.t5 0.0187
R453 OUT.n5 OUT.t3 0.0187
R454 OUT.n77 OUT.t0 0.0187
R455 OUT.n77 OUT.t38 0.0187
R456 OUT.n79 OUT.t12 0.0187
R457 OUT.n79 OUT.t27 0.0187
R458 OUT.n81 OUT.t6 0.0187
R459 OUT.n81 OUT.t28 0.0187
R460 OUT.n88 OUT.t22 0.0187
R461 OUT.n88 OUT.t82 0.0187
R462 OUT.n86 OUT.t34 0.0187
R463 OUT.n86 OUT.t21 0.0187
R464 OUT.n84 OUT.t10 0.0187
R465 OUT.n84 OUT.t9 0.0187
R466 OUT.n33 OUT.t67 0.01688
R467 OUT.n33 OUT.t49 0.01688
R468 OUT.n36 OUT.t63 0.01688
R469 OUT.n36 OUT.t45 0.01688
R470 OUT.n32 OUT.t77 0.01688
R471 OUT.n32 OUT.t54 0.01688
R472 OUT.n19 OUT.t58 0.01688
R473 OUT.n19 OUT.t70 0.01688
R474 OUT.n17 OUT.t53 0.01688
R475 OUT.n17 OUT.t65 0.01688
R476 OUT.n7 OUT.t60 0.01688
R477 OUT.n7 OUT.t80 0.01688
R478 OUT.n16 OUT.t62 0.01688
R479 OUT.n16 OUT.t72 0.01688
R480 OUT.n72 OUT.t61 0.01688
R481 OUT.n72 OUT.t66 0.01688
R482 OUT.n74 OUT.t73 0.01688
R483 OUT.n74 OUT.t81 0.01688
R484 OUT.n63 OUT.t76 0.01688
R485 OUT.n63 OUT.t44 0.01688
R486 OUT.n61 OUT.t71 0.01688
R487 OUT.n61 OUT.t41 0.01688
R488 OUT.n59 OUT.t42 0.01688
R489 OUT.n59 OUT.t48 0.01688
R490 OUT.n56 OUT.t50 0.01688
R491 OUT.n56 OUT.t55 0.01688
R492 OUT.n54 OUT.t47 0.01688
R493 OUT.n54 OUT.t52 0.01688
R494 OUT.n31 OUT.t57 0.01688
R495 OUT.n31 OUT.t59 0.01688
R496 OUT.n28 OUT.t69 0.01688
R497 OUT.n28 OUT.t78 0.01688
R498 OUT.n26 OUT.t64 0.01688
R499 OUT.n26 OUT.t75 0.01688
R500 OUT.n24 OUT.t79 0.01688
R501 OUT.n24 OUT.t43 0.01688
R502 OUT.n69 OUT.n65 0.00924149
R503 OUT.n103 OUT.n102 0.00923191
R504 OUT.n34 OUT.n0 0.00635957
R505 OUT.n47 OUT.n3 0.00478936
R506 OUT.n103 OUT.n3 0.00478936
R507 OUT.n102 OUT.n4 0.00478936
R508 OUT.n90 OUT.n4 0.00478936
R509 OUT.n91 OUT.n90 0.00478936
R510 OUT.n34 OUT.n21 0.00478936
R511 OUT.n70 OUT.n21 0.00478936
R512 OUT.n65 OUT.n58 0.00478936
R513 OUT.n58 OUT.n30 0.00478936
R514 OUT.n70 OUT.n69 0.00477979
R515 OUT.n91 OUT.n0 0.00293191
R516 OUT.n83 OUT.n76 0.000532943
R517 OUT.n107 OUT.n1 0.000532943
R518 OUT.n96 OUT.n95 0.000521962
R519 OUT.n76 OUT.n6 0.000510981
R520 OUT.n96 OUT.n6 0.000510981
R521 OUT.n95 OUT.n15 0.000510981
R522 OUT.n52 OUT.n15 0.000510981
R523 OUT.n52 OUT.n1 0.000510981
R524 ADJ.t35 ADJ.n4 620.038
R525 ADJ.t2 ADJ.n25 620.038
R526 ADJ.t11 ADJ.n35 620.038
R527 ADJ.n57 ADJ.t44 620.038
R528 ADJ.t31 ADJ.n69 620.006
R529 ADJ.t36 ADJ.n51 620.006
R530 ADJ.n14 ADJ.t9 620.006
R531 ADJ.t7 ADJ.n36 620.006
R532 ADJ.n14 ADJ.t3 619.74
R533 ADJ.n25 ADJ.t38 619.74
R534 ADJ.t28 ADJ.n15 619.74
R535 ADJ.t22 ADJ.n12 619.74
R536 ADJ.t30 ADJ.n9 619.74
R537 ADJ.t27 ADJ.n3 619.74
R538 ADJ.n68 ADJ.t13 619.74
R539 ADJ.n79 ADJ.t19 619.74
R540 ADJ.n69 ADJ.t34 619.74
R541 ADJ.t43 ADJ.n4 619.74
R542 ADJ.t5 ADJ.n35 619.74
R543 ADJ.n36 ADJ.t37 619.74
R544 ADJ.n48 ADJ.t20 619.74
R545 ADJ.n64 ADJ.t14 619.74
R546 ADJ.t15 ADJ.n58 619.74
R547 ADJ.t10 ADJ.n31 619.74
R548 ADJ.n57 ADJ.t21 619.74
R549 ADJ.n51 ADJ.t16 619.74
R550 ADJ.t32 ADJ.n30 619.74
R551 ADJ.n47 ADJ.t40 619.74
R552 ADJ.t3 ADJ.n13 614.254
R553 ADJ.n13 ADJ.t33 614.254
R554 ADJ.n24 ADJ.t33 614.254
R555 ADJ.t38 ADJ.n24 614.254
R556 ADJ.n20 ADJ.t28 614.254
R557 ADJ.t18 ADJ.n20 614.254
R558 ADJ.n21 ADJ.t18 614.254
R559 ADJ.n21 ADJ.t22 614.254
R560 ADJ.n17 ADJ.t30 614.254
R561 ADJ.n17 ADJ.t26 614.254
R562 ADJ.t26 ADJ.n16 614.254
R563 ADJ.n16 ADJ.t27 614.254
R564 ADJ.t13 ADJ.n67 614.254
R565 ADJ.n67 ADJ.t23 614.254
R566 ADJ.n78 ADJ.t23 614.254
R567 ADJ.t19 ADJ.n78 614.254
R568 ADJ.n74 ADJ.t34 614.254
R569 ADJ.t4 ADJ.n74 614.254
R570 ADJ.n75 ADJ.t4 614.254
R571 ADJ.n75 ADJ.t43 614.254
R572 ADJ.n70 ADJ.t35 614.254
R573 ADJ.t41 ADJ.n26 614.254
R574 ADJ.n26 ADJ.t2 614.254
R575 ADJ.n27 ADJ.t9 614.254
R576 ADJ.n27 ADJ.t41 614.254
R577 ADJ.n71 ADJ.t31 614.254
R578 ADJ.n71 ADJ.t39 614.254
R579 ADJ.t39 ADJ.n70 614.254
R580 ADJ.n41 ADJ.t5 614.254
R581 ADJ.n42 ADJ.t37 614.254
R582 ADJ.n42 ADJ.t8 614.254
R583 ADJ.t8 ADJ.n41 614.254
R584 ADJ.n62 ADJ.t20 614.254
R585 ADJ.t14 ADJ.n63 614.254
R586 ADJ.n63 ADJ.t24 614.254
R587 ADJ.t24 ADJ.n62 614.254
R588 ADJ.n59 ADJ.t15 614.254
R589 ADJ.n49 ADJ.t10 614.254
R590 ADJ.n49 ADJ.t17 614.254
R591 ADJ.n59 ADJ.t17 614.254
R592 ADJ.t21 ADJ.n56 614.254
R593 ADJ.n55 ADJ.t16 614.254
R594 ADJ.t25 ADJ.n55 614.254
R595 ADJ.n56 ADJ.t25 614.254
R596 ADJ.n45 ADJ.t32 614.254
R597 ADJ.t42 ADJ.n45 614.254
R598 ADJ.n46 ADJ.t42 614.254
R599 ADJ.t40 ADJ.n46 614.254
R600 ADJ.n38 ADJ.t11 614.254
R601 ADJ.n38 ADJ.t12 614.254
R602 ADJ.t12 ADJ.n37 614.254
R603 ADJ.n37 ADJ.t7 614.254
R604 ADJ.n53 ADJ.t36 614.254
R605 ADJ.n53 ADJ.t6 614.254
R606 ADJ.t6 ADJ.n52 614.254
R607 ADJ.n52 ADJ.t44 614.254
R608 ADJ.t29 ADJ.n86 101.537
R609 ADJ.t0 ADJ.n83 101.079
R610 ADJ.n87 ADJ.t29 101.079
R611 ADJ.n84 ADJ.t0 101.076
R612 ADJ.n65 ADJ.n29 15.7436
R613 ADJ.n82 ADJ.n2 14.7961
R614 ADJ.n29 ADJ.n2 14.6668
R615 ADJ.n54 ADJ.n53 5.13335
R616 ADJ.n52 ADJ.n34 5.13335
R617 ADJ.n37 ADJ.n8 5.02611
R618 ADJ.n72 ADJ.n71 5.02611
R619 ADJ.n28 ADJ.n27 5.02611
R620 ADJ.n26 ADJ.n11 5.02611
R621 ADJ.n24 ADJ.n23 5.02611
R622 ADJ.n13 ADJ.n10 5.02611
R623 ADJ.n22 ADJ.n21 5.02611
R624 ADJ.n20 ADJ.n19 5.02611
R625 ADJ.n16 ADJ.n5 5.02611
R626 ADJ.n18 ADJ.n17 5.02611
R627 ADJ.n78 ADJ.n77 5.02611
R628 ADJ.n67 ADJ.n7 5.02611
R629 ADJ.n76 ADJ.n75 5.02611
R630 ADJ.n74 ADJ.n73 5.02611
R631 ADJ.n70 ADJ.n6 5.02611
R632 ADJ.n39 ADJ.n38 5.02611
R633 ADJ.n43 ADJ.n42 5.02611
R634 ADJ.n41 ADJ.n40 5.02611
R635 ADJ.n46 ADJ.n33 5.02611
R636 ADJ.n63 ADJ.n32 5.02611
R637 ADJ.n62 ADJ.n61 5.02611
R638 ADJ.n50 ADJ.n49 5.02611
R639 ADJ.n60 ADJ.n59 5.02611
R640 ADJ.n55 ADJ.n54 5.02611
R641 ADJ.n56 ADJ.n34 5.02611
R642 ADJ.n45 ADJ.n44 5.02611
R643 ADJ.n65 ADJ.n64 2.82526
R644 ADJ.n81 ADJ.n1 2.35383
R645 ADJ.n86 ADJ.n85 1.5858
R646 ADJ.n85 ADJ.n0 1.5511
R647 ADJ.n82 ADJ.n81 0.8605
R648 ADJ ADJ.n87 0.800244
R649 ADJ.n84 ADJ.n1 0.649885
R650 ADJ.n83 ADJ.n82 0.533174
R651 ADJ.n48 ADJ.n1 0.471929
R652 ADJ.n85 ADJ.t1 0.470597
R653 ADJ.n39 ADJ.n6 0.437096
R654 ADJ.n72 ADJ.n8 0.437096
R655 ADJ.n87 ADJ.n0 0.401314
R656 ADJ.n66 ADJ.n65 0.321929
R657 ADJ.n81 ADJ.n80 0.321929
R658 ADJ.n79 ADJ.n4 0.298623
R659 ADJ.n12 ADJ.n3 0.298623
R660 ADJ.n25 ADJ.n12 0.298623
R661 ADJ.n48 ADJ.n47 0.298623
R662 ADJ.n47 ADJ.n35 0.298623
R663 ADJ.n58 ADJ.n57 0.298623
R664 ADJ.n58 ADJ.n48 0.298623
R665 ADJ.n80 ADJ.n79 0.295483
R666 ADJ.n15 ADJ.n14 0.26697
R667 ADJ.n15 ADJ.n9 0.26697
R668 ADJ.n69 ADJ.n68 0.26697
R669 ADJ.n36 ADJ.n30 0.26697
R670 ADJ.n64 ADJ.n30 0.26697
R671 ADJ.n64 ADJ.n31 0.26697
R672 ADJ.n51 ADJ.n31 0.26697
R673 ADJ.n68 ADJ.n66 0.26383
R674 ADJ.n11 ADJ.n2 0.148426
R675 ADJ.n29 ADJ.n28 0.148426
R676 ADJ.n83 ADJ.n0 0.1355
R677 ADJ.n86 ADJ.n84 0.120962
R678 ADJ.n23 ADJ.n11 0.107734
R679 ADJ.n23 ADJ.n22 0.107734
R680 ADJ.n22 ADJ.n5 0.107734
R681 ADJ.n77 ADJ.n5 0.107734
R682 ADJ.n77 ADJ.n76 0.107734
R683 ADJ.n76 ADJ.n6 0.107734
R684 ADJ.n40 ADJ.n39 0.107734
R685 ADJ.n40 ADJ.n33 0.107734
R686 ADJ.n61 ADJ.n33 0.107734
R687 ADJ.n61 ADJ.n60 0.107734
R688 ADJ.n60 ADJ.n34 0.107734
R689 ADJ.n28 ADJ.n10 0.107734
R690 ADJ.n19 ADJ.n10 0.107734
R691 ADJ.n19 ADJ.n18 0.107734
R692 ADJ.n18 ADJ.n7 0.107734
R693 ADJ.n73 ADJ.n7 0.107734
R694 ADJ.n73 ADJ.n72 0.107734
R695 ADJ.n43 ADJ.n8 0.107734
R696 ADJ.n44 ADJ.n43 0.107734
R697 ADJ.n44 ADJ.n32 0.107734
R698 ADJ.n50 ADJ.n32 0.107734
R699 ADJ.n54 ADJ.n50 0.107734
R700 ADJ.n80 ADJ.n3 0.00363953
R701 ADJ.n66 ADJ.n9 0.00363953
R702 VDD.t7 VDD.t13 4343.5
R703 VDD.t1 VDD.t7 4343.5
R704 VDD.n74 VDD.t1 2223.27
R705 VDD.n75 VDD.n3 180.601
R706 VDD.n92 VDD.n3 180.601
R707 VDD.n81 VDD.n8 180.601
R708 VDD.n8 VDD.n6 180.601
R709 VDD.n75 VDD.n7 147.525
R710 VDD.n6 VDD.n4 147.525
R711 VDD.n89 VDD.n3 135.8
R712 VDD.n89 VDD.n88 135.8
R713 VDD.n92 VDD.n4 135.8
R714 VDD.n81 VDD.n7 135.8
R715 VDD.n87 VDD.n86 135.8
R716 VDD.n86 VDD.n8 135.8
R717 VDD.n81 VDD.t50 119.879
R718 VDD.t0 VDD.n6 119.879
R719 VDD.t0 VDD.n5 119.683
R720 VDD.n74 VDD.t4 54.9597
R721 VDD.t22 VDD.n91 35.4234
R722 VDD.n54 VDD.n52 34.1113
R723 VDD.n31 VDD.n29 34.1107
R724 VDD.n66 VDD.n64 34.1107
R725 VDD.n39 VDD.n37 34.1085
R726 VDD.n46 VDD.n44 34.1085
R727 VDD.n60 VDD.n58 34.1074
R728 VDD.n88 VDD.n7 33.0755
R729 VDD.n87 VDD.n4 33.0755
R730 VDD.t4 VDD.t50 28.7682
R731 VDD.t0 VDD.t22 28.7682
R732 VDD.n92 VDD.t0 26.3889
R733 VDD.n42 VDD.n41 25.7991
R734 VDD.n35 VDD.n18 25.7912
R735 VDD.n50 VDD.n49 25.7893
R736 VDD.n67 VDD.n16 25.7873
R737 VDD.n32 VDD.n27 25.7854
R738 VDD.n56 VDD.n55 25.7854
R739 VDD.n91 VDD.n5 20.1034
R740 VDD.n90 VDD.t50 17.9501
R741 VDD.n19 VDD.n10 15.3535
R742 VDD.n80 VDD.n10 14.3237
R743 VDD.n91 VDD.n90 13.3893
R744 VDD.n88 VDD.n87 11.7255
R745 VDD.n20 VDD 11.1908
R746 VDD.n32 VDD.n31 6.59094
R747 VDD.n58 VDD.n56 6.59094
R748 VDD.n67 VDD.n66 6.58898
R749 VDD.n52 VDD.n50 6.58703
R750 VDD.n37 VDD.n35 6.58507
R751 VDD.n44 VDD.n42 6.57724
R752 VDD.n84 VDD.n82 4.0642
R753 VDD.n90 VDD.n89 3.71928
R754 VDD.n25 VDD.n24 3.34156
R755 VDD.n72 VDD.n71 3.08674
R756 VDD.n85 VDD.n9 3.06246
R757 VDD.n85 VDD.n84 3.06246
R758 VDD.n84 VDD.n83 2.52779
R759 VDD.n26 VDD.n21 2.48004
R760 VDD.n70 VDD.n13 2.29184
R761 VDD.n21 VDD.n20 1.65155
R762 VDD.n23 VDD.n22 1.6489
R763 VDD.n83 VDD.n2 1.5575
R764 VDD.n19 VDD.n13 1.52562
R765 VDD.n77 VDD.n11 1.5244
R766 VDD.n20 VDD.n19 1.03599
R767 VDD.n78 VDD.n1 0.98945
R768 VDD.n95 VDD.n1 0.98945
R769 VDD.n82 VDD.n80 0.970069
R770 VDD.n26 VDD.n25 0.862023
R771 VDD.n72 VDD.n70 0.795398
R772 VDD.n79 VDD.n78 0.695065
R773 VDD.n9 VDD.n2 0.695065
R774 VDD.n93 VDD.n2 0.6357
R775 VDD.n94 VDD.n93 0.6265
R776 VDD.n76 VDD.n0 0.380551
R777 VDD.n1 VDD.t23 0.303833
R778 VDD.n76 VDD.t5 0.303833
R779 VDD.n79 VDD.n77 0.27616
R780 VDD.n78 VDD.n9 0.262674
R781 VDD.n22 VDD 0.262078
R782 VDD.n80 VDD.n79 0.261707
R783 VDD VDD.n96 0.217474
R784 VDD.n83 VDD.n6 0.197375
R785 VDD.n93 VDD.n92 0.197375
R786 VDD.n76 VDD.n75 0.197375
R787 VDD.n75 VDD.n74 0.197375
R788 VDD.n82 VDD.n81 0.197375
R789 VDD.n86 VDD.n85 0.197375
R790 VDD.n86 VDD.n5 0.197375
R791 VDD.n89 VDD.n1 0.197375
R792 VDD.n95 VDD.n94 0.13595
R793 VDD.n96 VDD.n95 0.110525
R794 VDD.n77 VDD.n76 0.108972
R795 VDD.n33 VDD.n26 0.0547889
R796 VDD.n50 VDD.n15 0.0547889
R797 VDD.n56 VDD.n15 0.0505
R798 VDD.n68 VDD.n67 0.0505
R799 VDD.n42 VDD.n14 0.0505
R800 VDD.n35 VDD.n34 0.0505
R801 VDD.n33 VDD.n32 0.0505
R802 VDD.n22 VDD.n0 0.0499188
R803 VDD.n61 VDD.n54 0.0470525
R804 VDD.n29 VDD.n17 0.043625
R805 VDD.n64 VDD.n62 0.043625
R806 VDD.n24 VDD.t49 0.0431131
R807 VDD.n25 VDD.t10 0.0431131
R808 VDD.n21 VDD.t42 0.0431131
R809 VDD.n71 VDD.t40 0.0431131
R810 VDD.n72 VDD.t39 0.0431131
R811 VDD.n13 VDD.t44 0.0431131
R812 VDD.n40 VDD.n39 0.038
R813 VDD.n47 VDD.n46 0.038
R814 VDD.n61 VDD.n60 0.0351875
R815 VDD.n23 VDD.n17 0.0259588
R816 VDD.n94 VDD 0.0257
R817 VDD.n31 VDD.n30 0.0249131
R818 VDD.n29 VDD.n28 0.0249131
R819 VDD.n37 VDD.n36 0.0249131
R820 VDD.n39 VDD.n38 0.0249131
R821 VDD.n44 VDD.n43 0.0249131
R822 VDD.n46 VDD.n45 0.0249131
R823 VDD.n66 VDD.n65 0.0249131
R824 VDD.n64 VDD.n63 0.0249131
R825 VDD.n58 VDD.n57 0.0249131
R826 VDD.n60 VDD.n59 0.0249131
R827 VDD.n54 VDD.n53 0.0249131
R828 VDD.n52 VDD.n51 0.0249131
R829 VDD.n25 VDD.n12 0.0210046
R830 VDD.n72 VDD.n12 0.0210046
R831 VDD.n73 VDD.n72 0.0210046
R832 VDD.n73 VDD.n10 0.0210046
R833 VDD.n96 VDD.n0 0.0197986
R834 VDD.n51 VDD.t27 0.0187
R835 VDD.n51 VDD.t45 0.0187
R836 VDD.n53 VDD.t30 0.0187
R837 VDD.n53 VDD.t2 0.0187
R838 VDD.n28 VDD.t12 0.0187
R839 VDD.n28 VDD.t29 0.0187
R840 VDD.n30 VDD.t18 0.0187
R841 VDD.n30 VDD.t33 0.0187
R842 VDD.n27 VDD.t48 0.0187
R843 VDD.n27 VDD.t25 0.0187
R844 VDD.n38 VDD.t26 0.0187
R845 VDD.n38 VDD.t32 0.0187
R846 VDD.n36 VDD.t24 0.0187
R847 VDD.n36 VDD.t8 0.0187
R848 VDD.n18 VDD.t21 0.0187
R849 VDD.n18 VDD.t38 0.0187
R850 VDD.n45 VDD.t3 0.0187
R851 VDD.n45 VDD.t16 0.0187
R852 VDD.n43 VDD.t47 0.0187
R853 VDD.n43 VDD.t11 0.0187
R854 VDD.n41 VDD.t17 0.0187
R855 VDD.n41 VDD.t20 0.0187
R856 VDD.n63 VDD.t46 0.0187
R857 VDD.n63 VDD.t6 0.0187
R858 VDD.n65 VDD.t43 0.0187
R859 VDD.n65 VDD.t9 0.0187
R860 VDD.n16 VDD.t14 0.0187
R861 VDD.n16 VDD.t19 0.0187
R862 VDD.n59 VDD.t31 0.0187
R863 VDD.n59 VDD.t36 0.0187
R864 VDD.n57 VDD.t28 0.0187
R865 VDD.n57 VDD.t34 0.0187
R866 VDD.n55 VDD.t37 0.0187
R867 VDD.n55 VDD.t41 0.0187
R868 VDD.n49 VDD.t35 0.0187
R869 VDD.n49 VDD.t15 0.0187
R870 VDD.n70 VDD.n69 0.00883333
R871 VDD.n69 VDD.n68 0.007278
R872 VDD.n69 VDD.n14 0.00674189
R873 VDD.n34 VDD.n33 0.00478891
R874 VDD.n34 VDD.n14 0.00478891
R875 VDD.n68 VDD.n15 0.00478891
R876 VDD.n48 VDD.n11 0.00473203
R877 VDD.n62 VDD.n48 0.00406655
R878 VDD.n48 VDD.n47 0.00401084
R879 VDD.n24 VDD.n23 0.0031422
R880 VDD.n40 VDD.n17 0.00252126
R881 VDD.n47 VDD.n40 0.00252126
R882 VDD.n62 VDD.n61 0.00252126
R883 VDD.n71 VDD.n11 0.00172034
R884 VDD.t7 VDD.n12 0.00150004
R885 VDD.t7 VDD.n73 0.00150004
R886 a_30739_5010.n1 a_30739_5010.t3 39.1381
R887 a_30739_5010.n0 a_30739_5010.t1 36.2918
R888 a_30739_5010.t0 a_30739_5010.n1 3.29486
R889 a_30739_5010.n1 a_30739_5010.n0 0.643925
R890 a_30739_5010.n0 a_30739_5010.t2 0.608291
R891 MINUS MINUS.t0 50.8861
R892 a_30873_8186.t0 a_30873_8186.n0 3.08975
R893 a_30873_8186.n0 a_30873_8186.t2 0.551973
R894 a_30873_8186.n0 a_30873_8186.t1 0.545657
R895 PLUS PLUS.t0 53.5843
C0 PLUS ADJ 0.01871f
C1 OUT ADJ 58.5278f
C2 PLUS VDD 0.61561f
C3 MINUS ADJ 0
C4 OUT VDD 0.35828p
C5 MINUS VDD 0.56059f
C6 PLUS OUT 0
C7 VDD ADJ 0.10657p
C8 MINUS PLUS 0.27424f
C9 PLUS VSS 3.93904f
C10 MINUS VSS 4.22738f
C11 OUT VSS 0.49643p
C12 ADJ VSS 13.30631f
C13 VDD VSS 0.9838p
C14 PLUS.t0 VSS 1.62309f
C15 a_30873_8186.t1 VSS 1.48083f
C16 a_30873_8186.t2 VSS 1.47213f
C17 a_30873_8186.n0 VSS 6.7289f
C18 a_30873_8186.t0 VSS 2.81814f
C19 MINUS.t0 VSS 1.83269f
C20 a_30739_5010.t3 VSS 0.48774f
C21 a_30739_5010.t2 VSS 0.62068f
C22 a_30739_5010.t1 VSS 0.43386f
C23 a_30739_5010.n0 VSS 1.14289f
C24 a_30739_5010.n1 VSS 1.69797f
C25 a_30739_5010.t0 VSS 1.11687f
C26 VDD.n0 VSS 0.28161f
C27 VDD.t23 VSS 0.14226f
C28 VDD.n1 VSS 0.35592f
C29 VDD.n2 VSS 0.21733f
C30 VDD.n3 VSS 0.17235f
C31 VDD.n4 VSS 0.10964f
C32 VDD.n5 VSS 0.26449f
C33 VDD.n6 VSS 0.45855f
C34 VDD.t50 VSS 0.90884f
C35 VDD.n7 VSS 0.10964f
C36 VDD.n8 VSS 0.17235f
C37 VDD.n9 VSS 0.03907f
C38 VDD.n10 VSS 6.93115f
C39 VDD.n11 VSS 2.4395f
C40 VDD.t5 VSS 0.14226f
C41 VDD.t13 VSS 78.7837f
C42 VDD.n12 VSS 3.5516f
C43 VDD.t44 VSS 1.01768f
C44 VDD.n13 VSS 6.54263f
C45 VDD.n14 VSS 4.27663f
C46 VDD.n15 VSS 5.40276f
C47 VDD.t14 VSS 0.4301f
C48 VDD.t19 VSS 0.4301f
C49 VDD.n16 VSS 1.51055f
C50 VDD.n17 VSS 11.8093f
C51 VDD.t21 VSS 0.4301f
C52 VDD.t38 VSS 0.4301f
C53 VDD.n18 VSS 1.51058f
C54 VDD.n19 VSS 5.20137f
C55 VDD.n20 VSS 15.3164f
C56 VDD.t42 VSS 1.01768f
C57 VDD.n21 VSS 6.07568f
C58 VDD.t10 VSS 1.01768f
C59 VDD.n22 VSS 2.66338f
C60 VDD.n23 VSS 2.61366f
C61 VDD.t49 VSS 1.01768f
C62 VDD.n24 VSS 5.0017f
C63 VDD.n25 VSS 8.13183f
C64 VDD.n26 VSS 4.73083f
C65 VDD.t48 VSS 0.4301f
C66 VDD.t25 VSS 0.4301f
C67 VDD.n27 VSS 1.51053f
C68 VDD.t12 VSS 0.4301f
C69 VDD.t29 VSS 0.4301f
C70 VDD.n28 VSS 0.8602f
C71 VDD.n29 VSS 0.82073f
C72 VDD.t18 VSS 0.4301f
C73 VDD.t33 VSS 0.4301f
C74 VDD.n30 VSS 0.8602f
C75 VDD.n31 VSS 0.52642f
C76 VDD.n32 VSS 0.58968f
C77 VDD.n33 VSS 5.47438f
C78 VDD.n34 VSS 3.48351f
C79 VDD.n35 VSS 0.58961f
C80 VDD.t24 VSS 0.4301f
C81 VDD.t8 VSS 0.4301f
C82 VDD.n36 VSS 0.8602f
C83 VDD.n37 VSS 0.52646f
C84 VDD.t26 VSS 0.4301f
C85 VDD.t32 VSS 0.4301f
C86 VDD.n38 VSS 0.8602f
C87 VDD.n39 VSS 0.86345f
C88 VDD.n40 VSS 7.58915f
C89 VDD.t17 VSS 0.4301f
C90 VDD.t20 VSS 0.4301f
C91 VDD.n41 VSS 1.51065f
C92 VDD.n42 VSS 0.58952f
C93 VDD.t47 VSS 0.4301f
C94 VDD.t11 VSS 0.4301f
C95 VDD.n43 VSS 0.8602f
C96 VDD.n44 VSS 0.52647f
C97 VDD.t3 VSS 0.4301f
C98 VDD.t16 VSS 0.4301f
C99 VDD.n45 VSS 0.8602f
C100 VDD.n46 VSS 0.86345f
C101 VDD.n47 VSS 10.5358f
C102 VDD.n48 VSS 9.45918f
C103 VDD.t35 VSS 0.4301f
C104 VDD.t15 VSS 0.4301f
C105 VDD.n49 VSS 1.51056f
C106 VDD.n50 VSS 0.75426f
C107 VDD.t27 VSS 0.4301f
C108 VDD.t45 VSS 0.4301f
C109 VDD.n51 VSS 0.8602f
C110 VDD.n52 VSS 0.52642f
C111 VDD.t30 VSS 0.4301f
C112 VDD.t2 VSS 0.4301f
C113 VDD.n53 VSS 0.8602f
C114 VDD.n54 VSS 1.01887f
C115 VDD.t37 VSS 0.4301f
C116 VDD.t41 VSS 0.4301f
C117 VDD.n55 VSS 1.51053f
C118 VDD.n56 VSS 0.58968f
C119 VDD.t28 VSS 0.4301f
C120 VDD.t34 VSS 0.4301f
C121 VDD.n57 VSS 0.8602f
C122 VDD.n58 VSS 0.52646f
C123 VDD.t31 VSS 0.4301f
C124 VDD.t36 VSS 0.4301f
C125 VDD.n59 VSS 0.8602f
C126 VDD.n60 VSS 0.89002f
C127 VDD.n61 VSS 12.1257f
C128 VDD.n62 VSS 10.2736f
C129 VDD.t46 VSS 0.4301f
C130 VDD.t6 VSS 0.4301f
C131 VDD.n63 VSS 0.8602f
C132 VDD.n64 VSS 0.82073f
C133 VDD.t43 VSS 0.4301f
C134 VDD.t9 VSS 0.4301f
C135 VDD.n65 VSS 0.8602f
C136 VDD.n66 VSS 0.52643f
C137 VDD.n67 VSS 0.58966f
C138 VDD.n68 VSS 4.49435f
C139 VDD.n69 VSS 5.28747f
C140 VDD.n70 VSS 4.93657f
C141 VDD.t40 VSS 1.01768f
C142 VDD.n71 VSS 5.37657f
C143 VDD.t39 VSS 1.01768f
C144 VDD.n72 VSS 10.5618f
C145 VDD.n73 VSS 3.5516f
C146 VDD.t7 VSS 77.94771f
C147 VDD.t1 VSS 58.9231f
C148 VDD.t4 VSS 0.75128f
C149 VDD.n74 VSS 20.4424f
C150 VDD.n75 VSS 0.11236f
C151 VDD.n76 VSS 0.36201f
C152 VDD.n77 VSS 2.7633f
C153 VDD.n78 VSS 0.08816f
C154 VDD.n79 VSS 0.27417f
C155 VDD.n80 VSS 2.58235f
C156 VDD.n81 VSS 0.6063f
C157 VDD.n82 VSS 0.0495f
C158 VDD.n83 VSS 0.14582f
C159 VDD.n84 VSS 0.12324f
C160 VDD.n85 VSS 0.05954f
C161 VDD.n86 VSS 0.09242f
C162 VDD.n87 VSS 0.06146f
C163 VDD.n88 VSS 0.06146f
C164 VDD.n89 VSS 0.48101f
C165 VDD.n90 VSS 0.02172f
C166 VDD.n91 VSS 0.7196f
C167 VDD.t22 VSS 0.57598f
C168 VDD.t0 VSS 0.95419f
C169 VDD.n92 VSS 1.1139f
C170 VDD.n93 VSS 0.29339f
C171 VDD.n94 VSS 0.26373f
C172 VDD.n95 VSS 0.25934f
C173 VDD.n96 VSS 0.35123f
C174 ADJ.n0 VSS 0.11786f
C175 ADJ.n1 VSS 0.22005f
C176 ADJ.n2 VSS 3.64599f
C177 ADJ.n3 VSS 0.88061f
C178 ADJ.n4 VSS 1.77917f
C179 ADJ.t23 VSS 1.75524f
C180 ADJ.n5 VSS 0.07387f
C181 ADJ.n6 VSS 0.16755f
C182 ADJ.t34 VSS 1.76298f
C183 ADJ.n7 VSS 0.07387f
C184 ADJ.n8 VSS 0.16755f
C185 ADJ.n9 VSS 0.88155f
C186 ADJ.n10 VSS 0.07387f
C187 ADJ.t9 VSS 1.76336f
C188 ADJ.n11 VSS 0.08544f
C189 ADJ.n12 VSS 0.89195f
C190 ADJ.t33 VSS 1.75524f
C191 ADJ.n13 VSS 1.77217f
C192 ADJ.t3 VSS 1.76298f
C193 ADJ.n14 VSS 1.78203f
C194 ADJ.n15 VSS 0.89383f
C195 ADJ.t28 VSS 1.76298f
C196 ADJ.t30 VSS 1.76298f
C197 ADJ.t27 VSS 1.76298f
C198 ADJ.n16 VSS 1.77217f
C199 ADJ.t26 VSS 1.75524f
C200 ADJ.n17 VSS 1.77217f
C201 ADJ.n18 VSS 0.07387f
C202 ADJ.n19 VSS 0.07387f
C203 ADJ.n20 VSS 1.77217f
C204 ADJ.t18 VSS 1.75524f
C205 ADJ.t22 VSS 1.76298f
C206 ADJ.n21 VSS 1.77217f
C207 ADJ.n22 VSS 0.07387f
C208 ADJ.n23 VSS 0.07387f
C209 ADJ.n24 VSS 1.77217f
C210 ADJ.t38 VSS 1.76298f
C211 ADJ.n25 VSS 1.77917f
C212 ADJ.t2 VSS 1.76341f
C213 ADJ.n26 VSS 1.77217f
C214 ADJ.t41 VSS 1.75524f
C215 ADJ.n27 VSS 1.77217f
C216 ADJ.n28 VSS 0.08544f
C217 ADJ.n29 VSS 3.75721f
C218 ADJ.n30 VSS 0.89383f
C219 ADJ.n31 VSS 0.89383f
C220 ADJ.n32 VSS 0.07387f
C221 ADJ.t20 VSS 1.76298f
C222 ADJ.n33 VSS 0.07387f
C223 ADJ.n34 VSS 0.13073f
C224 ADJ.t17 VSS 1.75524f
C225 ADJ.n35 VSS 1.77917f
C226 ADJ.t32 VSS 1.76298f
C227 ADJ.t37 VSS 1.76298f
C228 ADJ.t5 VSS 1.76298f
C229 ADJ.n36 VSS 1.78203f
C230 ADJ.t7 VSS 1.76336f
C231 ADJ.n37 VSS 1.77217f
C232 ADJ.t12 VSS 1.75524f
C233 ADJ.t11 VSS 1.76341f
C234 ADJ.n38 VSS 1.77217f
C235 ADJ.n39 VSS 0.16755f
C236 ADJ.n40 VSS 0.07387f
C237 ADJ.n41 VSS 1.77217f
C238 ADJ.t8 VSS 1.75524f
C239 ADJ.n42 VSS 1.77217f
C240 ADJ.n43 VSS 0.07387f
C241 ADJ.n44 VSS 0.07387f
C242 ADJ.n45 VSS 1.77217f
C243 ADJ.t42 VSS 1.75524f
C244 ADJ.n46 VSS 1.77217f
C245 ADJ.t40 VSS 1.76298f
C246 ADJ.n47 VSS 0.89195f
C247 ADJ.n48 VSS 0.92265f
C248 ADJ.t44 VSS 1.76341f
C249 ADJ.t16 VSS 1.76298f
C250 ADJ.t10 VSS 1.76298f
C251 ADJ.n49 VSS 1.77217f
C252 ADJ.n50 VSS 0.07387f
C253 ADJ.n51 VSS 1.78203f
C254 ADJ.t36 VSS 1.76336f
C255 ADJ.n52 VSS 1.77339f
C256 ADJ.t6 VSS 1.75524f
C257 ADJ.n53 VSS 1.77338f
C258 ADJ.n54 VSS 0.13046f
C259 ADJ.n55 VSS 1.77217f
C260 ADJ.t25 VSS 1.75524f
C261 ADJ.n56 VSS 1.77217f
C262 ADJ.t21 VSS 1.76298f
C263 ADJ.n57 VSS 1.77917f
C264 ADJ.n58 VSS 0.89195f
C265 ADJ.t15 VSS 1.76298f
C266 ADJ.n59 VSS 1.77217f
C267 ADJ.n60 VSS 0.07387f
C268 ADJ.n61 VSS 0.07387f
C269 ADJ.n62 VSS 1.77217f
C270 ADJ.t24 VSS 1.75524f
C271 ADJ.n63 VSS 1.77217f
C272 ADJ.t14 VSS 1.76298f
C273 ADJ.n64 VSS 1.0903f
C274 ADJ.n65 VSS 1.94415f
C275 ADJ.n66 VSS 0.01243f
C276 ADJ.n67 VSS 1.77217f
C277 ADJ.t13 VSS 1.76298f
C278 ADJ.n68 VSS 0.89368f
C279 ADJ.n69 VSS 1.78203f
C280 ADJ.t31 VSS 1.76336f
C281 ADJ.t35 VSS 1.76341f
C282 ADJ.n70 VSS 1.77217f
C283 ADJ.t39 VSS 1.75524f
C284 ADJ.n71 VSS 1.77217f
C285 ADJ.n72 VSS 0.16755f
C286 ADJ.n73 VSS 0.07387f
C287 ADJ.n74 VSS 1.77217f
C288 ADJ.t4 VSS 1.75524f
C289 ADJ.t43 VSS 1.76298f
C290 ADJ.n75 VSS 1.77217f
C291 ADJ.n76 VSS 0.07387f
C292 ADJ.n77 VSS 0.07387f
C293 ADJ.n78 VSS 1.77217f
C294 ADJ.t19 VSS 1.76298f
C295 ADJ.n79 VSS 0.89183f
C296 ADJ.n80 VSS 0.01146f
C297 ADJ.n81 VSS 0.16966f
C298 ADJ.n82 VSS 1.88106f
C299 ADJ.n83 VSS 0.1651f
C300 ADJ.t0 VSS 0.28679f
C301 ADJ.n84 VSS 0.15154f
C302 ADJ.t1 VSS 0.3793f
C303 ADJ.n85 VSS 0.41068f
C304 ADJ.n86 VSS 0.25898f
C305 ADJ.t29 VSS 0.28746f
C306 ADJ.n87 VSS 0.19588f
C307 OUT.n0 VSS 8.38911f
C308 OUT.n1 VSS 0.02015f
C309 OUT.t40 VSS 1.79539f
C310 OUT.n2 VSS 1.93766f
C311 OUT.t20 VSS 1.81058f
C312 OUT.t31 VSS 3.13457f
C313 OUT.n3 VSS 5.177f
C314 OUT.n4 VSS 5.177f
C315 OUT.t5 VSS 0.63926f
C316 OUT.t3 VSS 0.63926f
C317 OUT.n5 VSS 1.27851f
C318 OUT.n6 VSS 0.1598f
C319 OUT.t60 VSS 0.63926f
C320 OUT.t80 VSS 0.63926f
C321 OUT.n7 VSS 1.27851f
C322 OUT.n8 VSS 1.45226f
C323 OUT.t16 VSS 0.63926f
C324 OUT.t14 VSS 0.63926f
C325 OUT.n9 VSS 1.39288f
C326 OUT.t36 VSS 0.63926f
C327 OUT.t24 VSS 0.63926f
C328 OUT.n10 VSS 2.25109f
C329 OUT.n11 VSS 0.75674f
C330 OUT.t4 VSS 0.63926f
C331 OUT.t39 VSS 0.63926f
C332 OUT.n12 VSS 1.27851f
C333 OUT.n13 VSS 0.75786f
C334 OUT.n14 VSS 1.45522f
C335 OUT.n15 VSS 0.01008f
C336 OUT.t13 VSS 1.60095f
C337 OUT.t18 VSS 3.13449f
C338 OUT.t62 VSS 0.63926f
C339 OUT.t72 VSS 0.63926f
C340 OUT.n16 VSS 2.25101f
C341 OUT.t53 VSS 0.63926f
C342 OUT.t65 VSS 0.63926f
C343 OUT.n17 VSS 1.27851f
C344 OUT.n18 VSS 0.75784f
C345 OUT.t58 VSS 0.63926f
C346 OUT.t70 VSS 0.63926f
C347 OUT.n19 VSS 2.25109f
C348 OUT.n20 VSS 0.7568f
C349 OUT.n21 VSS 5.177f
C350 OUT.t68 VSS 1.62033f
C351 OUT.n22 VSS 1.30112f
C352 OUT.t74 VSS 3.13452f
C353 OUT.n23 VSS 1.00038f
C354 OUT.t79 VSS 0.63926f
C355 OUT.t43 VSS 0.63926f
C356 OUT.n24 VSS 1.27851f
C357 OUT.n25 VSS 1.42062f
C358 OUT.t64 VSS 0.63926f
C359 OUT.t75 VSS 0.63926f
C360 OUT.n26 VSS 1.27851f
C361 OUT.n27 VSS 0.75786f
C362 OUT.t69 VSS 0.63926f
C363 OUT.t78 VSS 0.63926f
C364 OUT.n28 VSS 2.25101f
C365 OUT.n29 VSS 0.75685f
C366 OUT.n30 VSS 7.99734f
C367 OUT.t57 VSS 0.63926f
C368 OUT.t59 VSS 0.63926f
C369 OUT.n31 VSS 1.31375f
C370 OUT.t77 VSS 0.63926f
C371 OUT.t54 VSS 0.63926f
C372 OUT.n32 VSS 1.31375f
C373 OUT.t67 VSS 0.63926f
C374 OUT.t49 VSS 0.63926f
C375 OUT.n33 VSS 2.25111f
C376 OUT.n34 VSS 6.12458f
C377 OUT.n35 VSS 0.75678f
C378 OUT.t63 VSS 0.63926f
C379 OUT.t45 VSS 0.63926f
C380 OUT.n36 VSS 1.27851f
C381 OUT.n37 VSS 0.75783f
C382 OUT.n38 VSS 1.53453f
C383 OUT.t33 VSS 0.63926f
C384 OUT.t26 VSS 0.63926f
C385 OUT.n39 VSS 1.42385f
C386 OUT.t8 VSS 0.63926f
C387 OUT.t1 VSS 0.63926f
C388 OUT.n40 VSS 2.25114f
C389 OUT.t23 VSS 0.63926f
C390 OUT.t37 VSS 0.63926f
C391 OUT.n41 VSS 1.45204f
C392 OUT.n42 VSS 1.39589f
C393 OUT.t30 VSS 0.63926f
C394 OUT.t32 VSS 0.63926f
C395 OUT.n43 VSS 1.27851f
C396 OUT.n44 VSS 0.75782f
C397 OUT.t17 VSS 0.63926f
C398 OUT.t25 VSS 0.63926f
C399 OUT.n45 VSS 2.25106f
C400 OUT.n46 VSS 1.04253f
C401 OUT.n47 VSS 8.5082f
C402 OUT.n48 VSS 0.7567f
C403 OUT.t15 VSS 0.63926f
C404 OUT.t7 VSS 0.63926f
C405 OUT.n49 VSS 1.27851f
C406 OUT.n50 VSS 0.75782f
C407 OUT.n51 VSS 1.42417f
C408 OUT.n52 VSS 0.01008f
C409 OUT.n53 VSS 1.53453f
C410 OUT.t47 VSS 0.63926f
C411 OUT.t52 VSS 0.63926f
C412 OUT.n54 VSS 1.27851f
C413 OUT.n55 VSS 0.75783f
C414 OUT.t50 VSS 0.63926f
C415 OUT.t55 VSS 0.63926f
C416 OUT.n56 VSS 2.25111f
C417 OUT.n57 VSS 0.75678f
C418 OUT.n58 VSS 5.177f
C419 OUT.t42 VSS 0.63926f
C420 OUT.t48 VSS 0.63926f
C421 OUT.n59 VSS 1.34592f
C422 OUT.n60 VSS 1.50227f
C423 OUT.t71 VSS 0.63926f
C424 OUT.t41 VSS 0.63926f
C425 OUT.n61 VSS 1.27851f
C426 OUT.n62 VSS 0.75782f
C427 OUT.t76 VSS 0.63926f
C428 OUT.t44 VSS 0.63926f
C429 OUT.n63 VSS 2.25109f
C430 OUT.n64 VSS 0.7568f
C431 OUT.n65 VSS 7.86373f
C432 OUT.t56 VSS 1.62033f
C433 OUT.n66 VSS 2.11317f
C434 OUT.t46 VSS 1.62033f
C435 OUT.n67 VSS 1.30327f
C436 OUT.t51 VSS 3.13396f
C437 OUT.n68 VSS 0.76848f
C438 OUT.n69 VSS 7.85795f
C439 OUT.n70 VSS 5.17122f
C440 OUT.n71 VSS 0.75685f
C441 OUT.t61 VSS 0.63926f
C442 OUT.t66 VSS 0.63926f
C443 OUT.n72 VSS 1.27851f
C444 OUT.n73 VSS 0.75785f
C445 OUT.t73 VSS 0.63926f
C446 OUT.t81 VSS 0.63926f
C447 OUT.n74 VSS 1.27851f
C448 OUT.n75 VSS 1.39189f
C449 OUT.n76 VSS 0.19873f
C450 OUT.t0 VSS 0.63926f
C451 OUT.t38 VSS 0.63926f
C452 OUT.n77 VSS 2.25106f
C453 OUT.n78 VSS 0.75675f
C454 OUT.t12 VSS 0.63926f
C455 OUT.t27 VSS 0.63926f
C456 OUT.n79 VSS 1.27851f
C457 OUT.n80 VSS 0.75789f
C458 OUT.t6 VSS 0.63926f
C459 OUT.t28 VSS 0.63926f
C460 OUT.n81 VSS 1.27851f
C461 OUT.n82 VSS 1.39189f
C462 OUT.n83 VSS 0.10061p
C463 OUT.t10 VSS 0.63926f
C464 OUT.t9 VSS 0.63926f
C465 OUT.n84 VSS 1.27851f
C466 OUT.n85 VSS 1.40771f
C467 OUT.t34 VSS 0.63926f
C468 OUT.t21 VSS 0.63926f
C469 OUT.n86 VSS 1.27851f
C470 OUT.n87 VSS 0.75789f
C471 OUT.t22 VSS 0.63926f
C472 OUT.t82 VSS 0.63926f
C473 OUT.n88 VSS 2.25101f
C474 OUT.n89 VSS 0.75679f
C475 OUT.n90 VSS 5.177f
C476 OUT.n91 VSS 4.05609f
C477 OUT.n92 VSS 0.75845f
C478 OUT.t11 VSS 1.51258f
C479 OUT.n93 VSS 1.40895f
C480 OUT.n94 VSS 2.13237f
C481 OUT.n95 VSS 0.01511f
C482 OUT.n96 VSS 0.13308f
C483 OUT.n97 VSS 1.56986f
C484 OUT.t35 VSS 0.63926f
C485 OUT.t29 VSS 0.63926f
C486 OUT.n98 VSS 1.27851f
C487 OUT.n99 VSS 0.75795f
C488 OUT.t2 VSS 0.63926f
C489 OUT.t83 VSS 0.63926f
C490 OUT.n100 VSS 2.25103f
C491 OUT.n101 VSS 0.75677f
C492 OUT.n102 VSS 7.85795f
C493 OUT.n103 VSS 7.85795f
C494 OUT.n104 VSS 0.7584f
C495 OUT.t19 VSS 1.51258f
C496 OUT.n105 VSS 1.40878f
C497 OUT.n106 VSS 1.92221f
C498 OUT.n107 VSS 50.1114f
C499 a_31459_5010.t1 VSS 0.1447f
C500 a_31459_5010.n0 VSS 0.28422f
C501 a_31459_5010.n1 VSS 0.39314f
C502 a_31459_5010.t13 VSS 0.77747f
C503 a_31459_5010.n2 VSS 0.7843f
C504 a_31459_5010.t22 VSS 0.77406f
C505 a_31459_5010.n3 VSS 0.03258f
C506 a_31459_5010.n4 VSS 0.07389f
C507 a_31459_5010.t2 VSS 0.77747f
C508 a_31459_5010.n5 VSS 0.03258f
C509 a_31459_5010.n6 VSS 0.07389f
C510 a_31459_5010.n7 VSS 0.39314f
C511 a_31459_5010.n8 VSS 0.06036f
C512 a_31459_5010.t23 VSS 0.77747f
C513 a_31459_5010.n9 VSS 0.78212f
C514 a_31459_5010.t20 VSS 0.77406f
C515 a_31459_5010.n10 VSS 0.78212f
C516 a_31459_5010.t6 VSS 0.77767f
C517 a_31459_5010.n11 VSS 0.7843f
C518 a_31459_5010.t29 VSS 0.77747f
C519 a_31459_5010.n12 VSS 0.78153f
C520 a_31459_5010.t38 VSS 0.77406f
C521 a_31459_5010.t16 VSS 0.77767f
C522 a_31459_5010.n13 VSS 0.7843f
C523 a_31459_5010.t34 VSS 0.77747f
C524 a_31459_5010.n14 VSS 0.78153f
C525 a_31459_5010.n15 VSS 0.06047f
C526 a_31459_5010.n16 VSS 0.03258f
C527 a_31459_5010.t25 VSS 0.77747f
C528 a_31459_5010.n17 VSS 0.78153f
C529 a_31459_5010.t30 VSS 0.77406f
C530 a_31459_5010.n18 VSS 0.78153f
C531 a_31459_5010.n19 VSS 0.03258f
C532 a_31459_5010.n20 VSS 0.03258f
C533 a_31459_5010.n21 VSS 0.78153f
C534 a_31459_5010.t18 VSS 0.77406f
C535 a_31459_5010.n22 VSS 0.78153f
C536 a_31459_5010.t3 VSS 0.77747f
C537 a_31459_5010.n23 VSS 1.65262f
C538 a_31459_5010.n24 VSS 0.39314f
C539 a_31459_5010.n25 VSS 0.39314f
C540 a_31459_5010.t31 VSS 0.77406f
C541 a_31459_5010.n26 VSS 0.03258f
C542 a_31459_5010.n27 VSS 0.03258f
C543 a_31459_5010.t4 VSS 0.77747f
C544 a_31459_5010.n28 VSS 0.03258f
C545 a_31459_5010.n29 VSS 0.39314f
C546 a_31459_5010.n30 VSS 0.07389f
C547 a_31459_5010.t42 VSS 0.77406f
C548 a_31459_5010.n31 VSS 0.03258f
C549 a_31459_5010.n32 VSS 0.78153f
C550 a_31459_5010.t35 VSS 0.77747f
C551 a_31459_5010.n33 VSS 0.7843f
C552 a_31459_5010.t41 VSS 0.77767f
C553 a_31459_5010.n34 VSS 0.78153f
C554 a_31459_5010.t12 VSS 0.77406f
C555 a_31459_5010.n35 VSS 0.78153f
C556 a_31459_5010.t7 VSS 0.77767f
C557 a_31459_5010.n36 VSS 0.7843f
C558 a_31459_5010.t39 VSS 0.77747f
C559 a_31459_5010.n37 VSS 0.78153f
C560 a_31459_5010.n38 VSS 0.03258f
C561 a_31459_5010.t26 VSS 0.77747f
C562 a_31459_5010.n39 VSS 0.78153f
C563 a_31459_5010.t36 VSS 0.77406f
C564 a_31459_5010.t33 VSS 0.77747f
C565 a_31459_5010.n40 VSS 0.78153f
C566 a_31459_5010.n41 VSS 0.03258f
C567 a_31459_5010.n42 VSS 0.03258f
C568 a_31459_5010.n43 VSS 0.78153f
C569 a_31459_5010.t28 VSS 0.77747f
C570 a_31459_5010.n44 VSS 0.39314f
C571 a_31459_5010.t9 VSS 0.77767f
C572 a_31459_5010.t8 VSS 0.77406f
C573 a_31459_5010.n45 VSS 0.8392f
C574 a_31459_5010.n46 VSS 1.63749f
C575 a_31459_5010.n47 VSS 0.78153f
C576 a_31459_5010.t40 VSS 0.77747f
C577 a_31459_5010.n48 VSS 0.7843f
C578 a_31459_5010.t43 VSS 0.77767f
C579 a_31459_5010.n49 VSS 0.03546f
C580 a_31459_5010.n50 VSS 0.78153f
C581 a_31459_5010.t15 VSS 0.77406f
C582 a_31459_5010.n51 VSS 0.78153f
C583 a_31459_5010.n52 VSS 0.03546f
C584 a_31459_5010.n53 VSS 0.03258f
C585 a_31459_5010.n54 VSS 0.78153f
C586 a_31459_5010.t5 VSS 0.77747f
C587 a_31459_5010.n55 VSS 0.7843f
C588 a_31459_5010.n56 VSS 0.39314f
C589 a_31459_5010.t14 VSS 0.77747f
C590 a_31459_5010.n57 VSS 0.78153f
C591 a_31459_5010.t19 VSS 0.77406f
C592 a_31459_5010.n58 VSS 0.78153f
C593 a_31459_5010.n59 VSS 0.03258f
C594 a_31459_5010.n60 VSS 0.03258f
C595 a_31459_5010.n61 VSS 0.78153f
C596 a_31459_5010.t24 VSS 0.77747f
C597 a_31459_5010.n62 VSS 0.39314f
C598 a_31459_5010.n63 VSS 0.85781f
C599 a_31459_5010.n64 VSS 0.479f
C600 a_31459_5010.n65 VSS 0.78153f
C601 a_31459_5010.t10 VSS 0.77747f
C602 a_31459_5010.n66 VSS 0.39314f
C603 a_31459_5010.n67 VSS 0.7843f
C604 a_31459_5010.t27 VSS 0.77767f
C605 a_31459_5010.t32 VSS 0.77767f
C606 a_31459_5010.n68 VSS 0.78153f
C607 a_31459_5010.t37 VSS 0.77406f
C608 a_31459_5010.n69 VSS 0.78153f
C609 a_31459_5010.n70 VSS 0.07389f
C610 a_31459_5010.n71 VSS 0.03258f
C611 a_31459_5010.n72 VSS 0.78153f
C612 a_31459_5010.t17 VSS 0.77406f
C613 a_31459_5010.t11 VSS 0.77747f
C614 a_31459_5010.n73 VSS 0.78153f
C615 a_31459_5010.n74 VSS 0.03258f
C616 a_31459_5010.n75 VSS 0.03258f
C617 a_31459_5010.n76 VSS 0.78153f
C618 a_31459_5010.t21 VSS 0.77747f
C619 a_31459_5010.n77 VSS 0.39314f
C620 a_31459_5010.n78 VSS 0.39314f
C621 a_31459_5010.n79 VSS 0.32084f
C622 a_31459_5010.t0 VSS 0.21982f
.ends

