magic
tech gf180mcuD
magscale 1 10
timestamp 1763828743
<< nwell >>
rect 298 4675 62677 9333
rect 298 2536 1544 4675
<< pwell >>
rect 1544 2536 62677 4675
rect 298 0 62677 2536
<< mvnmos >>
rect 1877 4173 21877 4293
rect 22109 4173 42109 4293
rect 42341 4173 62341 4293
rect 1877 3949 21877 4069
rect 22109 3949 42109 4069
rect 42341 3949 62341 4069
rect 1877 3725 21877 3845
rect 22109 3725 42109 3845
rect 42341 3725 62341 3845
rect 1877 3501 21877 3621
rect 22109 3501 42109 3621
rect 42341 3501 62341 3621
rect 1877 3277 21877 3397
rect 22109 3277 42109 3397
rect 42341 3277 62341 3397
rect 1877 3053 21877 3173
rect 22109 3053 42109 3173
rect 42341 3053 62341 3173
rect 1877 2829 21877 2949
rect 22109 2829 42109 2949
rect 42341 2829 62341 2949
rect 717 272 837 2272
rect 1229 272 1349 2272
rect 1877 1917 21877 2037
rect 22109 1917 42109 2037
rect 42341 1917 62341 2037
rect 1877 1693 21877 1813
rect 22109 1693 42109 1813
rect 42341 1693 62341 1813
rect 1877 1469 21877 1589
rect 22109 1469 42109 1589
rect 42341 1469 62341 1589
rect 1877 1245 21877 1365
rect 22109 1245 42109 1365
rect 42341 1245 62341 1365
rect 1877 1021 21877 1141
rect 22109 1021 42109 1141
rect 42341 1021 62341 1141
rect 1877 797 21877 917
rect 22109 797 42109 917
rect 42341 797 62341 917
rect 1877 573 21877 693
rect 22109 573 42109 693
rect 42341 573 62341 693
<< mvpmos >>
rect 696 5968 816 8768
rect 1208 5968 1328 8768
rect 1880 8639 21880 8759
rect 22112 8639 42112 8759
rect 42344 8639 62344 8759
rect 1880 8415 21880 8535
rect 22112 8415 42112 8535
rect 42344 8415 62344 8535
rect 1880 8191 21880 8311
rect 22112 8191 42112 8311
rect 42344 8191 62344 8311
rect 1880 7967 21880 8087
rect 22112 7967 42112 8087
rect 42344 7967 62344 8087
rect 1880 7743 21880 7863
rect 22112 7743 42112 7863
rect 42344 7743 62344 7863
rect 1880 7519 21880 7639
rect 22112 7519 42112 7639
rect 42344 7519 62344 7639
rect 1880 7295 21880 7415
rect 22112 7295 42112 7415
rect 42344 7295 62344 7415
rect 562 2792 682 5592
rect 1074 2792 1194 5592
rect 1880 6383 21880 6503
rect 22112 6383 42112 6503
rect 42344 6383 62344 6503
rect 1880 6159 21880 6279
rect 22112 6159 42112 6279
rect 42344 6159 62344 6279
rect 1880 5935 21880 6055
rect 22112 5935 42112 6055
rect 42344 5935 62344 6055
rect 1880 5711 21880 5831
rect 22112 5711 42112 5831
rect 42344 5711 62344 5831
rect 1880 5487 21880 5607
rect 22112 5487 42112 5607
rect 42344 5487 62344 5607
rect 1880 5263 21880 5383
rect 22112 5263 42112 5383
rect 42344 5263 62344 5383
rect 1880 5039 21880 5159
rect 22112 5039 42112 5159
rect 42344 5039 62344 5159
<< mvndiff >>
rect 1877 4368 21877 4381
rect 1877 4322 1890 4368
rect 21864 4322 21877 4368
rect 1877 4293 21877 4322
rect 22109 4368 42109 4381
rect 22109 4322 22122 4368
rect 42096 4322 42109 4368
rect 22109 4293 42109 4322
rect 42341 4368 62341 4381
rect 42341 4322 42354 4368
rect 62328 4322 62341 4368
rect 42341 4293 62341 4322
rect 1877 4144 21877 4173
rect 1877 4098 1890 4144
rect 21864 4098 21877 4144
rect 1877 4069 21877 4098
rect 22109 4144 42109 4173
rect 22109 4098 22122 4144
rect 42096 4098 42109 4144
rect 22109 4069 42109 4098
rect 42341 4144 62341 4173
rect 42341 4098 42354 4144
rect 62328 4098 62341 4144
rect 42341 4069 62341 4098
rect 1877 3920 21877 3949
rect 1877 3874 1890 3920
rect 21864 3874 21877 3920
rect 1877 3845 21877 3874
rect 22109 3920 42109 3949
rect 22109 3874 22122 3920
rect 42096 3874 42109 3920
rect 22109 3845 42109 3874
rect 42341 3920 62341 3949
rect 42341 3874 42354 3920
rect 62328 3874 62341 3920
rect 42341 3845 62341 3874
rect 1877 3696 21877 3725
rect 1877 3650 1890 3696
rect 21864 3650 21877 3696
rect 1877 3621 21877 3650
rect 22109 3696 42109 3725
rect 22109 3650 22122 3696
rect 42096 3650 42109 3696
rect 22109 3621 42109 3650
rect 42341 3696 62341 3725
rect 42341 3650 42354 3696
rect 62328 3650 62341 3696
rect 42341 3621 62341 3650
rect 1877 3472 21877 3501
rect 1877 3426 1890 3472
rect 21864 3426 21877 3472
rect 1877 3397 21877 3426
rect 22109 3472 42109 3501
rect 22109 3426 22122 3472
rect 42096 3426 42109 3472
rect 22109 3397 42109 3426
rect 42341 3472 62341 3501
rect 42341 3426 42354 3472
rect 62328 3426 62341 3472
rect 42341 3397 62341 3426
rect 1877 3248 21877 3277
rect 1877 3202 1890 3248
rect 21864 3202 21877 3248
rect 1877 3173 21877 3202
rect 22109 3248 42109 3277
rect 22109 3202 22122 3248
rect 42096 3202 42109 3248
rect 22109 3173 42109 3202
rect 42341 3248 62341 3277
rect 42341 3202 42354 3248
rect 62328 3202 62341 3248
rect 42341 3173 62341 3202
rect 1877 3024 21877 3053
rect 1877 2978 1890 3024
rect 21864 2978 21877 3024
rect 1877 2949 21877 2978
rect 22109 3024 42109 3053
rect 22109 2978 22122 3024
rect 42096 2978 42109 3024
rect 22109 2949 42109 2978
rect 42341 3024 62341 3053
rect 42341 2978 42354 3024
rect 62328 2978 62341 3024
rect 42341 2949 62341 2978
rect 1877 2800 21877 2829
rect 1877 2754 1890 2800
rect 21864 2754 21877 2800
rect 1877 2741 21877 2754
rect 22109 2800 42109 2829
rect 22109 2754 22122 2800
rect 42096 2754 42109 2800
rect 22109 2741 42109 2754
rect 42341 2800 62341 2829
rect 42341 2754 42354 2800
rect 62328 2754 62341 2800
rect 42341 2741 62341 2754
rect 629 2259 717 2272
rect 629 285 642 2259
rect 688 285 717 2259
rect 629 272 717 285
rect 837 2259 925 2272
rect 837 285 866 2259
rect 912 285 925 2259
rect 837 272 925 285
rect 1141 2259 1229 2272
rect 1141 285 1154 2259
rect 1200 285 1229 2259
rect 1141 272 1229 285
rect 1349 2259 1437 2272
rect 1349 285 1378 2259
rect 1424 285 1437 2259
rect 1349 272 1437 285
rect 1877 2112 21877 2125
rect 1877 2066 1890 2112
rect 21864 2066 21877 2112
rect 1877 2037 21877 2066
rect 22109 2112 42109 2125
rect 22109 2066 22122 2112
rect 42096 2066 42109 2112
rect 22109 2037 42109 2066
rect 42341 2112 62341 2125
rect 42341 2066 42354 2112
rect 62328 2066 62341 2112
rect 42341 2037 62341 2066
rect 1877 1888 21877 1917
rect 1877 1842 1890 1888
rect 21864 1842 21877 1888
rect 1877 1813 21877 1842
rect 22109 1888 42109 1917
rect 22109 1842 22122 1888
rect 42096 1842 42109 1888
rect 22109 1813 42109 1842
rect 42341 1888 62341 1917
rect 42341 1842 42354 1888
rect 62328 1842 62341 1888
rect 42341 1813 62341 1842
rect 1877 1664 21877 1693
rect 1877 1618 1890 1664
rect 21864 1618 21877 1664
rect 1877 1589 21877 1618
rect 22109 1664 42109 1693
rect 22109 1618 22122 1664
rect 42096 1618 42109 1664
rect 22109 1589 42109 1618
rect 42341 1664 62341 1693
rect 42341 1618 42354 1664
rect 62328 1618 62341 1664
rect 42341 1589 62341 1618
rect 1877 1440 21877 1469
rect 1877 1394 1890 1440
rect 21864 1394 21877 1440
rect 1877 1365 21877 1394
rect 22109 1440 42109 1469
rect 22109 1394 22122 1440
rect 42096 1394 42109 1440
rect 22109 1365 42109 1394
rect 42341 1440 62341 1469
rect 42341 1394 42354 1440
rect 62328 1394 62341 1440
rect 42341 1365 62341 1394
rect 1877 1216 21877 1245
rect 1877 1170 1890 1216
rect 21864 1170 21877 1216
rect 1877 1141 21877 1170
rect 22109 1216 42109 1245
rect 22109 1170 22122 1216
rect 42096 1170 42109 1216
rect 22109 1141 42109 1170
rect 42341 1216 62341 1245
rect 42341 1170 42354 1216
rect 62328 1170 62341 1216
rect 42341 1141 62341 1170
rect 1877 992 21877 1021
rect 1877 946 1890 992
rect 21864 946 21877 992
rect 1877 917 21877 946
rect 22109 992 42109 1021
rect 22109 946 22122 992
rect 42096 946 42109 992
rect 22109 917 42109 946
rect 42341 992 62341 1021
rect 42341 946 42354 992
rect 62328 946 62341 992
rect 42341 917 62341 946
rect 1877 768 21877 797
rect 1877 722 1890 768
rect 21864 722 21877 768
rect 1877 693 21877 722
rect 22109 768 42109 797
rect 22109 722 22122 768
rect 42096 722 42109 768
rect 22109 693 42109 722
rect 42341 768 62341 797
rect 42341 722 42354 768
rect 62328 722 62341 768
rect 42341 693 62341 722
rect 1877 544 21877 573
rect 1877 498 1890 544
rect 21864 498 21877 544
rect 1877 485 21877 498
rect 22109 544 42109 573
rect 22109 498 22122 544
rect 42096 498 42109 544
rect 22109 485 42109 498
rect 42341 544 62341 573
rect 42341 498 42354 544
rect 62328 498 62341 544
rect 42341 485 62341 498
<< mvpdiff >>
rect 608 8755 696 8768
rect 608 5981 621 8755
rect 667 5981 696 8755
rect 608 5968 696 5981
rect 816 8755 904 8768
rect 816 5981 845 8755
rect 891 5981 904 8755
rect 816 5968 904 5981
rect 1120 8755 1208 8768
rect 1120 5981 1133 8755
rect 1179 5981 1208 8755
rect 1120 5968 1208 5981
rect 1328 8755 1416 8768
rect 1328 5981 1357 8755
rect 1403 5981 1416 8755
rect 1328 5968 1416 5981
rect 1880 8834 21880 8847
rect 1880 8788 1893 8834
rect 21867 8788 21880 8834
rect 1880 8759 21880 8788
rect 22112 8834 42112 8847
rect 22112 8788 22125 8834
rect 42099 8788 42112 8834
rect 22112 8759 42112 8788
rect 42344 8834 62344 8847
rect 42344 8788 42357 8834
rect 62331 8788 62344 8834
rect 42344 8759 62344 8788
rect 1880 8610 21880 8639
rect 1880 8564 1893 8610
rect 21867 8564 21880 8610
rect 1880 8535 21880 8564
rect 22112 8610 42112 8639
rect 22112 8564 22125 8610
rect 42099 8564 42112 8610
rect 22112 8535 42112 8564
rect 42344 8610 62344 8639
rect 42344 8564 42357 8610
rect 62331 8564 62344 8610
rect 42344 8535 62344 8564
rect 1880 8386 21880 8415
rect 1880 8340 1893 8386
rect 21867 8340 21880 8386
rect 1880 8311 21880 8340
rect 22112 8386 42112 8415
rect 22112 8340 22125 8386
rect 42099 8340 42112 8386
rect 22112 8311 42112 8340
rect 42344 8386 62344 8415
rect 42344 8340 42357 8386
rect 62331 8340 62344 8386
rect 42344 8311 62344 8340
rect 1880 8162 21880 8191
rect 1880 8116 1893 8162
rect 21867 8116 21880 8162
rect 1880 8087 21880 8116
rect 22112 8162 42112 8191
rect 22112 8116 22125 8162
rect 42099 8116 42112 8162
rect 22112 8087 42112 8116
rect 42344 8162 62344 8191
rect 42344 8116 42357 8162
rect 62331 8116 62344 8162
rect 42344 8087 62344 8116
rect 1880 7938 21880 7967
rect 1880 7892 1893 7938
rect 21867 7892 21880 7938
rect 1880 7863 21880 7892
rect 22112 7938 42112 7967
rect 22112 7892 22125 7938
rect 42099 7892 42112 7938
rect 22112 7863 42112 7892
rect 42344 7938 62344 7967
rect 42344 7892 42357 7938
rect 62331 7892 62344 7938
rect 42344 7863 62344 7892
rect 1880 7714 21880 7743
rect 1880 7668 1893 7714
rect 21867 7668 21880 7714
rect 1880 7639 21880 7668
rect 22112 7714 42112 7743
rect 22112 7668 22125 7714
rect 42099 7668 42112 7714
rect 22112 7639 42112 7668
rect 42344 7714 62344 7743
rect 42344 7668 42357 7714
rect 62331 7668 62344 7714
rect 42344 7639 62344 7668
rect 1880 7490 21880 7519
rect 1880 7444 1893 7490
rect 21867 7444 21880 7490
rect 1880 7415 21880 7444
rect 22112 7490 42112 7519
rect 22112 7444 22125 7490
rect 42099 7444 42112 7490
rect 22112 7415 42112 7444
rect 42344 7490 62344 7519
rect 42344 7444 42357 7490
rect 62331 7444 62344 7490
rect 42344 7415 62344 7444
rect 1880 7266 21880 7295
rect 1880 7220 1893 7266
rect 21867 7220 21880 7266
rect 1880 7207 21880 7220
rect 22112 7266 42112 7295
rect 22112 7220 22125 7266
rect 42099 7220 42112 7266
rect 22112 7207 42112 7220
rect 42344 7266 62344 7295
rect 42344 7220 42357 7266
rect 62331 7220 62344 7266
rect 42344 7207 62344 7220
rect 474 5579 562 5592
rect 474 2805 487 5579
rect 533 2805 562 5579
rect 474 2792 562 2805
rect 682 5579 770 5592
rect 682 2805 711 5579
rect 757 2805 770 5579
rect 682 2792 770 2805
rect 986 5579 1074 5592
rect 986 2805 999 5579
rect 1045 2805 1074 5579
rect 986 2792 1074 2805
rect 1194 5579 1282 5592
rect 1194 2805 1223 5579
rect 1269 2805 1282 5579
rect 1194 2792 1282 2805
rect 1880 6578 21880 6591
rect 1880 6532 1893 6578
rect 21867 6532 21880 6578
rect 1880 6503 21880 6532
rect 22112 6578 42112 6591
rect 22112 6532 22125 6578
rect 42099 6532 42112 6578
rect 22112 6503 42112 6532
rect 42344 6578 62344 6591
rect 42344 6532 42357 6578
rect 62331 6532 62344 6578
rect 42344 6503 62344 6532
rect 1880 6354 21880 6383
rect 1880 6308 1893 6354
rect 21867 6308 21880 6354
rect 1880 6279 21880 6308
rect 22112 6354 42112 6383
rect 22112 6308 22125 6354
rect 42099 6308 42112 6354
rect 22112 6279 42112 6308
rect 42344 6354 62344 6383
rect 42344 6308 42357 6354
rect 62331 6308 62344 6354
rect 42344 6279 62344 6308
rect 1880 6130 21880 6159
rect 1880 6084 1893 6130
rect 21867 6084 21880 6130
rect 1880 6055 21880 6084
rect 22112 6130 42112 6159
rect 22112 6084 22125 6130
rect 42099 6084 42112 6130
rect 22112 6055 42112 6084
rect 42344 6130 62344 6159
rect 42344 6084 42357 6130
rect 62331 6084 62344 6130
rect 42344 6055 62344 6084
rect 1880 5906 21880 5935
rect 1880 5860 1893 5906
rect 21867 5860 21880 5906
rect 1880 5831 21880 5860
rect 22112 5906 42112 5935
rect 22112 5860 22125 5906
rect 42099 5860 42112 5906
rect 22112 5831 42112 5860
rect 42344 5906 62344 5935
rect 42344 5860 42357 5906
rect 62331 5860 62344 5906
rect 42344 5831 62344 5860
rect 1880 5682 21880 5711
rect 1880 5636 1893 5682
rect 21867 5636 21880 5682
rect 1880 5607 21880 5636
rect 22112 5682 42112 5711
rect 22112 5636 22125 5682
rect 42099 5636 42112 5682
rect 22112 5607 42112 5636
rect 42344 5682 62344 5711
rect 42344 5636 42357 5682
rect 62331 5636 62344 5682
rect 42344 5607 62344 5636
rect 1880 5458 21880 5487
rect 1880 5412 1893 5458
rect 21867 5412 21880 5458
rect 1880 5383 21880 5412
rect 22112 5458 42112 5487
rect 22112 5412 22125 5458
rect 42099 5412 42112 5458
rect 22112 5383 42112 5412
rect 42344 5458 62344 5487
rect 42344 5412 42357 5458
rect 62331 5412 62344 5458
rect 42344 5383 62344 5412
rect 1880 5234 21880 5263
rect 1880 5188 1893 5234
rect 21867 5188 21880 5234
rect 1880 5159 21880 5188
rect 22112 5234 42112 5263
rect 22112 5188 22125 5234
rect 42099 5188 42112 5234
rect 22112 5159 42112 5188
rect 42344 5234 62344 5263
rect 42344 5188 42357 5234
rect 62331 5188 62344 5234
rect 42344 5159 62344 5188
rect 1880 5010 21880 5039
rect 1880 4964 1893 5010
rect 21867 4964 21880 5010
rect 1880 4951 21880 4964
rect 22112 5010 42112 5039
rect 22112 4964 22125 5010
rect 42099 4964 42112 5010
rect 22112 4951 42112 4964
rect 42344 5010 62344 5039
rect 42344 4964 42357 5010
rect 62331 4964 62344 5010
rect 42344 4951 62344 4964
<< mvndiffc >>
rect 1890 4322 21864 4368
rect 22122 4322 42096 4368
rect 42354 4322 62328 4368
rect 1890 4098 21864 4144
rect 22122 4098 42096 4144
rect 42354 4098 62328 4144
rect 1890 3874 21864 3920
rect 22122 3874 42096 3920
rect 42354 3874 62328 3920
rect 1890 3650 21864 3696
rect 22122 3650 42096 3696
rect 42354 3650 62328 3696
rect 1890 3426 21864 3472
rect 22122 3426 42096 3472
rect 42354 3426 62328 3472
rect 1890 3202 21864 3248
rect 22122 3202 42096 3248
rect 42354 3202 62328 3248
rect 1890 2978 21864 3024
rect 22122 2978 42096 3024
rect 42354 2978 62328 3024
rect 1890 2754 21864 2800
rect 22122 2754 42096 2800
rect 42354 2754 62328 2800
rect 642 285 688 2259
rect 866 285 912 2259
rect 1154 285 1200 2259
rect 1378 285 1424 2259
rect 1890 2066 21864 2112
rect 22122 2066 42096 2112
rect 42354 2066 62328 2112
rect 1890 1842 21864 1888
rect 22122 1842 42096 1888
rect 42354 1842 62328 1888
rect 1890 1618 21864 1664
rect 22122 1618 42096 1664
rect 42354 1618 62328 1664
rect 1890 1394 21864 1440
rect 22122 1394 42096 1440
rect 42354 1394 62328 1440
rect 1890 1170 21864 1216
rect 22122 1170 42096 1216
rect 42354 1170 62328 1216
rect 1890 946 21864 992
rect 22122 946 42096 992
rect 42354 946 62328 992
rect 1890 722 21864 768
rect 22122 722 42096 768
rect 42354 722 62328 768
rect 1890 498 21864 544
rect 22122 498 42096 544
rect 42354 498 62328 544
<< mvpdiffc >>
rect 621 5981 667 8755
rect 845 5981 891 8755
rect 1133 5981 1179 8755
rect 1357 5981 1403 8755
rect 1893 8788 21867 8834
rect 22125 8788 42099 8834
rect 42357 8788 62331 8834
rect 1893 8564 21867 8610
rect 22125 8564 42099 8610
rect 42357 8564 62331 8610
rect 1893 8340 21867 8386
rect 22125 8340 42099 8386
rect 42357 8340 62331 8386
rect 1893 8116 21867 8162
rect 22125 8116 42099 8162
rect 42357 8116 62331 8162
rect 1893 7892 21867 7938
rect 22125 7892 42099 7938
rect 42357 7892 62331 7938
rect 1893 7668 21867 7714
rect 22125 7668 42099 7714
rect 42357 7668 62331 7714
rect 1893 7444 21867 7490
rect 22125 7444 42099 7490
rect 42357 7444 62331 7490
rect 1893 7220 21867 7266
rect 22125 7220 42099 7266
rect 42357 7220 62331 7266
rect 487 2805 533 5579
rect 711 2805 757 5579
rect 999 2805 1045 5579
rect 1223 2805 1269 5579
rect 1893 6532 21867 6578
rect 22125 6532 42099 6578
rect 42357 6532 62331 6578
rect 1893 6308 21867 6354
rect 22125 6308 42099 6354
rect 42357 6308 62331 6354
rect 1893 6084 21867 6130
rect 22125 6084 42099 6130
rect 42357 6084 62331 6130
rect 1893 5860 21867 5906
rect 22125 5860 42099 5906
rect 42357 5860 62331 5906
rect 1893 5636 21867 5682
rect 22125 5636 42099 5682
rect 42357 5636 62331 5682
rect 1893 5412 21867 5458
rect 22125 5412 42099 5458
rect 42357 5412 62331 5458
rect 1893 5188 21867 5234
rect 22125 5188 42099 5234
rect 42357 5188 62331 5234
rect 1893 4964 21867 5010
rect 22125 4964 42099 5010
rect 42357 4964 62331 5010
<< mvpsubdiff >>
rect 1653 4512 62565 4525
rect 1653 4466 1769 4512
rect 62449 4466 62565 4512
rect 1653 4453 62565 4466
rect 1653 2669 1725 4453
rect 62493 2669 62565 4453
rect 1653 2656 62565 2669
rect 1653 2610 1769 2656
rect 62449 2610 62565 2656
rect 1653 2597 62565 2610
rect 485 2424 1581 2496
rect 485 2380 557 2424
rect 485 164 498 2380
rect 544 164 557 2380
rect 997 2380 1069 2424
rect 485 120 557 164
rect 997 164 1010 2380
rect 1056 164 1069 2380
rect 1509 2380 1581 2424
rect 997 120 1069 164
rect 1509 164 1522 2380
rect 1568 164 1581 2380
rect 1653 2256 62565 2269
rect 1653 2210 1769 2256
rect 62449 2210 62565 2256
rect 1653 2197 62565 2210
rect 1653 413 1725 2197
rect 62493 413 62565 2197
rect 1653 400 62565 413
rect 1653 354 1769 400
rect 62449 354 62565 400
rect 1653 341 62565 354
rect 1509 120 1581 164
rect 485 48 1581 120
<< mvnsubdiff >>
rect 464 8920 1560 8992
rect 464 8876 536 8920
rect 464 5860 477 8876
rect 523 5860 536 8876
rect 976 8876 1048 8920
rect 464 5816 536 5860
rect 976 5860 989 8876
rect 1035 5860 1048 8876
rect 1488 8876 1560 8920
rect 976 5816 1048 5860
rect 1488 5860 1501 8876
rect 1547 5860 1560 8876
rect 1656 8978 62568 8991
rect 1656 8932 1772 8978
rect 62452 8932 62568 8978
rect 1656 8919 62568 8932
rect 1656 7135 1728 8919
rect 62496 7135 62568 8919
rect 1656 7122 62568 7135
rect 1656 7076 1772 7122
rect 62452 7076 62568 7122
rect 1656 7063 62568 7076
rect 1488 5816 1560 5860
rect 330 5744 1560 5816
rect 1656 6722 62568 6735
rect 1656 6676 1772 6722
rect 62452 6676 62568 6722
rect 1656 6663 62568 6676
rect 330 5700 402 5744
rect 330 2684 343 5700
rect 389 2684 402 5700
rect 842 5700 914 5744
rect 330 2640 402 2684
rect 842 2684 855 5700
rect 901 2684 914 5700
rect 1354 5700 1426 5744
rect 842 2640 914 2684
rect 1354 2684 1367 5700
rect 1413 2684 1426 5700
rect 1656 4879 1728 6663
rect 62496 4879 62568 6663
rect 1656 4866 62568 4879
rect 1656 4820 1772 4866
rect 62452 4820 62568 4866
rect 1656 4807 62568 4820
rect 1354 2640 1426 2684
rect 330 2568 1426 2640
<< mvpsubdiffcont >>
rect 1769 4466 62449 4512
rect 1769 2610 62449 2656
rect 498 164 544 2380
rect 1010 164 1056 2380
rect 1522 164 1568 2380
rect 1769 2210 62449 2256
rect 1769 354 62449 400
<< mvnsubdiffcont >>
rect 477 5860 523 8876
rect 989 5860 1035 8876
rect 1501 5860 1547 8876
rect 1772 8932 62452 8978
rect 1772 7076 62452 7122
rect 1772 6676 62452 6722
rect 343 2684 389 5700
rect 855 2684 901 5700
rect 1367 2684 1413 5700
rect 1772 4820 62452 4866
<< polysilicon >>
rect 696 8847 816 8860
rect 696 8801 709 8847
rect 803 8801 816 8847
rect 696 8768 816 8801
rect 696 5935 816 5968
rect 696 5889 709 5935
rect 803 5889 816 5935
rect 696 5876 816 5889
rect 1208 8847 1328 8860
rect 1208 8801 1221 8847
rect 1315 8801 1328 8847
rect 1208 8768 1328 8801
rect 1208 5935 1328 5968
rect 1208 5889 1221 5935
rect 1315 5889 1328 5935
rect 1208 5876 1328 5889
rect 1788 8746 1880 8759
rect 1788 8652 1801 8746
rect 1847 8652 1880 8746
rect 1788 8639 1880 8652
rect 21880 8742 22112 8759
rect 21880 8656 21913 8742
rect 21959 8656 22033 8742
rect 22079 8656 22112 8742
rect 21880 8639 22112 8656
rect 42112 8742 42344 8759
rect 42112 8656 42145 8742
rect 42191 8656 42265 8742
rect 42311 8656 42344 8742
rect 42112 8639 42344 8656
rect 62344 8746 62436 8759
rect 62344 8652 62377 8746
rect 62423 8652 62436 8746
rect 62344 8639 62436 8652
rect 1788 8522 1880 8535
rect 1788 8428 1801 8522
rect 1847 8428 1880 8522
rect 1788 8415 1880 8428
rect 21880 8518 22112 8535
rect 21880 8432 21913 8518
rect 21959 8432 22033 8518
rect 22079 8432 22112 8518
rect 21880 8415 22112 8432
rect 42112 8518 42344 8535
rect 42112 8432 42145 8518
rect 42191 8432 42265 8518
rect 42311 8432 42344 8518
rect 42112 8415 42344 8432
rect 62344 8522 62436 8535
rect 62344 8428 62377 8522
rect 62423 8428 62436 8522
rect 62344 8415 62436 8428
rect 1788 8298 1880 8311
rect 1788 8204 1801 8298
rect 1847 8204 1880 8298
rect 1788 8191 1880 8204
rect 21880 8294 22112 8311
rect 21880 8208 21913 8294
rect 21959 8208 22033 8294
rect 22079 8208 22112 8294
rect 21880 8191 22112 8208
rect 42112 8294 42344 8311
rect 42112 8208 42145 8294
rect 42191 8208 42265 8294
rect 42311 8208 42344 8294
rect 42112 8191 42344 8208
rect 62344 8298 62436 8311
rect 62344 8204 62377 8298
rect 62423 8204 62436 8298
rect 62344 8191 62436 8204
rect 1788 8074 1880 8087
rect 1788 7980 1801 8074
rect 1847 7980 1880 8074
rect 1788 7967 1880 7980
rect 21880 8070 22112 8087
rect 21880 7984 21913 8070
rect 21959 7984 22033 8070
rect 22079 7984 22112 8070
rect 21880 7967 22112 7984
rect 42112 8070 42344 8087
rect 42112 7984 42145 8070
rect 42191 7984 42265 8070
rect 42311 7984 42344 8070
rect 42112 7967 42344 7984
rect 62344 8074 62436 8087
rect 62344 7980 62377 8074
rect 62423 7980 62436 8074
rect 62344 7967 62436 7980
rect 1788 7850 1880 7863
rect 1788 7756 1801 7850
rect 1847 7756 1880 7850
rect 1788 7743 1880 7756
rect 21880 7846 22112 7863
rect 21880 7760 21913 7846
rect 21959 7760 22033 7846
rect 22079 7760 22112 7846
rect 21880 7743 22112 7760
rect 42112 7846 42344 7863
rect 42112 7760 42145 7846
rect 42191 7760 42265 7846
rect 42311 7760 42344 7846
rect 42112 7743 42344 7760
rect 62344 7850 62436 7863
rect 62344 7756 62377 7850
rect 62423 7756 62436 7850
rect 62344 7743 62436 7756
rect 1788 7626 1880 7639
rect 1788 7532 1801 7626
rect 1847 7532 1880 7626
rect 1788 7519 1880 7532
rect 21880 7622 22112 7639
rect 21880 7536 21913 7622
rect 21959 7536 22033 7622
rect 22079 7536 22112 7622
rect 21880 7519 22112 7536
rect 42112 7622 42344 7639
rect 42112 7536 42145 7622
rect 42191 7536 42265 7622
rect 42311 7536 42344 7622
rect 42112 7519 42344 7536
rect 62344 7626 62436 7639
rect 62344 7532 62377 7626
rect 62423 7532 62436 7626
rect 62344 7519 62436 7532
rect 1788 7402 1880 7415
rect 1788 7308 1801 7402
rect 1847 7308 1880 7402
rect 1788 7295 1880 7308
rect 21880 7398 22112 7415
rect 21880 7312 21913 7398
rect 21959 7312 22033 7398
rect 22079 7312 22112 7398
rect 21880 7295 22112 7312
rect 42112 7398 42344 7415
rect 42112 7312 42145 7398
rect 42191 7312 42265 7398
rect 42311 7312 42344 7398
rect 42112 7295 42344 7312
rect 62344 7402 62436 7415
rect 62344 7308 62377 7402
rect 62423 7308 62436 7402
rect 62344 7295 62436 7308
rect 562 5671 682 5684
rect 562 5625 575 5671
rect 669 5625 682 5671
rect 562 5592 682 5625
rect 562 2759 682 2792
rect 562 2713 575 2759
rect 669 2713 682 2759
rect 562 2700 682 2713
rect 1074 5671 1194 5684
rect 1074 5625 1087 5671
rect 1181 5625 1194 5671
rect 1074 5592 1194 5625
rect 1074 2759 1194 2792
rect 1074 2713 1087 2759
rect 1181 2713 1194 2759
rect 1074 2700 1194 2713
rect 1788 6490 1880 6503
rect 1788 6396 1801 6490
rect 1847 6396 1880 6490
rect 1788 6383 1880 6396
rect 21880 6486 22112 6503
rect 21880 6400 21913 6486
rect 21959 6400 22033 6486
rect 22079 6400 22112 6486
rect 21880 6383 22112 6400
rect 42112 6486 42344 6503
rect 42112 6400 42145 6486
rect 42191 6400 42265 6486
rect 42311 6400 42344 6486
rect 42112 6383 42344 6400
rect 62344 6490 62436 6503
rect 62344 6396 62377 6490
rect 62423 6396 62436 6490
rect 62344 6383 62436 6396
rect 1788 6266 1880 6279
rect 1788 6172 1801 6266
rect 1847 6172 1880 6266
rect 1788 6159 1880 6172
rect 21880 6262 22112 6279
rect 21880 6176 21913 6262
rect 21959 6176 22033 6262
rect 22079 6176 22112 6262
rect 21880 6159 22112 6176
rect 42112 6262 42344 6279
rect 42112 6176 42145 6262
rect 42191 6176 42265 6262
rect 42311 6176 42344 6262
rect 42112 6159 42344 6176
rect 62344 6266 62436 6279
rect 62344 6172 62377 6266
rect 62423 6172 62436 6266
rect 62344 6159 62436 6172
rect 1788 6042 1880 6055
rect 1788 5948 1801 6042
rect 1847 5948 1880 6042
rect 1788 5935 1880 5948
rect 21880 6038 22112 6055
rect 21880 5952 21913 6038
rect 21959 5952 22033 6038
rect 22079 5952 22112 6038
rect 21880 5935 22112 5952
rect 42112 6038 42344 6055
rect 42112 5952 42145 6038
rect 42191 5952 42265 6038
rect 42311 5952 42344 6038
rect 42112 5935 42344 5952
rect 62344 6042 62436 6055
rect 62344 5948 62377 6042
rect 62423 5948 62436 6042
rect 62344 5935 62436 5948
rect 1788 5818 1880 5831
rect 1788 5724 1801 5818
rect 1847 5724 1880 5818
rect 1788 5711 1880 5724
rect 21880 5814 22112 5831
rect 21880 5728 21913 5814
rect 21959 5728 22033 5814
rect 22079 5728 22112 5814
rect 21880 5711 22112 5728
rect 42112 5814 42344 5831
rect 42112 5728 42145 5814
rect 42191 5728 42265 5814
rect 42311 5728 42344 5814
rect 42112 5711 42344 5728
rect 62344 5818 62436 5831
rect 62344 5724 62377 5818
rect 62423 5724 62436 5818
rect 62344 5711 62436 5724
rect 1788 5594 1880 5607
rect 1788 5500 1801 5594
rect 1847 5500 1880 5594
rect 1788 5487 1880 5500
rect 21880 5590 22112 5607
rect 21880 5504 21913 5590
rect 21959 5504 22033 5590
rect 22079 5504 22112 5590
rect 21880 5487 22112 5504
rect 42112 5590 42344 5607
rect 42112 5504 42145 5590
rect 42191 5504 42265 5590
rect 42311 5504 42344 5590
rect 42112 5487 42344 5504
rect 62344 5594 62436 5607
rect 62344 5500 62377 5594
rect 62423 5500 62436 5594
rect 62344 5487 62436 5500
rect 1788 5370 1880 5383
rect 1788 5276 1801 5370
rect 1847 5276 1880 5370
rect 1788 5263 1880 5276
rect 21880 5366 22112 5383
rect 21880 5280 21913 5366
rect 21959 5280 22033 5366
rect 22079 5280 22112 5366
rect 21880 5263 22112 5280
rect 42112 5366 42344 5383
rect 42112 5280 42145 5366
rect 42191 5280 42265 5366
rect 42311 5280 42344 5366
rect 42112 5263 42344 5280
rect 62344 5370 62436 5383
rect 62344 5276 62377 5370
rect 62423 5276 62436 5370
rect 62344 5263 62436 5276
rect 1788 5146 1880 5159
rect 1788 5052 1801 5146
rect 1847 5052 1880 5146
rect 1788 5039 1880 5052
rect 21880 5142 22112 5159
rect 21880 5056 21913 5142
rect 21959 5056 22033 5142
rect 22079 5056 22112 5142
rect 21880 5039 22112 5056
rect 42112 5142 42344 5159
rect 42112 5056 42145 5142
rect 42191 5056 42265 5142
rect 42311 5056 42344 5142
rect 42112 5039 42344 5056
rect 62344 5146 62436 5159
rect 62344 5052 62377 5146
rect 62423 5052 62436 5146
rect 62344 5039 62436 5052
rect 1785 4280 1877 4293
rect 1785 4186 1798 4280
rect 1844 4186 1877 4280
rect 1785 4173 1877 4186
rect 21877 4276 22109 4293
rect 21877 4190 21910 4276
rect 21956 4190 22030 4276
rect 22076 4190 22109 4276
rect 21877 4173 22109 4190
rect 42109 4276 42341 4293
rect 42109 4190 42142 4276
rect 42188 4190 42262 4276
rect 42308 4190 42341 4276
rect 42109 4173 42341 4190
rect 62341 4280 62433 4293
rect 62341 4186 62374 4280
rect 62420 4186 62433 4280
rect 62341 4173 62433 4186
rect 1785 4056 1877 4069
rect 1785 3962 1798 4056
rect 1844 3962 1877 4056
rect 1785 3949 1877 3962
rect 21877 4052 22109 4069
rect 21877 3966 21910 4052
rect 21956 3966 22030 4052
rect 22076 3966 22109 4052
rect 21877 3949 22109 3966
rect 42109 4052 42341 4069
rect 42109 3966 42142 4052
rect 42188 3966 42262 4052
rect 42308 3966 42341 4052
rect 42109 3949 42341 3966
rect 62341 4056 62433 4069
rect 62341 3962 62374 4056
rect 62420 3962 62433 4056
rect 62341 3949 62433 3962
rect 1785 3832 1877 3845
rect 1785 3738 1798 3832
rect 1844 3738 1877 3832
rect 1785 3725 1877 3738
rect 21877 3828 22109 3845
rect 21877 3742 21910 3828
rect 21956 3742 22030 3828
rect 22076 3742 22109 3828
rect 21877 3725 22109 3742
rect 42109 3828 42341 3845
rect 42109 3742 42142 3828
rect 42188 3742 42262 3828
rect 42308 3742 42341 3828
rect 42109 3725 42341 3742
rect 62341 3832 62433 3845
rect 62341 3738 62374 3832
rect 62420 3738 62433 3832
rect 62341 3725 62433 3738
rect 1785 3608 1877 3621
rect 1785 3514 1798 3608
rect 1844 3514 1877 3608
rect 1785 3501 1877 3514
rect 21877 3604 22109 3621
rect 21877 3518 21910 3604
rect 21956 3518 22030 3604
rect 22076 3518 22109 3604
rect 21877 3501 22109 3518
rect 42109 3604 42341 3621
rect 42109 3518 42142 3604
rect 42188 3518 42262 3604
rect 42308 3518 42341 3604
rect 42109 3501 42341 3518
rect 62341 3608 62433 3621
rect 62341 3514 62374 3608
rect 62420 3514 62433 3608
rect 62341 3501 62433 3514
rect 1785 3384 1877 3397
rect 1785 3290 1798 3384
rect 1844 3290 1877 3384
rect 1785 3277 1877 3290
rect 21877 3380 22109 3397
rect 21877 3294 21910 3380
rect 21956 3294 22030 3380
rect 22076 3294 22109 3380
rect 21877 3277 22109 3294
rect 42109 3380 42341 3397
rect 42109 3294 42142 3380
rect 42188 3294 42262 3380
rect 42308 3294 42341 3380
rect 42109 3277 42341 3294
rect 62341 3384 62433 3397
rect 62341 3290 62374 3384
rect 62420 3290 62433 3384
rect 62341 3277 62433 3290
rect 1785 3160 1877 3173
rect 1785 3066 1798 3160
rect 1844 3066 1877 3160
rect 1785 3053 1877 3066
rect 21877 3156 22109 3173
rect 21877 3070 21910 3156
rect 21956 3070 22030 3156
rect 22076 3070 22109 3156
rect 21877 3053 22109 3070
rect 42109 3156 42341 3173
rect 42109 3070 42142 3156
rect 42188 3070 42262 3156
rect 42308 3070 42341 3156
rect 42109 3053 42341 3070
rect 62341 3160 62433 3173
rect 62341 3066 62374 3160
rect 62420 3066 62433 3160
rect 62341 3053 62433 3066
rect 1785 2936 1877 2949
rect 1785 2842 1798 2936
rect 1844 2842 1877 2936
rect 1785 2829 1877 2842
rect 21877 2932 22109 2949
rect 21877 2846 21910 2932
rect 21956 2846 22030 2932
rect 22076 2846 22109 2932
rect 21877 2829 22109 2846
rect 42109 2932 42341 2949
rect 42109 2846 42142 2932
rect 42188 2846 42262 2932
rect 42308 2846 42341 2932
rect 42109 2829 42341 2846
rect 62341 2936 62433 2949
rect 62341 2842 62374 2936
rect 62420 2842 62433 2936
rect 62341 2829 62433 2842
rect 717 2351 837 2364
rect 717 2305 730 2351
rect 824 2305 837 2351
rect 717 2272 837 2305
rect 717 239 837 272
rect 717 193 730 239
rect 824 193 837 239
rect 717 180 837 193
rect 1229 2351 1349 2364
rect 1229 2305 1242 2351
rect 1336 2305 1349 2351
rect 1229 2272 1349 2305
rect 1229 239 1349 272
rect 1229 193 1242 239
rect 1336 193 1349 239
rect 1229 180 1349 193
rect 1785 2024 1877 2037
rect 1785 1930 1798 2024
rect 1844 1930 1877 2024
rect 1785 1917 1877 1930
rect 21877 2020 22109 2037
rect 21877 1934 21910 2020
rect 21956 1934 22030 2020
rect 22076 1934 22109 2020
rect 21877 1917 22109 1934
rect 42109 2020 42341 2037
rect 42109 1934 42142 2020
rect 42188 1934 42262 2020
rect 42308 1934 42341 2020
rect 42109 1917 42341 1934
rect 62341 2024 62433 2037
rect 62341 1930 62374 2024
rect 62420 1930 62433 2024
rect 62341 1917 62433 1930
rect 1785 1800 1877 1813
rect 1785 1706 1798 1800
rect 1844 1706 1877 1800
rect 1785 1693 1877 1706
rect 21877 1796 22109 1813
rect 21877 1710 21910 1796
rect 21956 1710 22030 1796
rect 22076 1710 22109 1796
rect 21877 1693 22109 1710
rect 42109 1796 42341 1813
rect 42109 1710 42142 1796
rect 42188 1710 42262 1796
rect 42308 1710 42341 1796
rect 42109 1693 42341 1710
rect 62341 1800 62433 1813
rect 62341 1706 62374 1800
rect 62420 1706 62433 1800
rect 62341 1693 62433 1706
rect 1785 1576 1877 1589
rect 1785 1482 1798 1576
rect 1844 1482 1877 1576
rect 1785 1469 1877 1482
rect 21877 1572 22109 1589
rect 21877 1486 21910 1572
rect 21956 1486 22030 1572
rect 22076 1486 22109 1572
rect 21877 1469 22109 1486
rect 42109 1572 42341 1589
rect 42109 1486 42142 1572
rect 42188 1486 42262 1572
rect 42308 1486 42341 1572
rect 42109 1469 42341 1486
rect 62341 1576 62433 1589
rect 62341 1482 62374 1576
rect 62420 1482 62433 1576
rect 62341 1469 62433 1482
rect 1785 1352 1877 1365
rect 1785 1258 1798 1352
rect 1844 1258 1877 1352
rect 1785 1245 1877 1258
rect 21877 1348 22109 1365
rect 21877 1262 21910 1348
rect 21956 1262 22030 1348
rect 22076 1262 22109 1348
rect 21877 1245 22109 1262
rect 42109 1348 42341 1365
rect 42109 1262 42142 1348
rect 42188 1262 42262 1348
rect 42308 1262 42341 1348
rect 42109 1245 42341 1262
rect 62341 1352 62433 1365
rect 62341 1258 62374 1352
rect 62420 1258 62433 1352
rect 62341 1245 62433 1258
rect 1785 1128 1877 1141
rect 1785 1034 1798 1128
rect 1844 1034 1877 1128
rect 1785 1021 1877 1034
rect 21877 1124 22109 1141
rect 21877 1038 21910 1124
rect 21956 1038 22030 1124
rect 22076 1038 22109 1124
rect 21877 1021 22109 1038
rect 42109 1124 42341 1141
rect 42109 1038 42142 1124
rect 42188 1038 42262 1124
rect 42308 1038 42341 1124
rect 42109 1021 42341 1038
rect 62341 1128 62433 1141
rect 62341 1034 62374 1128
rect 62420 1034 62433 1128
rect 62341 1021 62433 1034
rect 1785 904 1877 917
rect 1785 810 1798 904
rect 1844 810 1877 904
rect 1785 797 1877 810
rect 21877 900 22109 917
rect 21877 814 21910 900
rect 21956 814 22030 900
rect 22076 814 22109 900
rect 21877 797 22109 814
rect 42109 900 42341 917
rect 42109 814 42142 900
rect 42188 814 42262 900
rect 42308 814 42341 900
rect 42109 797 42341 814
rect 62341 904 62433 917
rect 62341 810 62374 904
rect 62420 810 62433 904
rect 62341 797 62433 810
rect 1785 680 1877 693
rect 1785 586 1798 680
rect 1844 586 1877 680
rect 1785 573 1877 586
rect 21877 676 22109 693
rect 21877 590 21910 676
rect 21956 590 22030 676
rect 22076 590 22109 676
rect 21877 573 22109 590
rect 42109 676 42341 693
rect 42109 590 42142 676
rect 42188 590 42262 676
rect 42308 590 42341 676
rect 42109 573 42341 590
rect 62341 680 62433 693
rect 62341 586 62374 680
rect 62420 586 62433 680
rect 62341 573 62433 586
<< polycontact >>
rect 709 8801 803 8847
rect 709 5889 803 5935
rect 1221 8801 1315 8847
rect 1221 5889 1315 5935
rect 1801 8652 1847 8746
rect 21913 8656 21959 8742
rect 22033 8656 22079 8742
rect 42145 8656 42191 8742
rect 42265 8656 42311 8742
rect 62377 8652 62423 8746
rect 1801 8428 1847 8522
rect 21913 8432 21959 8518
rect 22033 8432 22079 8518
rect 42145 8432 42191 8518
rect 42265 8432 42311 8518
rect 62377 8428 62423 8522
rect 1801 8204 1847 8298
rect 21913 8208 21959 8294
rect 22033 8208 22079 8294
rect 42145 8208 42191 8294
rect 42265 8208 42311 8294
rect 62377 8204 62423 8298
rect 1801 7980 1847 8074
rect 21913 7984 21959 8070
rect 22033 7984 22079 8070
rect 42145 7984 42191 8070
rect 42265 7984 42311 8070
rect 62377 7980 62423 8074
rect 1801 7756 1847 7850
rect 21913 7760 21959 7846
rect 22033 7760 22079 7846
rect 42145 7760 42191 7846
rect 42265 7760 42311 7846
rect 62377 7756 62423 7850
rect 1801 7532 1847 7626
rect 21913 7536 21959 7622
rect 22033 7536 22079 7622
rect 42145 7536 42191 7622
rect 42265 7536 42311 7622
rect 62377 7532 62423 7626
rect 1801 7308 1847 7402
rect 21913 7312 21959 7398
rect 22033 7312 22079 7398
rect 42145 7312 42191 7398
rect 42265 7312 42311 7398
rect 62377 7308 62423 7402
rect 575 5625 669 5671
rect 575 2713 669 2759
rect 1087 5625 1181 5671
rect 1087 2713 1181 2759
rect 1801 6396 1847 6490
rect 21913 6400 21959 6486
rect 22033 6400 22079 6486
rect 42145 6400 42191 6486
rect 42265 6400 42311 6486
rect 62377 6396 62423 6490
rect 1801 6172 1847 6266
rect 21913 6176 21959 6262
rect 22033 6176 22079 6262
rect 42145 6176 42191 6262
rect 42265 6176 42311 6262
rect 62377 6172 62423 6266
rect 1801 5948 1847 6042
rect 21913 5952 21959 6038
rect 22033 5952 22079 6038
rect 42145 5952 42191 6038
rect 42265 5952 42311 6038
rect 62377 5948 62423 6042
rect 1801 5724 1847 5818
rect 21913 5728 21959 5814
rect 22033 5728 22079 5814
rect 42145 5728 42191 5814
rect 42265 5728 42311 5814
rect 62377 5724 62423 5818
rect 1801 5500 1847 5594
rect 21913 5504 21959 5590
rect 22033 5504 22079 5590
rect 42145 5504 42191 5590
rect 42265 5504 42311 5590
rect 62377 5500 62423 5594
rect 1801 5276 1847 5370
rect 21913 5280 21959 5366
rect 22033 5280 22079 5366
rect 42145 5280 42191 5366
rect 42265 5280 42311 5366
rect 62377 5276 62423 5370
rect 1801 5052 1847 5146
rect 21913 5056 21959 5142
rect 22033 5056 22079 5142
rect 42145 5056 42191 5142
rect 42265 5056 42311 5142
rect 62377 5052 62423 5146
rect 1798 4186 1844 4280
rect 21910 4190 21956 4276
rect 22030 4190 22076 4276
rect 42142 4190 42188 4276
rect 42262 4190 42308 4276
rect 62374 4186 62420 4280
rect 1798 3962 1844 4056
rect 21910 3966 21956 4052
rect 22030 3966 22076 4052
rect 42142 3966 42188 4052
rect 42262 3966 42308 4052
rect 62374 3962 62420 4056
rect 1798 3738 1844 3832
rect 21910 3742 21956 3828
rect 22030 3742 22076 3828
rect 42142 3742 42188 3828
rect 42262 3742 42308 3828
rect 62374 3738 62420 3832
rect 1798 3514 1844 3608
rect 21910 3518 21956 3604
rect 22030 3518 22076 3604
rect 42142 3518 42188 3604
rect 42262 3518 42308 3604
rect 62374 3514 62420 3608
rect 1798 3290 1844 3384
rect 21910 3294 21956 3380
rect 22030 3294 22076 3380
rect 42142 3294 42188 3380
rect 42262 3294 42308 3380
rect 62374 3290 62420 3384
rect 1798 3066 1844 3160
rect 21910 3070 21956 3156
rect 22030 3070 22076 3156
rect 42142 3070 42188 3156
rect 42262 3070 42308 3156
rect 62374 3066 62420 3160
rect 1798 2842 1844 2936
rect 21910 2846 21956 2932
rect 22030 2846 22076 2932
rect 42142 2846 42188 2932
rect 42262 2846 42308 2932
rect 62374 2842 62420 2936
rect 730 2305 824 2351
rect 730 193 824 239
rect 1242 2305 1336 2351
rect 1242 193 1336 239
rect 1798 1930 1844 2024
rect 21910 1934 21956 2020
rect 22030 1934 22076 2020
rect 42142 1934 42188 2020
rect 42262 1934 42308 2020
rect 62374 1930 62420 2024
rect 1798 1706 1844 1800
rect 21910 1710 21956 1796
rect 22030 1710 22076 1796
rect 42142 1710 42188 1796
rect 42262 1710 42308 1796
rect 62374 1706 62420 1800
rect 1798 1482 1844 1576
rect 21910 1486 21956 1572
rect 22030 1486 22076 1572
rect 42142 1486 42188 1572
rect 42262 1486 42308 1572
rect 62374 1482 62420 1576
rect 1798 1258 1844 1352
rect 21910 1262 21956 1348
rect 22030 1262 22076 1348
rect 42142 1262 42188 1348
rect 42262 1262 42308 1348
rect 62374 1258 62420 1352
rect 1798 1034 1844 1128
rect 21910 1038 21956 1124
rect 22030 1038 22076 1124
rect 42142 1038 42188 1124
rect 42262 1038 42308 1124
rect 62374 1034 62420 1128
rect 1798 810 1844 904
rect 21910 814 21956 900
rect 22030 814 22076 900
rect 42142 814 42188 900
rect 42262 814 42308 900
rect 62374 810 62420 904
rect 1798 586 1844 680
rect 21910 590 21956 676
rect 22030 590 22076 676
rect 42142 590 42188 676
rect 42262 590 42308 676
rect 62374 586 62420 680
<< metal1 >>
rect 298 8978 62677 9333
rect 298 8933 1772 8978
rect 298 8876 523 8933
rect 298 5860 477 8876
rect 989 8876 1035 8933
rect 698 8856 814 8857
rect 698 8847 710 8856
rect 802 8847 814 8856
rect 698 8801 709 8847
rect 803 8801 814 8847
rect 621 8755 667 8766
rect 603 6103 615 8230
rect 621 5970 667 5981
rect 845 8755 989 8766
rect 891 5981 989 8755
rect 845 5970 989 5981
rect 698 5889 709 5935
rect 803 5889 814 5935
rect 698 5883 710 5889
rect 802 5883 814 5889
rect 698 5879 814 5883
rect 298 5803 523 5860
rect 1501 8932 1772 8933
rect 62452 8932 62677 8978
rect 1501 8876 62677 8932
rect 1210 8856 1326 8857
rect 1210 8847 1222 8856
rect 1314 8847 1326 8856
rect 1210 8801 1221 8847
rect 1315 8801 1326 8847
rect 1115 8755 1179 8766
rect 1115 8754 1133 8755
rect 1115 5982 1127 8754
rect 1115 5981 1133 5982
rect 1115 5970 1179 5981
rect 1357 8755 1501 8766
rect 1403 5981 1501 8755
rect 1357 5970 1501 5981
rect 1210 5889 1221 5935
rect 1315 5889 1326 5935
rect 1210 5883 1222 5889
rect 1314 5883 1326 5889
rect 1210 5879 1326 5883
rect 989 5803 1035 5860
rect 1547 8852 62677 8876
rect 1547 8840 32646 8852
rect 1547 8834 1902 8840
rect 21826 8834 32646 8840
rect 42012 8834 62677 8852
rect 1547 7122 1715 8834
rect 1882 8788 1893 8834
rect 21867 8788 22125 8834
rect 42099 8788 42357 8834
rect 62331 8788 62342 8834
rect 1761 8746 1847 8757
rect 1761 8739 1801 8746
rect 62377 8746 62463 8757
rect 1761 7309 1764 8739
rect 21902 8656 21913 8742
rect 22079 8656 22090 8742
rect 42134 8656 42145 8742
rect 42311 8656 42322 8742
rect 62423 8739 62463 8746
rect 1816 8641 1847 8652
rect 62377 8641 62407 8652
rect 22165 8616 31539 8628
rect 42416 8616 62262 8628
rect 1882 8564 1893 8610
rect 21867 8564 22125 8610
rect 42099 8564 42357 8610
rect 62331 8564 62342 8610
rect 62396 8533 62407 8641
rect 1816 8522 1847 8533
rect 62377 8522 62407 8533
rect 21902 8432 21913 8518
rect 22079 8432 22090 8518
rect 42134 8432 42145 8518
rect 42311 8432 42322 8518
rect 1816 8417 1847 8428
rect 62377 8417 62407 8428
rect 32646 8404 42012 8416
rect 1904 8392 21828 8404
rect 1882 8340 1893 8386
rect 21867 8340 22125 8386
rect 42099 8340 42357 8386
rect 62331 8340 62342 8386
rect 62396 8309 62407 8417
rect 1816 8298 1847 8309
rect 62377 8298 62407 8309
rect 21902 8208 21913 8294
rect 22079 8208 22090 8294
rect 42134 8208 42145 8294
rect 42311 8208 42322 8294
rect 1816 8193 1847 8204
rect 62377 8193 62407 8204
rect 22168 8168 31542 8180
rect 42417 8168 62263 8180
rect 1882 8116 1893 8162
rect 21867 8116 22125 8162
rect 42099 8116 42357 8162
rect 62331 8116 62342 8162
rect 62396 8085 62407 8193
rect 1816 8074 1847 8085
rect 62377 8074 62407 8085
rect 21902 7984 21913 8070
rect 22079 7984 22090 8070
rect 42134 7984 42145 8070
rect 42311 7984 42322 8070
rect 1816 7969 1847 7980
rect 62377 7969 62407 7980
rect 32643 7956 42009 7968
rect 1908 7944 21832 7956
rect 1882 7892 1893 7938
rect 21867 7892 22125 7938
rect 42099 7892 42357 7938
rect 62331 7892 62342 7938
rect 62396 7861 62407 7969
rect 1816 7850 1847 7861
rect 62377 7850 62407 7861
rect 21902 7760 21913 7846
rect 22079 7760 22090 7846
rect 42134 7760 42145 7846
rect 42311 7760 42322 7846
rect 1816 7745 1847 7756
rect 62377 7745 62407 7756
rect 22166 7720 31540 7732
rect 42418 7720 62264 7732
rect 1882 7668 1893 7714
rect 21867 7668 22125 7714
rect 42099 7668 42357 7714
rect 62331 7668 62342 7714
rect 62396 7637 62407 7745
rect 1816 7626 1847 7637
rect 62377 7626 62407 7637
rect 21902 7536 21913 7622
rect 22079 7536 22090 7622
rect 42134 7536 42145 7622
rect 42311 7536 42322 7622
rect 1816 7521 1847 7532
rect 62377 7521 62407 7532
rect 32639 7508 42005 7520
rect 1908 7496 21832 7508
rect 1882 7444 1893 7490
rect 21867 7444 22125 7490
rect 42099 7444 42357 7490
rect 62331 7444 62342 7490
rect 62396 7413 62407 7521
rect 1816 7402 1847 7413
rect 62377 7402 62407 7413
rect 21902 7312 21913 7398
rect 22079 7312 22090 7398
rect 42134 7312 42145 7398
rect 42311 7312 42322 7398
rect 1761 7308 1801 7309
rect 1761 7297 1847 7308
rect 62459 7309 62463 8739
rect 62423 7308 62463 7309
rect 62377 7297 62463 7308
rect 22168 7272 31542 7284
rect 42413 7272 62259 7284
rect 1882 7220 1893 7266
rect 21867 7220 22125 7266
rect 42099 7220 42357 7266
rect 62331 7220 62342 7266
rect 62509 7122 62677 8834
rect 1547 7076 1772 7122
rect 62452 7076 62677 7122
rect 1547 6722 1910 7076
rect 21834 6722 32640 7076
rect 42006 6722 62677 7076
rect 1547 6676 1772 6722
rect 62452 6676 62677 6722
rect 1547 6578 1910 6676
rect 21834 6584 32640 6676
rect 21835 6578 32640 6584
rect 42006 6578 62677 6676
rect 1547 5860 1715 6578
rect 1882 6532 1893 6578
rect 21867 6532 22125 6578
rect 42099 6532 42357 6578
rect 62331 6532 62342 6578
rect 1501 5803 1715 5860
rect 298 5757 1715 5803
rect 298 5700 389 5757
rect 298 2684 343 5700
rect 855 5700 901 5757
rect 564 5671 680 5681
rect 564 5625 575 5671
rect 669 5625 680 5671
rect 582 5600 653 5625
rect 487 5579 533 5590
rect 437 4199 487 4211
rect 437 2800 449 4199
rect 501 2800 533 2805
rect 437 2794 533 2800
rect 582 5042 589 5600
rect 641 5042 653 5600
rect 582 2759 653 5042
rect 711 5579 757 5590
rect 763 3061 775 5385
rect 711 2794 757 2805
rect 564 2713 575 2759
rect 669 2713 680 2759
rect 564 2703 680 2713
rect 298 2627 389 2684
rect 1367 5700 1715 5757
rect 1076 5671 1192 5681
rect 1076 5625 1087 5671
rect 1181 5625 1192 5671
rect 999 5579 1045 5590
rect 980 3056 992 5380
rect 1110 2991 1157 5625
rect 999 2794 1045 2805
rect 1093 2759 1105 2991
rect 1223 5579 1269 5590
rect 1275 3114 1287 5386
rect 1223 2794 1269 2805
rect 1076 2713 1087 2759
rect 1181 2713 1192 2759
rect 1076 2703 1088 2713
rect 1180 2703 1192 2713
rect 855 2627 901 2684
rect 1413 4866 1715 5700
rect 1761 6490 1847 6501
rect 1761 6489 1801 6490
rect 1761 5053 1764 6489
rect 62377 6490 62463 6501
rect 62423 6489 62463 6490
rect 21902 6400 21913 6486
rect 22079 6400 22090 6486
rect 42134 6400 42145 6486
rect 42311 6400 42322 6486
rect 1816 6385 1847 6396
rect 62377 6385 62407 6396
rect 22164 6360 31538 6372
rect 42421 6360 62267 6372
rect 1882 6308 1893 6354
rect 21867 6308 22125 6354
rect 42099 6308 42357 6354
rect 62331 6308 62342 6354
rect 62396 6277 62407 6385
rect 1816 6266 1847 6277
rect 62377 6266 62407 6277
rect 21902 6176 21913 6262
rect 22079 6176 22090 6262
rect 42134 6176 42145 6262
rect 42311 6176 42322 6262
rect 1816 6161 1847 6172
rect 62377 6161 62407 6172
rect 32645 6148 42011 6160
rect 1904 6136 21828 6148
rect 1882 6084 1893 6130
rect 21867 6084 22125 6130
rect 42099 6084 42357 6130
rect 62331 6084 62342 6130
rect 62396 6053 62407 6161
rect 1816 6042 1847 6053
rect 62377 6042 62407 6053
rect 21902 5952 21913 6038
rect 22079 5952 22090 6038
rect 42134 5952 42145 6038
rect 42311 5952 42322 6038
rect 1816 5937 1847 5948
rect 62377 5937 62407 5948
rect 22165 5912 31539 5924
rect 42426 5912 62272 5924
rect 1882 5860 1893 5906
rect 21867 5860 22125 5906
rect 42099 5860 42357 5906
rect 62331 5860 62342 5906
rect 62396 5829 62407 5937
rect 1816 5818 1847 5829
rect 62377 5818 62407 5829
rect 21902 5728 21913 5814
rect 22079 5728 22090 5814
rect 42134 5728 42145 5814
rect 42311 5728 42322 5814
rect 1816 5713 1847 5724
rect 62377 5713 62407 5724
rect 32646 5700 42012 5712
rect 1910 5688 21834 5700
rect 1882 5636 1893 5682
rect 21867 5636 22125 5682
rect 42099 5636 42357 5682
rect 62331 5636 62342 5682
rect 62396 5605 62407 5713
rect 1816 5594 1847 5605
rect 62377 5594 62407 5605
rect 21902 5504 21913 5590
rect 22079 5504 22090 5590
rect 42134 5504 42145 5590
rect 42311 5504 42322 5590
rect 1816 5489 1847 5500
rect 62377 5489 62407 5500
rect 22163 5464 31537 5476
rect 42428 5464 62274 5476
rect 1882 5412 1893 5458
rect 21867 5412 22125 5458
rect 42099 5412 42357 5458
rect 62331 5412 62342 5458
rect 62396 5381 62407 5489
rect 1816 5370 1847 5381
rect 62377 5370 62407 5381
rect 21902 5280 21913 5366
rect 22079 5280 22090 5366
rect 42134 5280 42145 5366
rect 42311 5280 42322 5366
rect 1816 5265 1847 5276
rect 62377 5265 62407 5276
rect 32644 5252 42010 5264
rect 1903 5240 21827 5252
rect 1882 5188 1893 5234
rect 21867 5188 22125 5234
rect 42099 5188 42357 5234
rect 62331 5188 62342 5234
rect 62396 5157 62407 5265
rect 1816 5146 1847 5157
rect 62377 5146 62407 5157
rect 21902 5056 21913 5142
rect 22079 5056 22090 5142
rect 42134 5056 42145 5142
rect 42311 5056 42322 5142
rect 1761 5052 1801 5053
rect 1761 5041 1847 5052
rect 62459 5053 62463 6489
rect 62423 5052 62463 5053
rect 62377 5041 62463 5052
rect 22165 5016 31539 5028
rect 42419 5016 62265 5028
rect 1882 4964 1893 5010
rect 21867 4964 22125 5010
rect 42099 4964 42357 5010
rect 62331 4964 62342 5010
rect 62509 4866 62677 6578
rect 1413 4820 1772 4866
rect 62452 4820 62677 4866
rect 1413 4675 62677 4820
rect 1367 2627 1413 2684
rect 298 2581 1413 2627
rect 1544 4628 2545 4629
rect 1544 4512 62677 4628
rect 1544 4466 1769 4512
rect 62449 4466 62677 4512
rect 1544 4387 62677 4466
rect 1544 4374 32662 4387
rect 1544 4368 1901 4374
rect 21823 4368 32662 4374
rect 42028 4368 62677 4387
rect 1544 2656 1712 4368
rect 1879 4322 1890 4368
rect 21864 4322 22122 4368
rect 42096 4322 42354 4368
rect 62328 4322 62339 4368
rect 1758 4280 1844 4291
rect 1758 4279 1798 4280
rect 62374 4280 62460 4291
rect 62420 4279 62460 4280
rect 21899 4190 21910 4276
rect 22076 4190 22087 4276
rect 42131 4190 42142 4276
rect 42308 4190 42319 4276
rect 1810 4175 1844 4186
rect 62374 4175 62408 4186
rect 22171 4150 31545 4162
rect 42417 4150 62263 4162
rect 1879 4098 1890 4144
rect 21864 4098 22122 4144
rect 42096 4098 42354 4144
rect 62328 4098 62339 4144
rect 1810 4056 1844 4067
rect 62374 4056 62408 4067
rect 21899 3966 21910 4052
rect 22076 3966 22087 4052
rect 42131 3966 42142 4052
rect 42308 3966 42319 4052
rect 1810 3951 1844 3962
rect 62374 3951 62408 3962
rect 32664 3939 42030 3951
rect 1907 3926 21831 3938
rect 21823 3920 21831 3926
rect 1879 3874 1890 3920
rect 21864 3874 22122 3920
rect 42096 3874 42354 3920
rect 62328 3874 62339 3920
rect 1810 3832 1844 3843
rect 62374 3832 62408 3843
rect 21899 3742 21910 3828
rect 22076 3742 22087 3828
rect 42131 3742 42142 3828
rect 42308 3742 42319 3828
rect 1810 3727 1844 3738
rect 62374 3727 62408 3738
rect 22170 3702 31544 3714
rect 42421 3702 62267 3714
rect 1879 3650 1890 3696
rect 21864 3650 22122 3696
rect 42096 3650 42354 3696
rect 62328 3650 62339 3696
rect 1810 3608 1844 3619
rect 62374 3608 62408 3619
rect 21899 3518 21910 3604
rect 22076 3518 22087 3604
rect 42131 3518 42142 3604
rect 42308 3518 42319 3604
rect 1810 3503 1844 3514
rect 62374 3503 62408 3514
rect 32664 3491 42030 3503
rect 1909 3478 21833 3490
rect 21823 3472 21833 3478
rect 1879 3426 1890 3472
rect 21864 3426 22122 3472
rect 42096 3426 42354 3472
rect 62328 3426 62339 3472
rect 1810 3384 1844 3395
rect 62374 3384 62408 3395
rect 21899 3294 21910 3380
rect 22076 3294 22087 3380
rect 42131 3294 42142 3380
rect 42308 3294 42319 3380
rect 1810 3279 1844 3290
rect 62374 3279 62408 3290
rect 22167 3254 31541 3266
rect 42423 3254 62269 3266
rect 1879 3202 1890 3248
rect 21864 3202 22122 3248
rect 42096 3202 42354 3248
rect 62328 3202 62339 3248
rect 1810 3160 1844 3171
rect 62374 3160 62408 3171
rect 21899 3070 21910 3156
rect 22076 3070 22087 3156
rect 42131 3070 42142 3156
rect 42308 3070 42319 3156
rect 1810 3055 1844 3066
rect 62374 3055 62408 3066
rect 32663 3043 42029 3055
rect 1905 3030 21829 3042
rect 21823 3024 21829 3030
rect 1879 2978 1890 3024
rect 21864 2978 22122 3024
rect 42096 2978 42354 3024
rect 62328 2978 62339 3024
rect 1810 2936 1844 2947
rect 62374 2936 62408 2947
rect 21899 2846 21910 2932
rect 22076 2846 22087 2932
rect 42131 2846 42142 2932
rect 42308 2846 42319 2932
rect 1758 2842 1798 2843
rect 1758 2831 1844 2842
rect 62420 2842 62460 2843
rect 62374 2831 62460 2842
rect 22168 2807 31542 2819
rect 42418 2806 62264 2818
rect 1879 2754 1890 2800
rect 21864 2754 22122 2800
rect 42096 2754 42354 2800
rect 62328 2754 62339 2800
rect 62506 2656 62677 4368
rect 1544 2610 1769 2656
rect 62449 2610 62677 2656
rect 1544 2483 1899 2610
rect 297 2437 1899 2483
rect 297 2380 544 2437
rect 297 164 498 2380
rect 1010 2380 1056 2437
rect 719 2351 835 2366
rect 719 2305 730 2351
rect 824 2305 835 2351
rect 719 2270 801 2305
rect 642 2259 801 2270
rect 688 2258 801 2259
rect 699 1301 801 2258
rect 688 285 801 1301
rect 642 274 801 285
rect 866 2259 1010 2270
rect 912 285 1010 2259
rect 866 274 1010 285
rect 719 239 801 274
rect 719 193 730 239
rect 824 193 835 239
rect 719 178 835 193
rect 297 107 544 164
rect 1522 2380 1899 2437
rect 1231 2351 1347 2366
rect 1231 2305 1242 2351
rect 1336 2305 1347 2351
rect 1056 2259 1200 2270
rect 1056 285 1154 2259
rect 1267 1392 1314 2305
rect 1251 1380 1314 1392
rect 1303 882 1314 1380
rect 1251 870 1314 882
rect 1056 274 1200 285
rect 1267 239 1314 870
rect 1378 2259 1424 2270
rect 1430 449 1442 2120
rect 1378 274 1424 285
rect 1231 193 1242 239
rect 1336 193 1347 239
rect 1231 178 1347 193
rect 1010 107 1056 164
rect 1568 2256 1899 2380
rect 21823 2256 32659 2610
rect 42025 2256 62677 2610
rect 1568 2210 1769 2256
rect 62449 2210 62677 2256
rect 1568 2112 1899 2210
rect 21823 2112 32659 2210
rect 42025 2131 62677 2210
rect 42026 2112 62677 2131
rect 1568 400 1712 2112
rect 1879 2066 1890 2112
rect 21864 2066 22122 2112
rect 42096 2066 42354 2112
rect 62328 2066 62339 2112
rect 1758 2024 1844 2035
rect 1758 2023 1798 2024
rect 62374 2024 62460 2035
rect 62420 2023 62460 2024
rect 21899 1934 21910 2020
rect 22076 1934 22087 2020
rect 42131 1934 42142 2020
rect 42308 1934 42319 2020
rect 1810 1919 1844 1930
rect 62374 1919 62408 1930
rect 22170 1894 31544 1906
rect 42416 1894 62262 1906
rect 1879 1842 1890 1888
rect 21864 1842 22122 1888
rect 42096 1842 42354 1888
rect 62328 1842 62339 1888
rect 1810 1800 1844 1811
rect 62374 1800 62408 1811
rect 21899 1710 21910 1796
rect 22076 1710 22087 1796
rect 42131 1710 42142 1796
rect 42308 1710 42319 1796
rect 1810 1695 1844 1706
rect 62374 1695 62408 1706
rect 32665 1683 42031 1695
rect 1903 1670 21827 1682
rect 21823 1664 21827 1670
rect 1879 1618 1890 1664
rect 21864 1618 22122 1664
rect 42096 1618 42354 1664
rect 62328 1618 62339 1664
rect 1810 1576 1844 1587
rect 62374 1576 62408 1587
rect 21899 1486 21910 1572
rect 22076 1486 22087 1572
rect 42131 1486 42142 1572
rect 42308 1486 42319 1572
rect 1810 1471 1844 1482
rect 62374 1471 62408 1482
rect 22171 1446 31545 1458
rect 42417 1446 62263 1458
rect 1879 1394 1890 1440
rect 21864 1394 22122 1440
rect 42096 1394 42354 1440
rect 62328 1394 62339 1440
rect 1810 1352 1844 1363
rect 62374 1352 62408 1363
rect 21899 1262 21910 1348
rect 22076 1262 22087 1348
rect 42131 1262 42142 1348
rect 42308 1262 42319 1348
rect 1810 1247 1844 1258
rect 62374 1247 62408 1258
rect 32675 1235 42041 1247
rect 1903 1222 21827 1234
rect 21823 1216 21827 1222
rect 1879 1170 1890 1216
rect 21864 1170 22122 1216
rect 42096 1170 42354 1216
rect 62328 1170 62339 1216
rect 1810 1128 1844 1139
rect 62374 1128 62408 1139
rect 21899 1038 21910 1124
rect 22076 1038 22087 1124
rect 42131 1038 42142 1124
rect 42308 1038 42319 1124
rect 1810 1023 1844 1034
rect 62374 1023 62408 1034
rect 22167 998 31541 1010
rect 42422 998 62268 1010
rect 1879 946 1890 992
rect 21864 946 22122 992
rect 42096 946 42354 992
rect 62328 946 62339 992
rect 1810 904 1844 915
rect 62374 904 62408 915
rect 21899 814 21910 900
rect 22076 814 22087 900
rect 42131 814 42142 900
rect 42308 814 42319 900
rect 1810 799 1844 810
rect 62374 799 62408 810
rect 32658 787 42024 799
rect 1891 774 21815 786
rect 1879 722 1890 768
rect 21864 722 22122 768
rect 42096 722 42354 768
rect 62328 722 62339 768
rect 1810 680 1844 691
rect 62374 680 62408 691
rect 21899 590 21910 676
rect 22076 590 22087 676
rect 42131 590 42142 676
rect 42308 590 42319 676
rect 1758 586 1798 587
rect 1758 575 1844 586
rect 62420 586 62460 587
rect 62374 575 62460 586
rect 22164 550 31538 562
rect 42413 550 62259 562
rect 1879 498 1890 544
rect 21864 498 22122 544
rect 42096 498 42354 544
rect 62328 498 62339 544
rect 62506 400 62677 2112
rect 1568 354 1769 400
rect 62449 354 62677 400
rect 1568 164 62677 354
rect 1522 107 62677 164
rect 297 1 62677 107
rect 498 0 62677 1
<< via1 >>
rect 710 8847 802 8856
rect 710 8804 802 8847
rect 615 6103 621 8230
rect 621 6103 667 8230
rect 710 5889 802 5935
rect 710 5883 802 5889
rect 1222 8847 1314 8856
rect 1222 8804 1314 8847
rect 1127 5982 1133 8754
rect 1133 5982 1179 8754
rect 1222 5889 1314 5935
rect 1222 5883 1314 5889
rect 1902 8834 21826 8840
rect 32646 8834 42012 8852
rect 1902 8788 21826 8834
rect 32646 8788 42012 8834
rect 1764 8652 1801 8739
rect 1801 8652 1816 8739
rect 21914 8656 21959 8742
rect 21959 8656 22033 8742
rect 22033 8656 22078 8742
rect 42146 8656 42191 8742
rect 42191 8656 42265 8742
rect 42265 8656 42310 8742
rect 1764 8522 1816 8652
rect 62407 8652 62423 8739
rect 62423 8652 62459 8739
rect 22165 8610 31539 8616
rect 42416 8610 62262 8616
rect 22165 8564 31539 8610
rect 42416 8564 62262 8610
rect 1764 8428 1801 8522
rect 1801 8428 1816 8522
rect 62407 8522 62459 8652
rect 21914 8432 21959 8518
rect 21959 8432 22033 8518
rect 22033 8432 22078 8518
rect 42146 8432 42191 8518
rect 42191 8432 42265 8518
rect 42265 8432 42310 8518
rect 1764 8298 1816 8428
rect 62407 8428 62423 8522
rect 62423 8428 62459 8522
rect 1904 8386 21828 8392
rect 32646 8386 42012 8404
rect 1904 8340 21828 8386
rect 32646 8340 42012 8386
rect 1764 8204 1801 8298
rect 1801 8204 1816 8298
rect 62407 8298 62459 8428
rect 21914 8208 21959 8294
rect 21959 8208 22033 8294
rect 22033 8208 22078 8294
rect 42146 8208 42191 8294
rect 42191 8208 42265 8294
rect 42265 8208 42310 8294
rect 1764 8074 1816 8204
rect 62407 8204 62423 8298
rect 62423 8204 62459 8298
rect 22168 8162 31542 8168
rect 42417 8162 62263 8168
rect 22168 8116 31542 8162
rect 42417 8116 62263 8162
rect 1764 7980 1801 8074
rect 1801 7980 1816 8074
rect 62407 8074 62459 8204
rect 21914 7984 21959 8070
rect 21959 7984 22033 8070
rect 22033 7984 22078 8070
rect 42146 7984 42191 8070
rect 42191 7984 42265 8070
rect 42265 7984 42310 8070
rect 1764 7850 1816 7980
rect 62407 7980 62423 8074
rect 62423 7980 62459 8074
rect 1908 7938 21832 7944
rect 32643 7938 42009 7956
rect 1908 7892 21832 7938
rect 32643 7892 42009 7938
rect 1764 7756 1801 7850
rect 1801 7756 1816 7850
rect 62407 7850 62459 7980
rect 21914 7760 21959 7846
rect 21959 7760 22033 7846
rect 22033 7760 22078 7846
rect 42146 7760 42191 7846
rect 42191 7760 42265 7846
rect 42265 7760 42310 7846
rect 1764 7626 1816 7756
rect 62407 7756 62423 7850
rect 62423 7756 62459 7850
rect 22166 7714 31540 7720
rect 42418 7714 62264 7720
rect 22166 7668 31540 7714
rect 42418 7668 62264 7714
rect 1764 7532 1801 7626
rect 1801 7532 1816 7626
rect 62407 7626 62459 7756
rect 21914 7536 21959 7622
rect 21959 7536 22033 7622
rect 22033 7536 22078 7622
rect 42146 7536 42191 7622
rect 42191 7536 42265 7622
rect 42265 7536 42310 7622
rect 1764 7402 1816 7532
rect 62407 7532 62423 7626
rect 62423 7532 62459 7626
rect 1908 7490 21832 7496
rect 32639 7490 42005 7508
rect 1908 7444 21832 7490
rect 32639 7444 42005 7490
rect 1764 7309 1801 7402
rect 1801 7309 1816 7402
rect 62407 7402 62459 7532
rect 21914 7312 21959 7398
rect 21959 7312 22033 7398
rect 22033 7312 22078 7398
rect 42146 7312 42191 7398
rect 42191 7312 42265 7398
rect 42265 7312 42310 7398
rect 62407 7309 62423 7402
rect 62423 7309 62459 7402
rect 22168 7266 31542 7272
rect 42413 7266 62259 7272
rect 22168 7220 31542 7266
rect 42413 7220 62259 7266
rect 1910 7076 21834 7115
rect 32640 7076 42006 7116
rect 1910 6722 21834 7076
rect 32640 6722 42006 7076
rect 1910 6676 21834 6722
rect 32640 6676 42006 6722
rect 1910 6584 21834 6676
rect 1910 6578 21835 6584
rect 32640 6578 42006 6676
rect 1910 6532 21835 6578
rect 32640 6532 42006 6578
rect 449 2805 487 4199
rect 487 2805 501 4199
rect 449 2800 501 2805
rect 589 5042 641 5600
rect 711 3061 757 5385
rect 757 3061 763 5385
rect 992 3056 999 5380
rect 999 3056 1044 5380
rect 1105 2759 1157 2991
rect 1223 3114 1269 5386
rect 1269 3114 1275 5386
rect 1088 2713 1180 2759
rect 1088 2703 1180 2713
rect 1764 6396 1801 6489
rect 1801 6396 1816 6489
rect 21914 6400 21959 6486
rect 21959 6400 22033 6486
rect 22033 6400 22078 6486
rect 42146 6400 42191 6486
rect 42191 6400 42265 6486
rect 42265 6400 42310 6486
rect 1764 6266 1816 6396
rect 62407 6396 62423 6489
rect 62423 6396 62459 6489
rect 22164 6354 31538 6360
rect 42421 6354 62267 6360
rect 22164 6308 31538 6354
rect 42421 6308 62267 6354
rect 1764 6172 1801 6266
rect 1801 6172 1816 6266
rect 62407 6266 62459 6396
rect 21914 6176 21959 6262
rect 21959 6176 22033 6262
rect 22033 6176 22078 6262
rect 42146 6176 42191 6262
rect 42191 6176 42265 6262
rect 42265 6176 42310 6262
rect 1764 6042 1816 6172
rect 62407 6172 62423 6266
rect 62423 6172 62459 6266
rect 1904 6130 21828 6136
rect 32645 6130 42011 6148
rect 1904 6084 21828 6130
rect 32645 6084 42011 6130
rect 1764 5948 1801 6042
rect 1801 5948 1816 6042
rect 62407 6042 62459 6172
rect 21914 5952 21959 6038
rect 21959 5952 22033 6038
rect 22033 5952 22078 6038
rect 42146 5952 42191 6038
rect 42191 5952 42265 6038
rect 42265 5952 42310 6038
rect 1764 5818 1816 5948
rect 62407 5948 62423 6042
rect 62423 5948 62459 6042
rect 22165 5906 31539 5912
rect 42426 5906 62272 5912
rect 22165 5860 31539 5906
rect 42426 5860 62272 5906
rect 1764 5724 1801 5818
rect 1801 5724 1816 5818
rect 62407 5818 62459 5948
rect 21914 5728 21959 5814
rect 21959 5728 22033 5814
rect 22033 5728 22078 5814
rect 42146 5728 42191 5814
rect 42191 5728 42265 5814
rect 42265 5728 42310 5814
rect 1764 5594 1816 5724
rect 62407 5724 62423 5818
rect 62423 5724 62459 5818
rect 1910 5682 21834 5688
rect 32646 5682 42012 5700
rect 1910 5636 21834 5682
rect 32646 5636 42012 5682
rect 1764 5500 1801 5594
rect 1801 5500 1816 5594
rect 62407 5594 62459 5724
rect 21914 5504 21959 5590
rect 21959 5504 22033 5590
rect 22033 5504 22078 5590
rect 42146 5504 42191 5590
rect 42191 5504 42265 5590
rect 42265 5504 42310 5590
rect 1764 5370 1816 5500
rect 62407 5500 62423 5594
rect 62423 5500 62459 5594
rect 22163 5458 31537 5464
rect 42428 5458 62274 5464
rect 22163 5412 31537 5458
rect 42428 5412 62274 5458
rect 1764 5276 1801 5370
rect 1801 5276 1816 5370
rect 62407 5370 62459 5500
rect 21914 5280 21959 5366
rect 21959 5280 22033 5366
rect 22033 5280 22078 5366
rect 42146 5280 42191 5366
rect 42191 5280 42265 5366
rect 42265 5280 42310 5366
rect 1764 5146 1816 5276
rect 62407 5276 62423 5370
rect 62423 5276 62459 5370
rect 1903 5234 21827 5240
rect 32644 5234 42010 5252
rect 1903 5188 21827 5234
rect 32644 5188 42010 5234
rect 1764 5053 1801 5146
rect 1801 5053 1816 5146
rect 62407 5146 62459 5276
rect 21914 5056 21959 5142
rect 21959 5056 22033 5142
rect 22033 5056 22078 5142
rect 42146 5056 42191 5142
rect 42191 5056 42265 5142
rect 42265 5056 42310 5142
rect 62407 5053 62423 5146
rect 62423 5053 62459 5146
rect 22165 5010 31539 5016
rect 42419 5010 62265 5016
rect 22165 4964 31539 5010
rect 42419 4964 62265 5010
rect 1901 4368 21823 4374
rect 32662 4368 42028 4387
rect 1901 4322 21823 4368
rect 32662 4322 42028 4368
rect 1758 4186 1798 4279
rect 1798 4186 1810 4279
rect 21911 4190 21956 4276
rect 21956 4190 22030 4276
rect 22030 4190 22075 4276
rect 42143 4190 42188 4276
rect 42188 4190 42262 4276
rect 42262 4190 42307 4276
rect 1758 4056 1810 4186
rect 62408 4186 62420 4279
rect 62420 4186 62460 4279
rect 22171 4144 31545 4150
rect 42417 4144 62263 4150
rect 22171 4098 31545 4144
rect 42417 4098 62263 4144
rect 1758 3962 1798 4056
rect 1798 3962 1810 4056
rect 62408 4056 62460 4186
rect 21911 3966 21956 4052
rect 21956 3966 22030 4052
rect 22030 3966 22075 4052
rect 42143 3966 42188 4052
rect 42188 3966 42262 4052
rect 42262 3966 42307 4052
rect 1758 3832 1810 3962
rect 62408 3962 62420 4056
rect 62420 3962 62460 4056
rect 1907 3920 21823 3926
rect 32664 3920 42030 3939
rect 1907 3874 21823 3920
rect 32664 3874 42030 3920
rect 1758 3738 1798 3832
rect 1798 3738 1810 3832
rect 62408 3832 62460 3962
rect 21911 3742 21956 3828
rect 21956 3742 22030 3828
rect 22030 3742 22075 3828
rect 42143 3742 42188 3828
rect 42188 3742 42262 3828
rect 42262 3742 42307 3828
rect 1758 3608 1810 3738
rect 62408 3738 62420 3832
rect 62420 3738 62460 3832
rect 22170 3696 31544 3702
rect 42421 3696 62267 3702
rect 22170 3650 31544 3696
rect 42421 3650 62267 3696
rect 1758 3514 1798 3608
rect 1798 3514 1810 3608
rect 62408 3608 62460 3738
rect 21911 3518 21956 3604
rect 21956 3518 22030 3604
rect 22030 3518 22075 3604
rect 42143 3518 42188 3604
rect 42188 3518 42262 3604
rect 42262 3518 42307 3604
rect 1758 3384 1810 3514
rect 62408 3514 62420 3608
rect 62420 3514 62460 3608
rect 1909 3472 21823 3478
rect 32664 3472 42030 3491
rect 1909 3426 21823 3472
rect 32664 3426 42030 3472
rect 1758 3290 1798 3384
rect 1798 3290 1810 3384
rect 62408 3384 62460 3514
rect 21911 3294 21956 3380
rect 21956 3294 22030 3380
rect 22030 3294 22075 3380
rect 42143 3294 42188 3380
rect 42188 3294 42262 3380
rect 42262 3294 42307 3380
rect 1758 3160 1810 3290
rect 62408 3290 62420 3384
rect 62420 3290 62460 3384
rect 22167 3248 31541 3254
rect 42423 3248 62269 3254
rect 22167 3202 31541 3248
rect 42423 3202 62269 3248
rect 1758 3066 1798 3160
rect 1798 3066 1810 3160
rect 62408 3160 62460 3290
rect 21911 3070 21956 3156
rect 21956 3070 22030 3156
rect 22030 3070 22075 3156
rect 42143 3070 42188 3156
rect 42188 3070 42262 3156
rect 42262 3070 42307 3156
rect 1758 2936 1810 3066
rect 62408 3066 62420 3160
rect 62420 3066 62460 3160
rect 1905 3024 21823 3030
rect 32663 3024 42029 3043
rect 1905 2978 21823 3024
rect 32663 2978 42029 3024
rect 1758 2843 1798 2936
rect 1798 2843 1810 2936
rect 62408 2936 62460 3066
rect 21911 2846 21956 2932
rect 21956 2846 22030 2932
rect 22030 2846 22075 2932
rect 42143 2846 42188 2932
rect 42188 2846 42262 2932
rect 42262 2846 42307 2932
rect 62408 2843 62420 2936
rect 62420 2843 62460 2936
rect 22168 2800 31542 2807
rect 42418 2800 62264 2806
rect 22168 2755 31542 2800
rect 42418 2754 62264 2800
rect 1899 2610 21823 2649
rect 32659 2610 42025 2650
rect 647 1301 688 2258
rect 688 1301 699 2258
rect 1251 882 1303 1380
rect 1378 449 1424 2120
rect 1424 449 1430 2120
rect 1899 2256 21823 2610
rect 32659 2256 42025 2610
rect 1899 2210 21823 2256
rect 32659 2210 42025 2256
rect 1899 2112 21823 2210
rect 32659 2131 42025 2210
rect 32659 2112 42026 2131
rect 1899 2066 21823 2112
rect 32659 2066 42026 2112
rect 1758 1930 1798 2023
rect 1798 1930 1810 2023
rect 21911 1934 21956 2020
rect 21956 1934 22030 2020
rect 22030 1934 22075 2020
rect 42143 1934 42188 2020
rect 42188 1934 42262 2020
rect 42262 1934 42307 2020
rect 1758 1800 1810 1930
rect 62408 1930 62420 2023
rect 62420 1930 62460 2023
rect 22170 1888 31544 1894
rect 42416 1888 62262 1894
rect 22170 1842 31544 1888
rect 42416 1842 62262 1888
rect 1758 1706 1798 1800
rect 1798 1706 1810 1800
rect 62408 1800 62460 1930
rect 21911 1710 21956 1796
rect 21956 1710 22030 1796
rect 22030 1710 22075 1796
rect 42143 1710 42188 1796
rect 42188 1710 42262 1796
rect 42262 1710 42307 1796
rect 1758 1576 1810 1706
rect 62408 1706 62420 1800
rect 62420 1706 62460 1800
rect 1903 1664 21823 1670
rect 32665 1664 42031 1683
rect 1903 1618 21823 1664
rect 32665 1618 42031 1664
rect 1758 1482 1798 1576
rect 1798 1482 1810 1576
rect 62408 1576 62460 1706
rect 21911 1486 21956 1572
rect 21956 1486 22030 1572
rect 22030 1486 22075 1572
rect 42143 1486 42188 1572
rect 42188 1486 42262 1572
rect 42262 1486 42307 1572
rect 1758 1352 1810 1482
rect 62408 1482 62420 1576
rect 62420 1482 62460 1576
rect 22171 1440 31545 1446
rect 42417 1440 62263 1446
rect 22171 1394 31545 1440
rect 42417 1394 62263 1440
rect 1758 1258 1798 1352
rect 1798 1258 1810 1352
rect 62408 1352 62460 1482
rect 21911 1262 21956 1348
rect 21956 1262 22030 1348
rect 22030 1262 22075 1348
rect 42143 1262 42188 1348
rect 42188 1262 42262 1348
rect 42262 1262 42307 1348
rect 1758 1128 1810 1258
rect 62408 1258 62420 1352
rect 62420 1258 62460 1352
rect 1903 1216 21823 1222
rect 32675 1216 42041 1235
rect 1903 1170 21823 1216
rect 32675 1170 42041 1216
rect 1758 1034 1798 1128
rect 1798 1034 1810 1128
rect 62408 1128 62460 1258
rect 21911 1038 21956 1124
rect 21956 1038 22030 1124
rect 22030 1038 22075 1124
rect 42143 1038 42188 1124
rect 42188 1038 42262 1124
rect 42262 1038 42307 1124
rect 1758 904 1810 1034
rect 62408 1034 62420 1128
rect 62420 1034 62460 1128
rect 22167 992 31541 998
rect 42422 992 62268 998
rect 22167 946 31541 992
rect 42422 946 62268 992
rect 1758 810 1798 904
rect 1798 810 1810 904
rect 62408 904 62460 1034
rect 21911 814 21956 900
rect 21956 814 22030 900
rect 22030 814 22075 900
rect 42143 814 42188 900
rect 42188 814 42262 900
rect 42262 814 42307 900
rect 1758 680 1810 810
rect 62408 810 62420 904
rect 62420 810 62460 904
rect 1891 768 21815 774
rect 32658 768 42024 787
rect 1891 722 21815 768
rect 32658 722 42024 768
rect 1758 587 1798 680
rect 1798 587 1810 680
rect 62408 680 62460 810
rect 21911 590 21956 676
rect 21956 590 22030 676
rect 22030 590 22075 676
rect 42143 590 42188 676
rect 42188 590 42262 676
rect 42262 590 42307 676
rect 62408 587 62420 680
rect 62420 587 62460 680
rect 22164 544 31538 550
rect 42413 544 62259 550
rect 22164 498 31538 544
rect 42413 498 62259 544
<< metal2 >>
rect 1737 8947 62477 9070
rect 1737 8884 1818 8947
rect 0 8856 1818 8884
rect 0 8804 710 8856
rect 802 8804 1222 8856
rect 1314 8804 1818 8856
rect 0 8799 1818 8804
rect 697 8798 1818 8799
rect 1098 8754 1181 8798
rect 582 8230 675 8240
rect 582 6103 615 8230
rect 667 6103 675 8230
rect 582 6094 675 6103
rect 582 5799 652 6094
rect 1098 5982 1127 8754
rect 1179 5982 1181 8754
rect 708 5939 817 5947
rect 1098 5939 1181 5982
rect 1737 8739 1818 8798
rect 1737 7309 1764 8739
rect 1816 7309 1818 8739
rect 1737 6489 1818 7309
rect 1737 5939 1764 6489
rect 708 5935 1764 5939
rect 708 5883 710 5935
rect 802 5883 1222 5935
rect 1314 5883 1764 5935
rect 708 5874 1764 5883
rect 708 5871 817 5874
rect 582 5727 777 5799
rect 562 5600 648 5612
rect 562 5182 589 5600
rect 0 5097 589 5182
rect 562 5042 589 5097
rect 641 5042 648 5600
rect 562 5030 648 5042
rect 704 5397 777 5727
rect 704 5385 1056 5397
rect 0 4267 647 4352
rect 423 4199 506 4211
rect 423 2800 449 4199
rect 501 2800 506 4199
rect 562 3420 647 4267
rect 562 2993 648 3420
rect 704 3061 711 5385
rect 763 5380 1056 5385
rect 763 3061 992 5380
rect 704 3056 992 3061
rect 1044 3056 1056 5380
rect 1215 5386 1290 5394
rect 1215 3114 1223 5386
rect 1275 3995 1290 5386
rect 1737 5053 1764 5874
rect 1816 5053 1818 6489
rect 1890 8840 21838 8865
rect 1890 8788 1902 8840
rect 21826 8788 21838 8840
rect 1890 8392 21838 8788
rect 1890 8340 1904 8392
rect 21828 8340 21838 8392
rect 1890 7944 21838 8340
rect 1890 7892 1908 7944
rect 21832 7892 21838 7944
rect 1890 7496 21838 7892
rect 1890 7444 1908 7496
rect 21832 7444 21838 7496
rect 1890 7115 21838 7444
rect 1890 6532 1910 7115
rect 21834 6584 21838 7115
rect 21835 6532 21838 6584
rect 1890 6136 21838 6532
rect 1890 6084 1904 6136
rect 21828 6084 21838 6136
rect 1890 5688 21838 6084
rect 1890 5636 1910 5688
rect 21834 5636 21838 5688
rect 1890 5240 21838 5636
rect 1890 5188 1903 5240
rect 21827 5188 21838 5240
rect 1890 5164 21838 5188
rect 21902 8742 22090 8947
rect 21902 8656 21914 8742
rect 22078 8656 22090 8742
rect 32627 8852 42028 8874
rect 32627 8788 32646 8852
rect 42012 8788 42028 8852
rect 21902 8518 22090 8656
rect 21902 8432 21914 8518
rect 22078 8432 22090 8518
rect 21902 8294 22090 8432
rect 21902 8208 21914 8294
rect 22078 8208 22090 8294
rect 21902 8070 22090 8208
rect 21902 7984 21914 8070
rect 22078 7984 22090 8070
rect 21902 7846 22090 7984
rect 21902 7760 21914 7846
rect 22078 7760 22090 7846
rect 21902 7622 22090 7760
rect 21902 7536 21914 7622
rect 22078 7536 22090 7622
rect 21902 7398 22090 7536
rect 21902 7312 21914 7398
rect 22078 7312 22090 7398
rect 21902 6486 22090 7312
rect 21902 6400 21914 6486
rect 22078 6400 22090 6486
rect 21902 6262 22090 6400
rect 21902 6176 21914 6262
rect 22078 6176 22090 6262
rect 21902 6038 22090 6176
rect 21902 5952 21914 6038
rect 22078 5952 22090 6038
rect 21902 5814 22090 5952
rect 21902 5728 21914 5814
rect 22078 5728 22090 5814
rect 21902 5590 22090 5728
rect 21902 5504 21914 5590
rect 22078 5504 22090 5590
rect 21902 5366 22090 5504
rect 21902 5280 21914 5366
rect 22078 5280 22090 5366
rect 1737 5016 1818 5053
rect 21902 5142 22090 5280
rect 21902 5056 21914 5142
rect 22078 5056 22090 5142
rect 21902 5045 22090 5056
rect 22150 8616 31550 8679
rect 22150 8564 22165 8616
rect 31539 8564 31550 8616
rect 22150 8168 31550 8564
rect 22150 8116 22168 8168
rect 31542 8116 31550 8168
rect 22150 7720 31550 8116
rect 22150 7668 22166 7720
rect 31540 7668 31550 7720
rect 22150 7272 31550 7668
rect 22150 7220 22168 7272
rect 31542 7220 31550 7272
rect 22150 6360 31550 7220
rect 22150 6308 22164 6360
rect 31538 6308 31550 6360
rect 22150 5912 31550 6308
rect 22150 5860 22165 5912
rect 31539 5860 31550 5912
rect 22150 5464 31550 5860
rect 22150 5412 22163 5464
rect 31537 5412 31550 5464
rect 22150 5016 31550 5412
rect 32627 8404 42028 8788
rect 32627 8340 32646 8404
rect 42012 8340 42028 8404
rect 32627 7956 42028 8340
rect 32627 7892 32643 7956
rect 42009 7892 42028 7956
rect 32627 7508 42028 7892
rect 32627 7444 32639 7508
rect 42005 7444 42028 7508
rect 32627 7116 42028 7444
rect 32627 6532 32640 7116
rect 42006 6532 42028 7116
rect 32627 6148 42028 6532
rect 32627 6084 32645 6148
rect 42011 6084 42028 6148
rect 32627 5700 42028 6084
rect 32627 5636 32646 5700
rect 42012 5636 42028 5700
rect 32627 5252 42028 5636
rect 32627 5188 32644 5252
rect 42010 5188 42028 5252
rect 32627 5176 42028 5188
rect 42134 8742 42322 8947
rect 42134 8656 42146 8742
rect 42310 8656 42322 8742
rect 62396 8739 62477 8947
rect 42134 8518 42322 8656
rect 42134 8432 42146 8518
rect 42310 8432 42322 8518
rect 42134 8294 42322 8432
rect 42134 8208 42146 8294
rect 42310 8208 42322 8294
rect 42134 8070 42322 8208
rect 42134 7984 42146 8070
rect 42310 7984 42322 8070
rect 42134 7846 42322 7984
rect 42134 7760 42146 7846
rect 42310 7760 42322 7846
rect 42134 7622 42322 7760
rect 42134 7536 42146 7622
rect 42310 7536 42322 7622
rect 42134 7398 42322 7536
rect 42134 7312 42146 7398
rect 42310 7312 42322 7398
rect 42134 6486 42322 7312
rect 42134 6400 42146 6486
rect 42310 6400 42322 6486
rect 42134 6262 42322 6400
rect 42134 6176 42146 6262
rect 42310 6176 42322 6262
rect 42134 6038 42322 6176
rect 42134 5952 42146 6038
rect 42310 5952 42322 6038
rect 42134 5814 42322 5952
rect 42134 5728 42146 5814
rect 42310 5728 42322 5814
rect 42134 5590 42322 5728
rect 42134 5504 42146 5590
rect 42310 5504 42322 5590
rect 42134 5366 42322 5504
rect 42134 5280 42146 5366
rect 42310 5280 42322 5366
rect 42134 5142 42322 5280
rect 42134 5056 42146 5142
rect 42310 5056 42322 5142
rect 42134 5046 42322 5056
rect 42392 8616 62299 8679
rect 42392 8564 42416 8616
rect 62262 8564 62299 8616
rect 42392 8168 62299 8564
rect 42392 8116 42417 8168
rect 62263 8116 62299 8168
rect 42392 7720 62299 8116
rect 42392 7668 42418 7720
rect 62264 7668 62299 7720
rect 42392 7272 62299 7668
rect 42392 7220 42413 7272
rect 62259 7220 62299 7272
rect 42392 6360 62299 7220
rect 42392 6308 42421 6360
rect 62267 6308 62299 6360
rect 42392 5912 62299 6308
rect 42392 5860 42426 5912
rect 62272 5860 62299 5912
rect 42392 5464 62299 5860
rect 42392 5412 42428 5464
rect 62274 5412 62299 5464
rect 22150 4964 22165 5016
rect 31539 4990 31550 5016
rect 42392 5016 62299 5412
rect 42392 4990 42419 5016
rect 31539 4964 42419 4990
rect 62265 4964 62299 5016
rect 62396 7309 62407 8739
rect 62459 7309 62477 8739
rect 62396 6489 62477 7309
rect 62396 5053 62407 6489
rect 62459 5053 62477 6489
rect 62396 5008 62477 5053
rect 22150 4482 62299 4964
rect 1883 4374 21825 4408
rect 1883 4322 1901 4374
rect 21823 4322 21825 4374
rect 1691 4279 1814 4305
rect 1691 3995 1758 4279
rect 1275 3437 1758 3995
rect 1275 3114 1290 3437
rect 1215 3106 1290 3114
rect 704 3049 1056 3056
rect 562 2991 1169 2993
rect 562 2899 1105 2991
rect 423 2392 506 2800
rect 1075 2764 1105 2899
rect 1066 2759 1105 2764
rect 1157 2764 1169 2991
rect 1691 2843 1758 3437
rect 1810 2843 1814 4279
rect 1157 2759 1200 2764
rect 1066 2703 1088 2759
rect 1180 2703 1200 2759
rect 1066 2696 1200 2703
rect 423 2309 709 2392
rect 626 2258 709 2309
rect 626 1301 647 2258
rect 699 1388 709 2258
rect 1369 2120 1444 2128
rect 699 1380 1313 1388
rect 699 1301 1251 1380
rect 626 1293 1251 1301
rect 1234 882 1251 1293
rect 1303 882 1313 1380
rect 1234 874 1313 882
rect 1369 449 1378 2120
rect 1430 2078 1444 2120
rect 1691 2078 1814 2843
rect 1430 2023 1814 2078
rect 1430 1520 1758 2023
rect 1430 449 1444 1520
rect 1369 441 1444 449
rect 1691 587 1758 1520
rect 1810 587 1814 2023
rect 1883 3926 21825 4322
rect 1883 3874 1907 3926
rect 21823 3874 21825 3926
rect 1883 3478 21825 3874
rect 1883 3426 1909 3478
rect 21823 3426 21825 3478
rect 1883 3030 21825 3426
rect 1883 2978 1905 3030
rect 21823 2978 21825 3030
rect 1883 2649 21825 2978
rect 1883 2066 1899 2649
rect 21823 2066 21825 2649
rect 1883 1670 21825 2066
rect 1883 1618 1903 1670
rect 21823 1618 21825 1670
rect 1883 1222 21825 1618
rect 1883 1170 1903 1222
rect 21823 1170 21825 1222
rect 1883 774 21825 1170
rect 1883 722 1891 774
rect 21815 722 21825 774
rect 1883 707 21825 722
rect 21899 4276 22087 4311
rect 21899 4190 21911 4276
rect 22075 4190 22087 4276
rect 21899 4052 22087 4190
rect 21899 3966 21911 4052
rect 22075 3966 22087 4052
rect 21899 3828 22087 3966
rect 21899 3742 21911 3828
rect 22075 3742 22087 3828
rect 21899 3604 22087 3742
rect 21899 3518 21911 3604
rect 22075 3518 22087 3604
rect 21899 3380 22087 3518
rect 21899 3294 21911 3380
rect 22075 3294 22087 3380
rect 21899 3156 22087 3294
rect 21899 3070 21911 3156
rect 22075 3070 22087 3156
rect 21899 2932 22087 3070
rect 21899 2846 21911 2932
rect 22075 2846 22087 2932
rect 21899 2020 22087 2846
rect 21899 1934 21911 2020
rect 22075 1934 22087 2020
rect 21899 1796 22087 1934
rect 21899 1710 21911 1796
rect 22075 1710 22087 1796
rect 21899 1572 22087 1710
rect 21899 1486 21911 1572
rect 22075 1486 22087 1572
rect 21899 1348 22087 1486
rect 21899 1262 21911 1348
rect 22075 1262 22087 1348
rect 21899 1124 22087 1262
rect 21899 1038 21911 1124
rect 22075 1038 22087 1124
rect 21899 900 22087 1038
rect 21899 814 21911 900
rect 22075 814 22087 900
rect 1691 423 1814 587
rect 21899 676 22087 814
rect 21899 590 21911 676
rect 22075 590 22087 676
rect 21899 423 22087 590
rect 22150 4150 31550 4482
rect 22150 4098 22171 4150
rect 31545 4098 31550 4150
rect 22150 3702 31550 4098
rect 22150 3650 22170 3702
rect 31544 3650 31550 3702
rect 22150 3254 31550 3650
rect 22150 3202 22167 3254
rect 31541 3202 31550 3254
rect 22150 2807 31550 3202
rect 22150 2755 22168 2807
rect 31542 2755 31550 2807
rect 22150 1894 31550 2755
rect 22150 1842 22170 1894
rect 31544 1842 31550 1894
rect 22150 1446 31550 1842
rect 22150 1394 22171 1446
rect 31545 1394 31550 1446
rect 22150 998 31550 1394
rect 22150 946 22167 998
rect 31541 946 31550 998
rect 22150 550 31550 946
rect 32651 4387 42052 4396
rect 32651 4322 32662 4387
rect 42028 4322 42052 4387
rect 32651 3939 42052 4322
rect 32651 3874 32664 3939
rect 42030 3874 42052 3939
rect 32651 3491 42052 3874
rect 32651 3426 32664 3491
rect 42030 3426 42052 3491
rect 32651 3043 42052 3426
rect 32651 2978 32663 3043
rect 42029 2978 42052 3043
rect 32651 2650 42052 2978
rect 32651 2066 32659 2650
rect 42025 2131 42052 2650
rect 42026 2066 42052 2131
rect 32651 1683 42052 2066
rect 32651 1618 32665 1683
rect 42031 1618 42052 1683
rect 32651 1235 42052 1618
rect 32651 1170 32675 1235
rect 42041 1170 42052 1235
rect 32651 787 42052 1170
rect 32651 722 32658 787
rect 42024 722 42052 787
rect 32651 700 42052 722
rect 42131 4276 42319 4310
rect 42131 4190 42143 4276
rect 42307 4190 42319 4276
rect 42131 4052 42319 4190
rect 42131 3966 42143 4052
rect 42307 3966 42319 4052
rect 42131 3828 42319 3966
rect 42131 3742 42143 3828
rect 42307 3742 42319 3828
rect 42131 3604 42319 3742
rect 42131 3518 42143 3604
rect 42307 3518 42319 3604
rect 42131 3380 42319 3518
rect 42131 3294 42143 3380
rect 42307 3294 42319 3380
rect 42131 3156 42319 3294
rect 42131 3070 42143 3156
rect 42307 3070 42319 3156
rect 42131 2932 42319 3070
rect 42131 2846 42143 2932
rect 42307 2846 42319 2932
rect 42131 2020 42319 2846
rect 42131 1934 42143 2020
rect 42307 1934 42319 2020
rect 42131 1796 42319 1934
rect 42131 1710 42143 1796
rect 42307 1710 42319 1796
rect 42131 1572 42319 1710
rect 42131 1486 42143 1572
rect 42307 1486 42319 1572
rect 42131 1348 42319 1486
rect 42131 1262 42143 1348
rect 42307 1262 42319 1348
rect 42131 1124 42319 1262
rect 42131 1038 42143 1124
rect 42307 1038 42319 1124
rect 42131 900 42319 1038
rect 42131 814 42143 900
rect 42307 814 42319 900
rect 22150 498 22164 550
rect 31538 498 31550 550
rect 22150 483 31550 498
rect 42131 676 42319 814
rect 42131 590 42143 676
rect 42307 590 42319 676
rect 42131 423 42319 590
rect 42392 4150 62299 4482
rect 42392 4098 42417 4150
rect 62263 4098 62299 4150
rect 42392 3702 62299 4098
rect 42392 3650 42421 3702
rect 62267 3650 62299 3702
rect 42392 3254 62299 3650
rect 42392 3202 42423 3254
rect 62269 3202 62299 3254
rect 42392 2806 62299 3202
rect 42392 2754 42418 2806
rect 62264 2754 62299 2806
rect 42392 1894 62299 2754
rect 42392 1842 42416 1894
rect 62262 1842 62299 1894
rect 42392 1446 62299 1842
rect 42392 1394 42417 1446
rect 62263 1394 62299 1446
rect 42392 998 62299 1394
rect 42392 946 42422 998
rect 62268 946 62299 998
rect 42392 550 62299 946
rect 42392 498 42413 550
rect 62259 498 62299 550
rect 42392 483 62299 498
rect 62401 4279 62482 4305
rect 62401 2843 62408 4279
rect 62460 2843 62482 4279
rect 62401 2023 62482 2843
rect 62401 587 62408 2023
rect 62460 587 62482 2023
rect 62401 423 62482 587
rect 1691 300 62482 423
<< labels >>
flabel metal2 0 4267 286 4352 0 FreeSans 200 0 0 0 PLUS
port 1 nsew signal input
flabel metal2 0 5097 286 5182 0 FreeSans 200 0 0 0 MINUS
port 2 nsew signal input
flabel metal2 0 8799 286 8884 0 FreeSans 200 0 0 0 ADJ
port 3 nsew signal input
flabel metal1 298 9122 62677 9333 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 1613 0 62677 211 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal2 42392 483 62299 8679 0 FreeSans 200 0 0 0 OUT
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 62677 9333
<< end >>
