magic
tech gf180mcuD
magscale 1 10
timestamp 1763254865
<< pwell >>
rect 1023 10276 1331 11672
rect 2019 10276 2327 11672
rect 3015 10276 3323 11672
rect 4011 10276 4319 11672
rect 5007 10276 5315 11672
rect 6003 10276 6311 11672
rect 6999 10276 7307 11672
rect 7995 10276 8303 11672
rect 8991 10276 9299 11672
rect 9987 10276 10295 11672
rect 10982 10276 11290 11672
rect 11979 10276 12913 11672
rect 12823 9588 12913 10276
rect 335 9465 12913 9588
rect 335 9118 2266 9465
rect 335 8644 1023 9118
rect 991 6418 1055 8612
rect 2258 6386 2266 9118
rect 1023 5412 2266 6386
rect 991 3944 1050 5380
rect 335 0 1018 3912
rect 1706 2732 2266 5412
rect 2258 0 2266 2732
<< mvpsubdiff >>
rect 991 6418 1055 8612
rect 991 3944 1050 5380
<< metal1 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 11672 212 12102
rect 64759 12100 64971 12118
rect 201 11627 12909 11672
rect 201 10185 380 11627
rect 580 11423 778 11425
rect 580 11371 592 11423
rect 766 11371 778 11423
rect 580 11369 778 11371
rect 201 9679 426 10185
rect 592 10031 681 10397
rect 978 10231 1376 11627
rect 1576 11423 1774 11425
rect 1576 11371 1588 11423
rect 1762 11371 1774 11423
rect 1576 11369 1774 11371
rect 592 10022 771 10031
rect 1588 10030 1668 10443
rect 1974 10231 2372 11627
rect 2572 11423 2770 11425
rect 2572 11371 2584 11423
rect 2758 11371 2770 11423
rect 2572 11369 2770 11371
rect 2575 10030 2638 10397
rect 2970 10231 3368 11627
rect 3568 11423 3766 11425
rect 3568 11371 3580 11423
rect 3754 11371 3766 11423
rect 3568 11369 3766 11371
rect 3571 10030 3634 10397
rect 3966 10231 4364 11627
rect 4564 11423 4762 11425
rect 4564 11371 4576 11423
rect 4750 11371 4762 11423
rect 4564 11369 4762 11371
rect 4566 10030 4629 10397
rect 4962 10231 5360 11627
rect 5560 11423 5758 11425
rect 5560 11371 5572 11423
rect 5746 11371 5758 11423
rect 5560 11369 5758 11371
rect 5562 10030 5625 10397
rect 5958 10231 6356 11627
rect 6556 11423 6754 11425
rect 6556 11371 6568 11423
rect 6742 11371 6754 11423
rect 6556 11369 6754 11371
rect 6558 10030 6621 10397
rect 6954 10231 7352 11627
rect 7552 11423 7750 11425
rect 7552 11371 7564 11423
rect 7738 11371 7750 11423
rect 7552 11369 7750 11371
rect 7553 10030 7616 10397
rect 7950 10231 8348 11627
rect 8548 11423 8746 11425
rect 8548 11371 8560 11423
rect 8734 11371 8746 11423
rect 8548 11369 8746 11371
rect 8549 10030 8612 10397
rect 8946 10231 9344 11627
rect 9544 11423 9742 11425
rect 9544 11371 9556 11423
rect 9730 11371 9742 11423
rect 9544 11369 9742 11371
rect 592 9842 601 10022
rect 762 9842 771 10022
rect 592 9834 771 9842
rect 1164 9834 1668 10030
rect 2206 9834 2638 10030
rect 3202 9834 3634 10030
rect 4198 9834 4629 10030
rect 5194 9834 5625 10030
rect 6190 9834 6621 10030
rect 7186 9834 7616 10030
rect 8182 9834 8612 10030
rect 9178 9834 9556 10030
rect 9602 9834 9665 10397
rect 9942 10231 10340 11627
rect 10540 11423 10738 11425
rect 10540 11371 10552 11423
rect 10726 11371 10738 11423
rect 10540 11369 10738 11371
rect 10174 9834 10552 10030
rect 10598 9834 10661 10397
rect 10938 10231 11336 11627
rect 11536 11423 11734 11425
rect 11536 11371 11548 11423
rect 11722 11371 11734 11423
rect 11536 11369 11734 11371
rect 11536 10397 11548 10449
rect 11661 10397 11673 10449
rect 11934 10231 12909 11627
rect 11548 10030 11600 10032
rect 11170 10020 11600 10030
rect 11170 9845 11548 10020
rect 11170 9834 11600 9845
rect 12566 9834 12732 10030
rect 11548 9833 11600 9834
rect 201 9633 380 9679
rect 12778 9633 12909 10231
rect 201 9471 12909 9633
rect 201 8599 1080 9471
rect 1212 9326 2280 9334
rect 64759 9333 64773 12100
rect 1212 9148 1272 9326
rect 1462 9148 2280 9326
rect 1212 9134 2280 9148
rect 1811 8867 2027 8880
rect 1268 8815 1280 8867
rect 1454 8815 1466 8867
rect 1811 8815 1823 8867
rect 2014 8815 2027 8867
rect 1811 8803 2027 8815
rect 201 3957 380 8599
rect 580 8341 592 8393
rect 766 8341 778 8393
rect 581 5182 777 5184
rect 572 5180 787 5182
rect 572 5100 584 5180
rect 775 5100 787 5180
rect 978 5161 1068 8599
rect 1268 6630 1280 6689
rect 1454 6630 1466 6689
rect 1821 6477 2017 6643
rect 1267 6339 1467 6350
rect 1267 6164 1278 6339
rect 1456 6258 1467 6339
rect 1456 6164 2013 6258
rect 1267 6065 2013 6164
rect 572 5097 787 5100
rect 581 4169 777 5097
rect 973 3957 1068 5161
rect 1262 5160 1462 5162
rect 1262 5108 1275 5160
rect 1449 5108 1462 5160
rect 1262 5107 1462 5108
rect 1813 4343 2013 6065
rect 1813 4215 1822 4343
rect 2002 4215 2013 4343
rect 1813 4201 2013 4215
rect 201 45 1063 3957
rect 2094 2483 2184 6431
rect 64644 4675 64773 9333
rect 1815 2429 1827 2481
rect 2001 2429 2013 2481
rect 2094 2332 2265 2483
rect 1261 251 1275 303
rect 1449 251 1461 303
rect 1816 91 2012 257
rect 2213 45 2265 2332
rect 201 16 2265 45
rect 0 0 2265 16
rect 64759 14 64773 4675
rect 64959 14 64971 12100
rect 64759 1 64971 14
<< via1 >>
rect 15 16 201 12102
rect 592 11371 766 11423
rect 1588 11371 1762 11423
rect 2584 11371 2758 11423
rect 3580 11371 3754 11423
rect 4576 11371 4750 11423
rect 5572 11371 5746 11423
rect 6568 11371 6742 11423
rect 7564 11371 7738 11423
rect 8560 11371 8734 11423
rect 9556 11371 9730 11423
rect 601 9842 762 10022
rect 10552 11371 10726 11423
rect 11548 11371 11722 11423
rect 11548 10397 11661 10449
rect 11548 9845 11600 10020
rect 1272 9148 1462 9326
rect 1280 8815 1454 8867
rect 1823 8815 2014 8867
rect 592 8341 766 8393
rect 584 5100 775 5180
rect 1280 6630 1454 6689
rect 1278 6164 1456 6339
rect 1275 5108 1449 5160
rect 1822 4215 2002 4343
rect 1827 2429 2001 2481
rect 1275 251 1449 303
rect 64773 14 64959 12100
<< metal2 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 16 212 12102
rect 580 11423 778 12117
rect 580 11371 592 11423
rect 766 11371 778 11423
rect 580 11369 778 11371
rect 1576 11423 1774 12117
rect 1576 11371 1588 11423
rect 1762 11371 1774 11423
rect 1576 11369 1774 11371
rect 2572 11423 2770 12117
rect 2572 11371 2584 11423
rect 2758 11371 2770 11423
rect 2572 11369 2770 11371
rect 3568 11423 3766 12117
rect 3568 11371 3580 11423
rect 3754 11371 3766 11423
rect 3568 11369 3766 11371
rect 4564 11423 4762 12117
rect 4564 11371 4576 11423
rect 4750 11371 4762 11423
rect 4564 11369 4762 11371
rect 5560 11423 5758 12117
rect 5560 11371 5572 11423
rect 5746 11371 5758 11423
rect 5560 11369 5758 11371
rect 6556 11423 6754 12117
rect 6556 11371 6568 11423
rect 6742 11371 6754 11423
rect 6556 11369 6754 11371
rect 7552 11423 7750 12117
rect 7552 11371 7564 11423
rect 7738 11371 7750 11423
rect 7552 11369 7750 11371
rect 8548 11423 8746 12117
rect 8548 11371 8560 11423
rect 8734 11371 8746 11423
rect 8548 11369 8746 11371
rect 9544 11423 9742 12117
rect 9544 11371 9556 11423
rect 9730 11371 9742 11423
rect 9544 11369 9742 11371
rect 10540 11423 10738 12117
rect 10540 11371 10552 11423
rect 10726 11371 10738 11423
rect 10540 11369 10738 11371
rect 11536 11423 11734 12117
rect 51536 11510 51733 12118
rect 11536 11371 11548 11423
rect 11722 11371 11734 11423
rect 11536 11369 11734 11371
rect 51535 11369 51733 11510
rect 64759 12100 64971 12118
rect 51535 10998 51732 11369
rect 51535 10774 51536 10998
rect 51731 10774 51732 10998
rect 51535 10761 51732 10774
rect 11524 10449 11673 10453
rect 11524 10397 11548 10449
rect 11661 10397 11673 10449
rect 11524 10384 11673 10397
rect 578 10022 779 10051
rect 578 9842 601 10022
rect 762 9842 779 10022
rect 578 8393 779 9842
rect 11524 10020 11610 10384
rect 11524 9845 11548 10020
rect 11600 9845 11610 10020
rect 11524 9821 11610 9845
rect 1264 9326 1468 9338
rect 1264 9148 1272 9326
rect 1462 9148 1468 9326
rect 1264 8867 1468 9148
rect 1264 8815 1280 8867
rect 1454 8815 1468 8867
rect 1264 8810 1468 8815
rect 1808 8867 1968 8884
rect 1808 8815 1823 8867
rect 1808 8799 1968 8815
rect 578 8341 592 8393
rect 766 8341 779 8393
rect 578 8337 779 8341
rect 1267 6689 1467 6695
rect 1267 6630 1280 6689
rect 1454 6630 1467 6689
rect 1267 6339 1467 6630
rect 1267 6164 1278 6339
rect 1456 6164 1467 6339
rect 1267 6152 1467 6164
rect 572 5180 1968 5182
rect 572 5100 584 5180
rect 775 5160 1968 5180
rect 775 5108 1275 5160
rect 1449 5108 1968 5160
rect 775 5100 1968 5108
rect 572 5097 1968 5100
rect 1814 4343 2013 4352
rect 1814 4215 1822 4343
rect 2002 4215 2013 4343
rect 1814 2481 2013 4215
rect 1814 2429 1827 2481
rect 2001 2429 2013 2481
rect 1814 2427 2013 2429
rect 1261 303 1462 309
rect 1261 251 1275 303
rect 1449 251 1462 303
rect 1261 231 1462 251
rect 24450 231 24640 238
rect 1261 227 24640 231
rect 1261 113 24460 227
rect 24630 113 24640 227
rect 1261 108 24640 113
rect 24450 103 24640 108
rect 0 0 212 16
rect 64759 14 64773 12100
rect 64959 14 64971 12100
rect 64759 1 64971 14
<< via2 >>
rect 15 16 201 12102
rect 51536 10774 51731 10998
rect 51556 7464 52428 8364
rect 24456 485 24656 839
rect 24460 113 24630 227
rect 64773 14 64959 12100
<< metal3 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 16 212 12102
rect 64759 12100 64971 12118
rect 51535 10998 51732 11008
rect 51535 10774 51536 10998
rect 51731 10774 51732 10998
rect 51535 8385 51732 10774
rect 51535 8364 52452 8385
rect 51535 7464 51556 8364
rect 52428 7464 52452 8364
rect 51535 7435 52452 7464
rect 24456 839 24656 849
rect 24456 238 24656 485
rect 24450 227 24656 238
rect 24450 113 24460 227
rect 24630 113 24656 227
rect 24450 108 24656 113
rect 24450 103 24640 108
rect 0 0 212 16
rect 64759 14 64773 12100
rect 64959 14 64971 12100
rect 64759 1 64971 14
<< via3 >>
rect 15 16 201 12102
rect 64773 14 64959 12100
<< metal4 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 16 212 12102
rect 0 0 212 16
rect 64759 12100 64971 12118
rect 64759 14 64773 12100
rect 64959 14 64971 12100
rect 64759 1 64971 14
use opamp_chonky  x1
timestamp 1762910833
transform 1 0 1968 0 1 0
box 0 0 62677 9333
use ppolyf_u_1k_6p0_QZFH4C  XR1
timestamp 1763231934
transform 1 0 11635 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR2
timestamp 1763231934
transform 1 0 10639 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR3
timestamp 1763231934
transform 1 0 9643 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR4
timestamp 1763231934
transform 1 0 8647 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR5
timestamp 1763231934
transform 1 0 7651 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR6
timestamp 1763231934
transform 1 0 6655 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR7
timestamp 1763231934
transform 1 0 5659 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR8
timestamp 1763231934
transform 1 0 4663 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR9
timestamp 1763231934
transform 1 0 3667 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR10
timestamp 1763231934
transform 1 0 2671 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR11
timestamp 1763231934
transform 1 0 1675 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR12
timestamp 1763231934
transform 1 0 679 0 1 10906
box -344 -766 344 766
use ppolyf_u_1k_6p0_QZFH4C  XR13
timestamp 1763231934
transform 0 1 12057 -1 0 9932
box -344 -766 344 766
use ppolyf_u_1k_6p0_YUFH2C  XR14
timestamp 1763231934
transform 0 1 10861 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR15
timestamp 1763231934
transform 0 1 9865 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR16
timestamp 1763231934
transform 0 1 8869 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR17
timestamp 1763231934
transform 0 1 7873 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR18
timestamp 1763231934
transform 0 1 6877 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR19
timestamp 1763231934
transform 0 1 5881 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR20
timestamp 1763231934
transform 0 1 4885 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR21
timestamp 1763231934
transform 0 1 3889 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR22
timestamp 1763231934
transform 0 1 2893 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR23
timestamp 1763231934
transform 0 1 1897 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_YUFH2C  XR24
timestamp 1763231934
transform 0 1 901 -1 0 9932
box -344 -566 344 566
use ppolyf_u_1k_6p0_KPKJWY  XR26
timestamp 1762910469
transform 1 0 1919 0 1 7752
box -344 -1366 344 1366
use ppolyf_u_1k_6p0_KPKJWY  XR27
timestamp 1762910469
transform 1 0 1914 0 1 1366
box -344 -1366 344 1366
use ppolyf_u_1k_6p0_KPKJWY  XR28
timestamp 1762910469
transform 1 0 1367 0 1 7752
box -344 -1366 344 1366
use ppolyf_u_1k_6p0_QRJAJP  XR29
timestamp 1763230762
transform 1 0 1362 0 1 2706
box -344 -2706 344 2706
use ppolyf_u_1k_6p0_LRJJWQ  XR30
timestamp 1762910469
transform 1 0 679 0 1 6278
box -344 -2366 344 2366
<< labels >>
flabel metal2 51536 11369 51733 12118 0 FreeSans 200 0 0 0 OUT
port 1 nsew signal output
flabel metal2 11536 11369 11734 12117 0 FreeSans 200 0 0 0 D0
port 2 nsew signal input
flabel metal2 10540 11369 10738 12117 0 FreeSans 200 0 0 0 D1
port 3 nsew signal input
flabel metal2 9544 11369 9742 12117 0 FreeSans 200 0 0 0 D2
port 4 nsew signal input
flabel metal2 8548 11369 8746 12117 0 FreeSans 200 0 0 0 D3
port 5 nsew signal input
flabel metal2 7552 11369 7750 12117 0 FreeSans 200 0 0 0 D4
port 6 nsew signal input
flabel metal2 6556 11369 6754 12117 0 FreeSans 200 0 0 0 D5
port 7 nsew signal input
flabel metal2 5560 11369 5758 12117 0 FreeSans 200 0 0 0 D6
port 8 nsew signal input
flabel metal2 4564 11369 4762 12117 0 FreeSans 200 0 0 0 D7
port 9 nsew signal input
flabel metal2 3568 11369 3766 12117 0 FreeSans 200 0 0 0 D8
port 10 nsew signal input
flabel metal2 2572 11369 2770 12117 0 FreeSans 200 0 0 0 D9
port 11 nsew signal input
flabel metal2 1576 11369 1774 12117 0 FreeSans 200 0 0 0 D10
port 12 nsew signal input
flabel metal2 580 11369 778 12117 0 FreeSans 200 0 0 0 D11
port 13 nsew signal input
flabel metal4 64759 1 64971 12118 0 FreeSans 400 0 0 0 VDD
port 14 nsew power bidirectional
flabel metal4 0 0 212 12117 0 FreeSans 400 0 0 0 VSS
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 64971 12118
<< end >>
