* NGSPICE file created from flattened.ext - technology: gf180mcuD

.subckt r2r_dac_buffered_spice OUT D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 VDD VSS
X0 VDD.t48 x1.ADJ.t3 OUT.t34 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X1 x1.PLUS.t0 VSS.t7 VSS.t6 ppolyf_u_1k_6p0 r_width=1u r_length=10u
X2 VDD.t47 x1.ADJ.t4 OUT.t10 VDD.t4 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X3 a_6081_9832# a_7077_9832# VSS.t27 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X4 VSS.t53 a_3162_2792.t2 OUT.t69 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X5 OUT.t61 a_3162_2792.t3 VSS.t42 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X6 OUT.t62 a_3162_2792.t4 VSS.t43 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X7 OUT.t76 a_3162_2792.t5 VSS.t64 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X8 VDD.t46 x1.ADJ.t5 OUT.t8 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X9 OUT.t23 x1.ADJ.t6 VDD.t45 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X10 VSS.t65 a_3162_2792.t6 OUT.t77 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X11 VSS.t71 a_3162_2792.t7 OUT.t82 VSS.t2 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X12 x1.ADJ.t2 VSS.t29 VSS.t28 ppolyf_u_1k_6p0 r_width=1u r_length=10u
X13 VDD.t44 x1.ADJ.t7 OUT.t17 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X14 OUT.t11 x1.ADJ.t8 VDD.t43 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X15 OUT.t24 x1.ADJ.t9 VDD.t42 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X16 VDD.t41 x1.ADJ.t10 OUT.t18 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X17 D4.t0 a_7077_9832# VSS.t50 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X18 VSS.t72 a_3162_2792.t8 OUT.t83 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X19 OUT.t59 a_3162_2792.t9 VSS.t40 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X20 OUT.t60 a_3162_2792.t10 VSS.t41 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X21 VSS.t47 a_3162_2792.t11 OUT.t65 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X22 x1.MINUS.t1 OUT.t84 VSS.t80 ppolyf_u_1k_6p0 r_width=1u r_length=23.4u
X23 VSS.t48 a_3162_2792.t12 OUT.t66 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X24 VDD.t40 x1.ADJ.t11 OUT.t22 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X25 OUT.t13 x1.ADJ.t12 VDD.t39 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X26 VDD.t38 x1.ADJ.t13 OUT.t19 VDD.t9 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X27 OUT.t70 a_3162_2792.t13 VSS.t54 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X28 D8.t0 a_3093_9832# VSS.t73 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X29 VSS.t55 a_3162_2792.t14 OUT.t71 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X30 VDD.t29 x1.ADJ.t14 OUT.t25 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X31 VSS.t36 a_3162_2792.t15 OUT.t55 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X32 VSS.t37 a_3162_2792.t16 OUT.t56 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X33 OUT.t74 a_3162_2792.t17 VSS.t62 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X34 OUT.t75 a_3162_2792.t18 VSS.t63 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X35 VSS.t69 a_3162_2792.t19 OUT.t80 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X36 OUT.t28 x1.ADJ.t15 VDD.t37 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X37 a_10065_9832# a_11061_9832# VSS.t30 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X38 VSS.t70 a_3162_2792.t20 OUT.t81 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X39 a_579_8278# a_1101_9832# VSS.t79 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X40 a_5085_9832# a_6081_9832# VSS.t33 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X41 VSS.t38 a_3162_2792.t21 OUT.t57 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X42 OUT.t58 a_3162_2792.t22 VSS.t39 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X43 OUT.t29 x1.ADJ.t16 VDD.t36 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X44 VDD.t35 x1.ADJ.t17 OUT.t44 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X45 D7.t0 a_4089_9832# VSS.t26 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X46 D1.t0 a_10065_9832# VSS.t66 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X47 VSS.t45 a_3162_2792.t23 OUT.t63 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X48 OUT.t64 a_3162_2792.t24 VSS.t46 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X49 VSS.t51 a_3162_2792.t25 OUT.t67 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X50 OUT.t68 a_3162_2792.t26 VSS.t52 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X51 VDD.t34 x1.ADJ.t18 OUT.t6 VDD.t0 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X52 a_4089_9832# a_5085_9832# VSS.t56 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X53 VDD.t33 x1.ADJ.t19 OUT.t14 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X54 OUT.t53 a_3162_2792.t27 VSS.t34 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X55 a_2576_5968.t2 x1.MINUS.t2 a_2442_2792.t2 VDD.t51 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X56 VSS.t76 a_2442_2792.t0 a_2442_2792.t1 VSS.t75 nfet_05v0 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=0.6u
X57 OUT.t15 x1.ADJ.t20 VDD.t32 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X58 OUT.t54 a_3162_2792.t28 VSS.t35 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X59 VSS.t60 a_3162_2792.t29 OUT.t72 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X60 a_3093_9832# a_4089_9832# VSS.t9 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X61 VDD.t31 x1.ADJ.t21 OUT.t39 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X62 OUT.t5 x1.ADJ.t22 VDD.t30 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X63 D11.t0 a_579_8278# VSS.t25 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X64 a_579_8278# x1.MINUS.t0 VSS.t11 ppolyf_u_1k_6p0 r_width=1u r_length=20u
X65 VDD.t28 x1.ADJ.t23 a_2576_5968.t0 VDD.t27 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X66 D0.t0 a_11061_9832# VSS.t44 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X67 VDD.t26 x1.ADJ.t24 OUT.t41 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X68 OUT.t4 x1.ADJ.t25 VDD.t14 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X69 VDD.t49 x1.PLUS.t1 VSS.t57 ppolyf_u_1k_6p0 r_width=1u r_length=10u
X70 a_9069_9832# a_10065_9832# VSS.t49 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X71 VSS.t61 a_3162_2792.t30 OUT.t73 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X72 OUT.t20 x1.ADJ.t26 VDD.t25 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X73 VDD.t24 x1.ADJ.t27 OUT.t40 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X74 D3.t0 a_8073_9832# VSS.t15 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X75 VDD.t23 x1.ADJ.t28 OUT.t45 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X76 VSS.t67 a_3162_2792.t31 OUT.t78 VSS.t13 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X77 OUT.t30 x1.ADJ.t29 VDD.t22 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X78 VDD.t21 x1.ADJ.t30 OUT.t35 VDD.t4 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X79 D10.t0 a_1101_9832# VSS.t19 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X80 VSS.t68 a_3162_2792.t32 OUT.t79 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X81 OUT.t47 a_3162_2792.t33 VSS.t17 VSS.t2 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X82 VDD.t20 x1.ADJ.t31 OUT.t43 VDD.t9 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X83 a_8073_9832# a_9069_9832# VSS.t24 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X84 VDD.t19 x1.ADJ.t32 OUT.t36 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X85 OUT.t27 x1.ADJ.t33 VDD.t18 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X86 VDD.t17 x1.ADJ.t34 OUT.t9 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X87 OUT.t7 x1.ADJ.t35 VDD.t16 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X88 OUT.t48 a_3162_2792.t34 VSS.t18 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X89 OUT.t51 a_3162_2792.t35 VSS.t22 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X90 VSS.t23 a_3162_2792.t36 OUT.t52 VSS.t0 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X91 D2.t0 a_9069_9832# VSS.t5 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X92 VSS.t20 a_3162_2792.t37 OUT.t49 VSS.t13 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X93 a_3162_2792.t0 x1.PLUS.t2 a_2576_5968.t1 VDD.t50 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X94 D9.t0 a_2097_9832# VSS.t4 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X95 D6.t0 a_5085_9832# VSS.t32 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X96 VDD.t15 x1.ADJ.t36 OUT.t33 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X97 a_2097_9832# a_3093_9832# VSS.t10 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X98 a_3162_2792.t1 a_2442_2792.t3 VSS.t78 VSS.t77 nfet_05v0 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=0.6u
X99 OUT.t50 a_3162_2792.t38 VSS.t21 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X100 VDD.t13 x1.ADJ.t0 x1.ADJ.t1 VDD.t12 pfet_05v0 ad=6.16p pd=28.88u as=6.16p ps=28.88u w=14u l=0.6u
X101 OUT.t2 a_3162_2792.t39 VSS.t12 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X102 VSS.t14 a_3162_2792.t40 OUT.t3 VSS.t13 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X103 OUT.t26 x1.ADJ.t37 VDD.t11 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X104 OUT.t31 x1.ADJ.t38 VDD.t10 VDD.t9 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X105 a_1101_9832# a_2097_9832# VSS.t8 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X106 VSS.t1 a_3162_2792.t41 OUT.t0 VSS.t0 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X107 VSS.t3 a_3162_2792.t42 OUT.t1 VSS.t2 nfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X108 VDD.t8 x1.ADJ.t39 OUT.t42 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=44p ps=0.20088m w=100u l=0.6u
X109 OUT.t16 x1.ADJ.t40 VDD.t7 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X110 a_7077_9832# a_8073_9832# VSS.t31 ppolyf_u_1k_6p0 r_width=1u r_length=2u
X111 D5.t0 a_6081_9832# VSS.t74 ppolyf_u_1k_6p0 r_width=1u r_length=4u
X112 VSS.t16 a_3162_2792.t43 OUT.t46 VSS.t0 nfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X113 OUT.t32 x1.ADJ.t41 VDD.t6 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X114 VDD.t5 x1.ADJ.t42 OUT.t21 VDD.t4 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X115 VDD.t3 x1.ADJ.t43 OUT.t38 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X116 OUT.t37 x1.ADJ.t44 VDD.t2 VDD.t0 pfet_05v0 ad=26p pd=0.10052m as=26p ps=0.10052m w=100u l=0.6u
X117 VDD.t1 x1.ADJ.t45 OUT.t12 VDD.t0 pfet_05v0 ad=44p pd=0.20088m as=26p ps=0.10052m w=100u l=0.6u
X118 a_11061_9832# VSS.t59 VSS.t58 ppolyf_u_1k_6p0 r_width=1u r_length=4u
R0 x1.ADJ.t30 x1.ADJ.n25 620.038
R1 x1.ADJ.t32 x1.ADJ.n4 620.038
R2 x1.ADJ.n57 x1.ADJ.t24 620.038
R3 x1.ADJ.n42 x1.ADJ.t4 620.038
R4 x1.ADJ.n14 x1.ADJ.t45 620.006
R5 x1.ADJ.t39 x1.ADJ.n52 620.006
R6 x1.ADJ.t5 x1.ADJ.n69 620.006
R7 x1.ADJ.t18 x1.ADJ.n39 620.006
R8 x1.ADJ.t29 x1.ADJ.n42 619.74
R9 x1.ADJ.n39 x1.ADJ.t44 619.74
R10 x1.ADJ.t19 x1.ADJ.n35 619.74
R11 x1.ADJ.t36 x1.ADJ.n30 619.74
R12 x1.ADJ.n50 x1.ADJ.t15 619.74
R13 x1.ADJ.n64 x1.ADJ.t33 619.74
R14 x1.ADJ.t7 x1.ADJ.n58 619.74
R15 x1.ADJ.t21 x1.ADJ.n31 619.74
R16 x1.ADJ.n69 x1.ADJ.t40 619.74
R17 x1.ADJ.t25 x1.ADJ.n4 619.74
R18 x1.ADJ.n68 x1.ADJ.t17 619.74
R19 x1.ADJ.n79 x1.ADJ.t42 619.74
R20 x1.ADJ.t22 x1.ADJ.n9 619.74
R21 x1.ADJ.t8 x1.ADJ.n3 619.74
R22 x1.ADJ.n25 x1.ADJ.t20 619.74
R23 x1.ADJ.n14 x1.ADJ.t37 619.74
R24 x1.ADJ.t28 x1.ADJ.n12 619.74
R25 x1.ADJ.t43 x1.ADJ.n15 619.74
R26 x1.ADJ.n52 x1.ADJ.t16 619.74
R27 x1.ADJ.n57 x1.ADJ.t41 619.74
R28 x1.ADJ.n43 x1.ADJ.t12 614.254
R29 x1.ADJ.n43 x1.ADJ.t29 614.254
R30 x1.ADJ.n38 x1.ADJ.t12 614.254
R31 x1.ADJ.t44 x1.ADJ.n38 614.254
R32 x1.ADJ.n46 x1.ADJ.t3 614.254
R33 x1.ADJ.n46 x1.ADJ.t19 614.254
R34 x1.ADJ.t3 x1.ADJ.n45 614.254
R35 x1.ADJ.n45 x1.ADJ.t36 614.254
R36 x1.ADJ.n49 x1.ADJ.t38 614.254
R37 x1.ADJ.t15 x1.ADJ.n49 614.254
R38 x1.ADJ.n63 x1.ADJ.t38 614.254
R39 x1.ADJ.t33 x1.ADJ.n63 614.254
R40 x1.ADJ.t34 x1.ADJ.n59 614.254
R41 x1.ADJ.n59 x1.ADJ.t7 614.254
R42 x1.ADJ.n60 x1.ADJ.t34 614.254
R43 x1.ADJ.n60 x1.ADJ.t21 614.254
R44 x1.ADJ.n74 x1.ADJ.t40 614.254
R45 x1.ADJ.t9 x1.ADJ.n74 614.254
R46 x1.ADJ.n75 x1.ADJ.t9 614.254
R47 x1.ADJ.n75 x1.ADJ.t25 614.254
R48 x1.ADJ.t17 x1.ADJ.n67 614.254
R49 x1.ADJ.n67 x1.ADJ.t27 614.254
R50 x1.ADJ.n78 x1.ADJ.t27 614.254
R51 x1.ADJ.t42 x1.ADJ.n78 614.254
R52 x1.ADJ.n17 x1.ADJ.t22 614.254
R53 x1.ADJ.n17 x1.ADJ.t35 614.254
R54 x1.ADJ.t35 x1.ADJ.n16 614.254
R55 x1.ADJ.n16 x1.ADJ.t8 614.254
R56 x1.ADJ.n24 x1.ADJ.t6 614.254
R57 x1.ADJ.t20 x1.ADJ.n24 614.254
R58 x1.ADJ.t37 x1.ADJ.n13 614.254
R59 x1.ADJ.n13 x1.ADJ.t6 614.254
R60 x1.ADJ.n21 x1.ADJ.t11 614.254
R61 x1.ADJ.n21 x1.ADJ.t28 614.254
R62 x1.ADJ.n20 x1.ADJ.t43 614.254
R63 x1.ADJ.t11 x1.ADJ.n20 614.254
R64 x1.ADJ.n27 x1.ADJ.t45 614.254
R65 x1.ADJ.n27 x1.ADJ.t13 614.254
R66 x1.ADJ.t13 x1.ADJ.n26 614.254
R67 x1.ADJ.n26 x1.ADJ.t30 614.254
R68 x1.ADJ.t14 x1.ADJ.n70 614.254
R69 x1.ADJ.n70 x1.ADJ.t32 614.254
R70 x1.ADJ.n71 x1.ADJ.t5 614.254
R71 x1.ADJ.n71 x1.ADJ.t14 614.254
R72 x1.ADJ.t16 x1.ADJ.n51 614.254
R73 x1.ADJ.n51 x1.ADJ.t26 614.254
R74 x1.ADJ.n56 x1.ADJ.t26 614.254
R75 x1.ADJ.t41 x1.ADJ.n56 614.254
R76 x1.ADJ.n54 x1.ADJ.t24 614.254
R77 x1.ADJ.n41 x1.ADJ.t31 614.254
R78 x1.ADJ.t4 x1.ADJ.n41 614.254
R79 x1.ADJ.t31 x1.ADJ.n40 614.254
R80 x1.ADJ.n40 x1.ADJ.t18 614.254
R81 x1.ADJ.n53 x1.ADJ.t39 614.254
R82 x1.ADJ.t10 x1.ADJ.n53 614.254
R83 x1.ADJ.n54 x1.ADJ.t10 614.254
R84 x1.ADJ.t23 x1.ADJ.n86 101.537
R85 x1.ADJ.n87 x1.ADJ.t23 101.079
R86 x1.ADJ.t0 x1.ADJ.n83 101.079
R87 x1.ADJ.n84 x1.ADJ.t0 101.076
R88 x1.ADJ.n65 x1.ADJ.n29 15.7436
R89 x1.ADJ.n82 x1.ADJ.n2 14.7961
R90 x1.ADJ.n29 x1.ADJ.n2 14.6668
R91 x1.ADJ x1.ADJ.t2 9.44369
R92 x1.ADJ.n53 x1.ADJ.n33 5.13335
R93 x1.ADJ.n55 x1.ADJ.n54 5.13335
R94 x1.ADJ.n41 x1.ADJ.n36 5.02611
R95 x1.ADJ.n56 x1.ADJ.n55 5.02611
R96 x1.ADJ.n40 x1.ADJ.n8 5.02611
R97 x1.ADJ.n44 x1.ADJ.n43 5.02611
R98 x1.ADJ.n38 x1.ADJ.n37 5.02611
R99 x1.ADJ.n47 x1.ADJ.n46 5.02611
R100 x1.ADJ.n45 x1.ADJ.n32 5.02611
R101 x1.ADJ.n49 x1.ADJ.n48 5.02611
R102 x1.ADJ.n63 x1.ADJ.n62 5.02611
R103 x1.ADJ.n59 x1.ADJ.n34 5.02611
R104 x1.ADJ.n61 x1.ADJ.n60 5.02611
R105 x1.ADJ.n72 x1.ADJ.n71 5.02611
R106 x1.ADJ.n70 x1.ADJ.n6 5.02611
R107 x1.ADJ.n76 x1.ADJ.n75 5.02611
R108 x1.ADJ.n74 x1.ADJ.n73 5.02611
R109 x1.ADJ.n78 x1.ADJ.n77 5.02611
R110 x1.ADJ.n67 x1.ADJ.n7 5.02611
R111 x1.ADJ.n16 x1.ADJ.n5 5.02611
R112 x1.ADJ.n18 x1.ADJ.n17 5.02611
R113 x1.ADJ.n26 x1.ADJ.n11 5.02611
R114 x1.ADJ.n28 x1.ADJ.n27 5.02611
R115 x1.ADJ.n13 x1.ADJ.n10 5.02611
R116 x1.ADJ.n24 x1.ADJ.n23 5.02611
R117 x1.ADJ.n20 x1.ADJ.n19 5.02611
R118 x1.ADJ.n22 x1.ADJ.n21 5.02611
R119 x1.ADJ.n51 x1.ADJ.n33 5.02611
R120 x1.ADJ.n65 x1.ADJ.n64 2.82526
R121 x1.ADJ.n81 x1.ADJ.n1 2.35383
R122 x1.ADJ.n86 x1.ADJ.n85 1.5858
R123 x1.ADJ.n85 x1.ADJ.n0 1.5511
R124 x1.ADJ.n82 x1.ADJ.n81 0.8605
R125 x1.ADJ x1.ADJ.n87 0.800244
R126 x1.ADJ.n84 x1.ADJ.n1 0.649885
R127 x1.ADJ.n83 x1.ADJ.n82 0.533174
R128 x1.ADJ.n50 x1.ADJ.n1 0.471929
R129 x1.ADJ.n85 x1.ADJ.t1 0.470597
R130 x1.ADJ.n72 x1.ADJ.n8 0.437096
R131 x1.ADJ.n36 x1.ADJ.n6 0.437096
R132 x1.ADJ.n87 x1.ADJ.n0 0.401314
R133 x1.ADJ.n66 x1.ADJ.n65 0.321929
R134 x1.ADJ.n81 x1.ADJ.n80 0.321929
R135 x1.ADJ.n25 x1.ADJ.n12 0.298623
R136 x1.ADJ.n12 x1.ADJ.n3 0.298623
R137 x1.ADJ.n79 x1.ADJ.n4 0.298623
R138 x1.ADJ.n58 x1.ADJ.n57 0.298623
R139 x1.ADJ.n58 x1.ADJ.n50 0.298623
R140 x1.ADJ.n50 x1.ADJ.n35 0.298623
R141 x1.ADJ.n42 x1.ADJ.n35 0.298623
R142 x1.ADJ.n80 x1.ADJ.n79 0.295483
R143 x1.ADJ.n15 x1.ADJ.n9 0.26697
R144 x1.ADJ.n15 x1.ADJ.n14 0.26697
R145 x1.ADJ.n69 x1.ADJ.n68 0.26697
R146 x1.ADJ.n39 x1.ADJ.n30 0.26697
R147 x1.ADJ.n64 x1.ADJ.n30 0.26697
R148 x1.ADJ.n64 x1.ADJ.n31 0.26697
R149 x1.ADJ.n52 x1.ADJ.n31 0.26697
R150 x1.ADJ.n68 x1.ADJ.n66 0.26383
R151 x1.ADJ.n29 x1.ADJ.n28 0.148426
R152 x1.ADJ.n11 x1.ADJ.n2 0.148426
R153 x1.ADJ.n83 x1.ADJ.n0 0.1355
R154 x1.ADJ.n86 x1.ADJ.n84 0.120962
R155 x1.ADJ.n28 x1.ADJ.n10 0.107734
R156 x1.ADJ.n19 x1.ADJ.n10 0.107734
R157 x1.ADJ.n19 x1.ADJ.n18 0.107734
R158 x1.ADJ.n18 x1.ADJ.n7 0.107734
R159 x1.ADJ.n73 x1.ADJ.n7 0.107734
R160 x1.ADJ.n73 x1.ADJ.n72 0.107734
R161 x1.ADJ.n37 x1.ADJ.n8 0.107734
R162 x1.ADJ.n37 x1.ADJ.n32 0.107734
R163 x1.ADJ.n62 x1.ADJ.n32 0.107734
R164 x1.ADJ.n62 x1.ADJ.n61 0.107734
R165 x1.ADJ.n61 x1.ADJ.n33 0.107734
R166 x1.ADJ.n23 x1.ADJ.n11 0.107734
R167 x1.ADJ.n23 x1.ADJ.n22 0.107734
R168 x1.ADJ.n22 x1.ADJ.n5 0.107734
R169 x1.ADJ.n77 x1.ADJ.n5 0.107734
R170 x1.ADJ.n77 x1.ADJ.n76 0.107734
R171 x1.ADJ.n76 x1.ADJ.n6 0.107734
R172 x1.ADJ.n44 x1.ADJ.n36 0.107734
R173 x1.ADJ.n47 x1.ADJ.n44 0.107734
R174 x1.ADJ.n48 x1.ADJ.n47 0.107734
R175 x1.ADJ.n48 x1.ADJ.n34 0.107734
R176 x1.ADJ.n55 x1.ADJ.n34 0.107734
R177 x1.ADJ.n80 x1.ADJ.n3 0.00363953
R178 x1.ADJ.n66 x1.ADJ.n9 0.00363953
R179 OUT.n63 OUT.n61 34.1284
R180 OUT.n44 OUT.n42 34.1273
R181 OUT.n82 OUT.n80 34.1273
R182 OUT.n76 OUT.n74 34.1267
R183 OUT.n37 OUT.n35 34.1262
R184 OUT.n71 OUT.n70 34.1245
R185 OUT.n87 OUT.n86 34.1245
R186 OUT.n97 OUT.n95 34.1225
R187 OUT.n16 OUT.n15 34.1225
R188 OUT.n48 OUT.n47 34.1206
R189 OUT.n11 OUT.n10 34.1206
R190 OUT.n27 OUT.n25 34.1186
R191 OUT.n93 OUT.n92 34.1167
R192 OUT.n53 OUT.n51 34.1147
R193 OUT.n58 OUT.n57 34.1147
R194 OUT.n20 OUT.n19 34.1089
R195 OUT.n66 OUT.t84 29.5912
R196 OUT.n59 OUT.t77 26.7643
R197 OUT.n21 OUT.t36 26.7629
R198 OUT.n99 OUT.n98 26.7616
R199 OUT.n2 OUT.n1 26.7616
R200 OUT.n33 OUT.n32 26.7596
R201 OUT.n8 OUT.n7 26.7596
R202 OUT.n49 OUT.t41 26.757
R203 OUT.n84 OUT.n83 26.7538
R204 OUT.n23 OUT.n22 26.7538
R205 OUT.n90 OUT.n18 26.7447
R206 OUT.n29 OUT.n28 26.7408
R207 OUT.n55 OUT.n54 26.7388
R208 OUT.n46 OUT.n45 26.7388
R209 OUT.n68 OUT.n40 26.7369
R210 OUT.n65 OUT.n64 26.7349
R211 OUT.n88 OUT.t71 26.6707
R212 OUT.n65 OUT.n63 7.71659
R213 OUT.n70 OUT.n68 7.71464
R214 OUT.n55 OUT.n53 7.71268
R215 OUT.n46 OUT.n44 7.71268
R216 OUT.n49 OUT.n48 7.71268
R217 OUT.n29 OUT.n27 7.71072
R218 OUT.n59 OUT.n58 7.70877
R219 OUT.n92 OUT.n90 7.70681
R220 OUT.n21 OUT.n20 7.70681
R221 OUT.n84 OUT.n82 7.7029
R222 OUT.n74 OUT.n23 7.7029
R223 OUT.n35 OUT.n33 7.69703
R224 OUT.n10 OUT.n8 7.69703
R225 OUT.n99 OUT.n97 7.69507
R226 OUT.n15 OUT.n2 7.69507
R227 OUT.n88 OUT.n87 7.59954
R228 OUT OUT.n100 1.97295
R229 OUT OUT.n0 0.109596
R230 OUT.n19 OUT.t8 0.0543631
R231 OUT.n57 OUT.t81 0.0534887
R232 OUT.n67 OUT.n59 0.0505
R233 OUT.n85 OUT.n23 0.0505
R234 OUT.n100 OUT.n2 0.0505
R235 OUT.n8 OUT.n3 0.0505
R236 OUT.n89 OUT.n88 0.0505
R237 OUT.n85 OUT.n84 0.0505
R238 OUT.n33 OUT.n3 0.0505
R239 OUT.n100 OUT.n99 0.0505
R240 OUT.n56 OUT.n49 0.0505
R241 OUT.n66 OUT.n65 0.0505
R242 OUT.n56 OUT.n46 0.0505
R243 OUT.n68 OUT.n67 0.0505
R244 OUT.n89 OUT.n21 0.0505
R245 OUT.n30 OUT.n29 0.0505
R246 OUT.n90 OUT.n89 0.0505
R247 OUT.n56 OUT.n55 0.0505
R248 OUT.n87 OUT.t73 0.0464575
R249 OUT.n86 OUT.t63 0.0464575
R250 OUT.n58 OUT.t55 0.0464575
R251 OUT.n47 OUT.t42 0.0459256
R252 OUT.n20 OUT.t25 0.0431131
R253 OUT.n48 OUT.t18 0.0431131
R254 OUT.n61 OUT.n31 0.0339259
R255 OUT.n11 OUT.n6 0.03289
R256 OUT.n51 OUT.n50 0.0319444
R257 OUT.n95 OUT.n4 0.0314837
R258 OUT.n16 OUT.n13 0.0314837
R259 OUT.n42 OUT.n31 0.0310915
R260 OUT.n80 OUT.n78 0.0310915
R261 OUT.n93 OUT.n17 0.0305381
R262 OUT.n97 OUT.n96 0.0300775
R263 OUT.n37 OUT.n36 0.0300775
R264 OUT.n35 OUT.n34 0.0300775
R265 OUT.n80 OUT.n79 0.0300775
R266 OUT.n82 OUT.n81 0.0300775
R267 OUT.n10 OUT.n9 0.0300775
R268 OUT.n15 OUT.n14 0.0300775
R269 OUT.n76 OUT.n75 0.0300775
R270 OUT.n74 OUT.n73 0.0300775
R271 OUT.n77 OUT.n76 0.0296852
R272 OUT.n25 OUT.n24 0.0291319
R273 OUT.n72 OUT.n37 0.028279
R274 OUT.n53 OUT.n52 0.0249131
R275 OUT.n92 OUT.n91 0.0249131
R276 OUT.n27 OUT.n26 0.0249131
R277 OUT.n71 OUT.n39 0.0249131
R278 OUT.n70 OUT.n69 0.0249131
R279 OUT.n42 OUT.n41 0.0249131
R280 OUT.n44 OUT.n43 0.0249131
R281 OUT.n61 OUT.n60 0.0249131
R282 OUT.n63 OUT.n62 0.0249131
R283 OUT.n57 OUT.n0 0.0240602
R284 OUT.n94 OUT.n16 0.0240602
R285 OUT.n12 OUT.n11 0.0240602
R286 OUT.n86 OUT.n5 0.0240602
R287 OUT.n95 OUT.n94 0.0240602
R288 OUT.n47 OUT.n38 0.0240602
R289 OUT.n72 OUT.n71 0.0240602
R290 OUT.n19 OUT.n0 0.0240602
R291 OUT.n25 OUT.n5 0.0240602
R292 OUT.n94 OUT.n93 0.0240602
R293 OUT.n51 OUT.n12 0.0240602
R294 OUT.n54 OUT.t35 0.0187
R295 OUT.n54 OUT.t15 0.0187
R296 OUT.n52 OUT.t19 0.0187
R297 OUT.n52 OUT.t23 0.0187
R298 OUT.n50 OUT.t12 0.0187
R299 OUT.n50 OUT.t26 0.0187
R300 OUT.n18 OUT.t45 0.0187
R301 OUT.n18 OUT.t11 0.0187
R302 OUT.n91 OUT.t22 0.0187
R303 OUT.n91 OUT.t7 0.0187
R304 OUT.n17 OUT.t38 0.0187
R305 OUT.n17 OUT.t5 0.0187
R306 OUT.n28 OUT.t21 0.0187
R307 OUT.n28 OUT.t4 0.0187
R308 OUT.n26 OUT.t40 0.0187
R309 OUT.n26 OUT.t24 0.0187
R310 OUT.n24 OUT.t44 0.0187
R311 OUT.n24 OUT.t16 0.0187
R312 OUT.n40 OUT.t10 0.0187
R313 OUT.n40 OUT.t30 0.0187
R314 OUT.n69 OUT.t43 0.0187
R315 OUT.n69 OUT.t13 0.0187
R316 OUT.n39 OUT.t6 0.0187
R317 OUT.n39 OUT.t37 0.0187
R318 OUT.n45 OUT.t14 0.0187
R319 OUT.n45 OUT.t28 0.0187
R320 OUT.n43 OUT.t34 0.0187
R321 OUT.n43 OUT.t31 0.0187
R322 OUT.n41 OUT.t33 0.0187
R323 OUT.n41 OUT.t27 0.0187
R324 OUT.n64 OUT.t17 0.0187
R325 OUT.n64 OUT.t32 0.0187
R326 OUT.n62 OUT.t9 0.0187
R327 OUT.n62 OUT.t20 0.0187
R328 OUT.n60 OUT.t39 0.0187
R329 OUT.n60 OUT.t29 0.0187
R330 OUT.n98 OUT.t49 0.01688
R331 OUT.n98 OUT.t74 0.01688
R332 OUT.n96 OUT.t82 0.01688
R333 OUT.n96 OUT.t47 0.01688
R334 OUT.n4 OUT.t0 0.01688
R335 OUT.n4 OUT.t68 0.01688
R336 OUT.n32 OUT.t65 0.01688
R337 OUT.n32 OUT.t62 0.01688
R338 OUT.n34 OUT.t72 0.01688
R339 OUT.n34 OUT.t58 0.01688
R340 OUT.n36 OUT.t80 0.01688
R341 OUT.n36 OUT.t60 0.01688
R342 OUT.n83 OUT.t3 0.01688
R343 OUT.n83 OUT.t51 0.01688
R344 OUT.n81 OUT.t66 0.01688
R345 OUT.n81 OUT.t76 0.01688
R346 OUT.n79 OUT.t46 0.01688
R347 OUT.n79 OUT.t2 0.01688
R348 OUT.n7 OUT.t78 0.01688
R349 OUT.n7 OUT.t48 0.01688
R350 OUT.n9 OUT.t1 0.01688
R351 OUT.n9 OUT.t61 0.01688
R352 OUT.n6 OUT.t52 0.01688
R353 OUT.n6 OUT.t50 0.01688
R354 OUT.n1 OUT.t56 0.01688
R355 OUT.n1 OUT.t59 0.01688
R356 OUT.n14 OUT.t79 0.01688
R357 OUT.n14 OUT.t54 0.01688
R358 OUT.n13 OUT.t67 0.01688
R359 OUT.n13 OUT.t75 0.01688
R360 OUT.n22 OUT.t69 0.01688
R361 OUT.n22 OUT.t70 0.01688
R362 OUT.n73 OUT.t57 0.01688
R363 OUT.n73 OUT.t64 0.01688
R364 OUT.n75 OUT.t83 0.01688
R365 OUT.n75 OUT.t53 0.01688
R366 OUT.n78 OUT.n31 0.000532943
R367 OUT.n12 OUT.n0 0.000532943
R368 OUT.n89 OUT.n3 0.000521962
R369 OUT.n72 OUT.n38 0.000521962
R370 OUT.n100 OUT.n3 0.000510981
R371 OUT.n89 OUT.n85 0.000510981
R372 OUT.n85 OUT.n30 0.000510981
R373 OUT.n56 OUT.n30 0.000510981
R374 OUT.n67 OUT.n56 0.000510981
R375 OUT.n67 OUT.n66 0.000510981
R376 OUT.n78 OUT.n77 0.000510981
R377 OUT.n77 OUT.n72 0.000510981
R378 OUT.n38 OUT.n5 0.000510981
R379 OUT.n94 OUT.n5 0.000510981
R380 OUT.n94 OUT.n12 0.000510981
R381 VDD.t9 VDD.t0 4343.5
R382 VDD.t9 VDD.t4 4343.5
R383 VDD.n25 VDD.t4 2223.27
R384 VDD.n27 VDD.n26 180.601
R385 VDD.n33 VDD.n27 180.601
R386 VDD.n23 VDD.n17 180.601
R387 VDD.n36 VDD.n17 180.601
R388 VDD.n26 VDD.n21 147.525
R389 VDD.n36 VDD.n34 147.525
R390 VDD.n27 VDD.n19 135.8
R391 VDD.n20 VDD.n19 135.8
R392 VDD.n34 VDD.n33 135.8
R393 VDD.n23 VDD.n21 135.8
R394 VDD.n38 VDD.n16 135.8
R395 VDD.n38 VDD.n17 135.8
R396 VDD.t50 VDD.n23 119.879
R397 VDD.t51 VDD.n36 119.879
R398 VDD.n37 VDD.t51 119.683
R399 VDD.n25 VDD.t12 54.9597
R400 VDD.t27 VDD.n18 35.4234
R401 VDD.n51 VDD.n49 34.1113
R402 VDD.n87 VDD.n85 34.1107
R403 VDD.n65 VDD.n63 34.1107
R404 VDD.n79 VDD.n77 34.1085
R405 VDD.n72 VDD.n70 34.1085
R406 VDD.n57 VDD.n55 34.1074
R407 VDD.n21 VDD.n20 33.0755
R408 VDD.n34 VDD.n16 33.0755
R409 VDD.t12 VDD.t50 28.7682
R410 VDD.t51 VDD.t27 28.7682
R411 VDD.t51 VDD.n33 26.3889
R412 VDD.n73 VDD.n10 25.7991
R413 VDD.n80 VDD.n75 25.7912
R414 VDD.n52 VDD.n47 25.7893
R415 VDD.n61 VDD.n46 25.7873
R416 VDD.n83 VDD.n7 25.7854
R417 VDD.n58 VDD.n53 25.7854
R418 VDD.n37 VDD.n18 20.1034
R419 VDD.t50 VDD.n24 17.9501
R420 VDD.n95 VDD.n94 14.5582
R421 VDD.n94 VDD.n2 14.3237
R422 VDD.n24 VDD.n18 13.3893
R423 VDD.n20 VDD.n16 11.7255
R424 VDD VDD.n97 11.1908
R425 VDD VDD.t49 11.0951
R426 VDD.n85 VDD.n83 6.59094
R427 VDD.n58 VDD.n57 6.59094
R428 VDD.n63 VDD.n61 6.58898
R429 VDD.n52 VDD.n51 6.58703
R430 VDD.n80 VDD.n79 6.58507
R431 VDD.n73 VDD.n72 6.57724
R432 VDD.n22 VDD.n15 4.0642
R433 VDD.n24 VDD.n19 3.71928
R434 VDD.n91 VDD.n90 3.34156
R435 VDD.n11 VDD.n3 3.08674
R436 VDD.n40 VDD.n39 3.06246
R437 VDD.n39 VDD.n15 3.06246
R438 VDD.n95 VDD 2.62963
R439 VDD.n35 VDD.n15 2.52779
R440 VDD.n4 VDD.n0 2.48004
R441 VDD.n8 VDD.n1 2.29184
R442 VDD.n97 VDD.n0 1.65155
R443 VDD.n89 VDD.n5 1.6489
R444 VDD.n35 VDD.n14 1.5575
R445 VDD.n96 VDD.n1 1.52562
R446 VDD.n44 VDD.n43 1.5244
R447 VDD.n30 VDD.n13 0.98945
R448 VDD.n41 VDD.n13 0.98945
R449 VDD.n22 VDD.n2 0.970069
R450 VDD.n91 VDD.n4 0.862023
R451 VDD.n8 VDD.n3 0.795398
R452 VDD.n42 VDD.n41 0.695065
R453 VDD.n40 VDD.n14 0.695065
R454 VDD.n32 VDD.n14 0.6357
R455 VDD.n32 VDD.n31 0.6265
R456 VDD.n97 VDD.n96 0.424107
R457 VDD.n28 VDD.n12 0.380551
R458 VDD.n12 VDD.t13 0.303833
R459 VDD.n13 VDD.t28 0.303833
R460 VDD.n43 VDD.n42 0.27616
R461 VDD.n41 VDD.n40 0.262674
R462 VDD.n5 VDD 0.262078
R463 VDD.n42 VDD.n2 0.261707
R464 VDD.n29 VDD 0.217474
R465 VDD.n36 VDD.n35 0.197375
R466 VDD.n33 VDD.n32 0.197375
R467 VDD.n19 VDD.n13 0.197375
R468 VDD.n39 VDD.n38 0.197375
R469 VDD.n38 VDD.n37 0.197375
R470 VDD.n23 VDD.n22 0.197375
R471 VDD.n26 VDD.n12 0.197375
R472 VDD.n26 VDD.n25 0.197375
R473 VDD.n31 VDD.n30 0.13595
R474 VDD.n96 VDD.n95 0.132454
R475 VDD.n30 VDD.n29 0.110525
R476 VDD.n43 VDD.n12 0.108972
R477 VDD.n82 VDD.n4 0.0547889
R478 VDD.n59 VDD.n52 0.0547889
R479 VDD.n59 VDD.n58 0.0505
R480 VDD.n61 VDD.n60 0.0505
R481 VDD.n74 VDD.n73 0.0505
R482 VDD.n81 VDD.n80 0.0505
R483 VDD.n83 VDD.n82 0.0505
R484 VDD.n28 VDD.n5 0.0499188
R485 VDD.n49 VDD.n45 0.0470525
R486 VDD.n88 VDD.n87 0.043625
R487 VDD.n66 VDD.n65 0.043625
R488 VDD.n90 VDD.t21 0.0431131
R489 VDD.n91 VDD.t38 0.0431131
R490 VDD.n0 VDD.t1 0.0431131
R491 VDD.n11 VDD.t47 0.0431131
R492 VDD.n3 VDD.t20 0.0431131
R493 VDD.n1 VDD.t34 0.0431131
R494 VDD.n77 VDD.n6 0.038
R495 VDD.n70 VDD.n68 0.038
R496 VDD.n55 VDD.n45 0.0351875
R497 VDD.n89 VDD.n88 0.0259588
R498 VDD.n31 VDD 0.0256961
R499 VDD.n87 VDD.n86 0.0249131
R500 VDD.n85 VDD.n84 0.0249131
R501 VDD.n77 VDD.n76 0.0249131
R502 VDD.n79 VDD.n78 0.0249131
R503 VDD.n70 VDD.n69 0.0249131
R504 VDD.n72 VDD.n71 0.0249131
R505 VDD.n65 VDD.n64 0.0249131
R506 VDD.n63 VDD.n62 0.0249131
R507 VDD.n55 VDD.n54 0.0249131
R508 VDD.n57 VDD.n56 0.0249131
R509 VDD.n51 VDD.n50 0.0249131
R510 VDD.n49 VDD.n48 0.0249131
R511 VDD.n92 VDD.n91 0.0205046
R512 VDD.n94 VDD.n93 0.0205046
R513 VDD.n93 VDD.n3 0.0205046
R514 VDD.n92 VDD.n3 0.0205046
R515 VDD.n29 VDD.n28 0.0197986
R516 VDD.n48 VDD.t6 0.0187
R517 VDD.n48 VDD.t26 0.0187
R518 VDD.n50 VDD.t25 0.0187
R519 VDD.n50 VDD.t41 0.0187
R520 VDD.n84 VDD.t45 0.0187
R521 VDD.n84 VDD.t40 0.0187
R522 VDD.n86 VDD.t32 0.0187
R523 VDD.n86 VDD.t23 0.0187
R524 VDD.n7 VDD.t11 0.0187
R525 VDD.n7 VDD.t3 0.0187
R526 VDD.n78 VDD.t16 0.0187
R527 VDD.n78 VDD.t24 0.0187
R528 VDD.n76 VDD.t43 0.0187
R529 VDD.n76 VDD.t5 0.0187
R530 VDD.n75 VDD.t30 0.0187
R531 VDD.n75 VDD.t35 0.0187
R532 VDD.n71 VDD.t42 0.0187
R533 VDD.n71 VDD.t29 0.0187
R534 VDD.n69 VDD.t14 0.0187
R535 VDD.n69 VDD.t19 0.0187
R536 VDD.n10 VDD.t7 0.0187
R537 VDD.n10 VDD.t46 0.0187
R538 VDD.n62 VDD.t39 0.0187
R539 VDD.n62 VDD.t48 0.0187
R540 VDD.n64 VDD.t22 0.0187
R541 VDD.n64 VDD.t33 0.0187
R542 VDD.n46 VDD.t2 0.0187
R543 VDD.n46 VDD.t15 0.0187
R544 VDD.n56 VDD.t10 0.0187
R545 VDD.n56 VDD.t17 0.0187
R546 VDD.n54 VDD.t37 0.0187
R547 VDD.n54 VDD.t44 0.0187
R548 VDD.n53 VDD.t18 0.0187
R549 VDD.n53 VDD.t31 0.0187
R550 VDD.n47 VDD.t36 0.0187
R551 VDD.n47 VDD.t8 0.0187
R552 VDD.n9 VDD.n8 0.00883333
R553 VDD.n60 VDD.n9 0.007278
R554 VDD.n74 VDD.n9 0.00674189
R555 VDD.n82 VDD.n81 0.00478891
R556 VDD.n81 VDD.n74 0.00478891
R557 VDD.n60 VDD.n59 0.00478891
R558 VDD.n67 VDD.n44 0.00473203
R559 VDD.n67 VDD.n66 0.00406655
R560 VDD.n68 VDD.n67 0.00401084
R561 VDD.n90 VDD.n89 0.0031422
R562 VDD.n88 VDD.n6 0.00252126
R563 VDD.n68 VDD.n6 0.00252126
R564 VDD.n66 VDD.n45 0.00252126
R565 VDD.n44 VDD.n11 0.00172034
R566 VDD.n93 VDD.t9 0.00100004
R567 VDD.t9 VDD.n92 0.00100004
R568 x1.PLUS.n0 x1.PLUS.t2 53.5367
R569 x1.PLUS.n1 x1.PLUS.t1 13.9911
R570 x1.PLUS x1.PLUS.t0 10.2104
R571 x1.PLUS.n0 x1.PLUS 0.0481471
R572 x1.PLUS.n1 x1.PLUS.n0 0.0140678
R573 x1.PLUS x1.PLUS.n1 0.00592714
R574 VSS.t58 VSS.t0 115295
R575 VSS.t0 VSS.t2 14065
R576 VSS.t2 VSS.t13 14065
R577 VSS.n264 VSS.t13 7182.67
R578 VSS.n261 VSS.n259 383.183
R579 VSS.n259 VSS.t6 353.707
R580 VSS.n255 VSS.t6 353.707
R581 VSS.n255 VSS.t80 353.707
R582 VSS.t77 VSS.n263 328.077
R583 VSS.n263 VSS.t75 328.077
R584 VSS.t75 VSS.n261 328.077
R585 VSS.n264 VSS.t77 327.49
R586 VSS.n165 VSS.n85 324.418
R587 VSS.n163 VSS.n76 324.418
R588 VSS.n179 VSS.n72 324.418
R589 VSS.n177 VSS.n63 324.418
R590 VSS.n192 VSS.n60 324.418
R591 VSS.n190 VSS.n51 324.418
R592 VSS.n206 VSS.n47 324.418
R593 VSS.n204 VSS.n38 324.418
R594 VSS.n219 VSS.n35 324.418
R595 VSS.n217 VSS.n28 324.418
R596 VSS.n249 VSS.t25 322.483
R597 VSS.n153 VSS.t44 322.084
R598 VSS.t44 VSS.n85 322.084
R599 VSS.t66 VSS.n163 322.084
R600 VSS.t5 VSS.n72 322.084
R601 VSS.t15 VSS.n177 322.084
R602 VSS.t50 VSS.n60 322.084
R603 VSS.t74 VSS.n190 322.084
R604 VSS.t32 VSS.n47 322.084
R605 VSS.t26 VSS.n204 322.084
R606 VSS.t73 VSS.n35 322.084
R607 VSS.t4 VSS.n217 322.084
R608 VSS.t19 VSS.n17 322.084
R609 VSS.n254 VSS.n17 310.413
R610 VSS.n278 VSS.n8 306.639
R611 VSS.n257 VSS.n11 303.723
R612 VSS.n244 VSS.n243 270.084
R613 VSS.n244 VSS.n7 270.084
R614 VSS.t30 VSS.t66 259.067
R615 VSS.t49 VSS.t5 259.067
R616 VSS.t24 VSS.t15 259.067
R617 VSS.t31 VSS.t50 259.067
R618 VSS.t27 VSS.t74 259.067
R619 VSS.t33 VSS.t32 259.067
R620 VSS.t56 VSS.t26 259.067
R621 VSS.t9 VSS.t73 259.067
R622 VSS.t10 VSS.t4 259.067
R623 VSS.t8 VSS.t19 259.067
R624 VSS.t25 VSS.t79 259.067
R625 VSS.n165 VSS.n164 193.716
R626 VSS.n172 VSS.n76 193.716
R627 VSS.n179 VSS.n178 193.716
R628 VSS.n186 VSS.n63 193.716
R629 VSS.n192 VSS.n191 193.716
R630 VSS.n199 VSS.n51 193.716
R631 VSS.n206 VSS.n205 193.716
R632 VSS.n213 VSS.n38 193.716
R633 VSS.n219 VSS.n218 193.716
R634 VSS.n226 VSS.n28 193.716
R635 VSS.n253 VSS.n18 193.716
R636 VSS.n154 VSS.n152 182.389
R637 VSS.n82 VSS.n81 182.389
R638 VSS.n171 VSS.n77 182.389
R639 VSS.n69 VSS.n68 182.389
R640 VSS.n185 VSS.n64 182.389
R641 VSS.n57 VSS.n56 182.389
R642 VSS.n198 VSS.n52 182.389
R643 VSS.n44 VSS.n43 182.389
R644 VSS.n212 VSS.n39 182.389
R645 VSS.n32 VSS.n31 182.389
R646 VSS.n225 VSS.n22 182.389
R647 VSS.n250 VSS.n249 182.389
R648 VSS.n258 VSS.n257 176.362
R649 VSS.n258 VSS.n8 176.362
R650 VSS.n240 VSS.n231 176.362
R651 VSS.n232 VSS.n231 176.362
R652 VSS.n153 VSS.t58 170.377
R653 VSS.n265 VSS.n15 161.779
R654 VSS.n260 VSS.n15 161.779
R655 VSS.n260 VSS.n16 161.779
R656 VSS.n265 VSS.n16 161.779
R657 VSS.t28 VSS.n231 132.171
R658 VSS.n244 VSS.t11 132.082
R659 VSS.n238 VSS.t28 131.97
R660 VSS.n238 VSS.t57 131.97
R661 VSS.n276 VSS.t11 131.97
R662 VSS.n257 VSS.n256 122.695
R663 VSS.n256 VSS.n8 122.695
R664 VSS.n240 VSS.n239 122.695
R665 VSS.n239 VSS.n232 122.695
R666 VSS.n278 VSS.n7 121.603
R667 VSS.n262 VSS.n15 112.001
R668 VSS.n262 VSS.n16 112.001
R669 VSS.n248 VSS.n23 95.0838
R670 VSS.n243 VSS.n240 93.962
R671 VSS.n275 VSS.n11 88.5474
R672 VSS.t80 VSS.n254 79.7444
R673 VSS.n161 VSS.n160 67.8616
R674 VSS.n154 VSS.n149 64.3616
R675 VSS.n167 VSS.n82 64.3616
R676 VSS.n168 VSS.n81 64.3616
R677 VSS.n171 VSS.n78 64.3616
R678 VSS.n77 VSS.n70 64.3616
R679 VSS.n181 VSS.n69 64.3616
R680 VSS.n182 VSS.n68 64.3616
R681 VSS.n185 VSS.n65 64.3616
R682 VSS.n64 VSS.n58 64.3616
R683 VSS.n194 VSS.n57 64.3616
R684 VSS.n195 VSS.n56 64.3616
R685 VSS.n198 VSS.n53 64.3616
R686 VSS.n52 VSS.n45 64.3616
R687 VSS.n208 VSS.n44 64.3616
R688 VSS.n209 VSS.n43 64.3616
R689 VSS.n212 VSS.n40 64.3616
R690 VSS.n39 VSS.n33 64.3616
R691 VSS.n221 VSS.n32 64.3616
R692 VSS.n222 VSS.n31 64.3616
R693 VSS.n225 VSS.n29 64.3616
R694 VSS.n22 VSS.n19 64.3616
R695 VSS.n250 VSS.n20 64.3616
R696 VSS.n249 VSS.n23 64.3616
R697 VSS.n152 VSS.n83 64.3616
R698 VSS.n164 VSS.t30 63.0167
R699 VSS.t49 VSS.n172 63.0167
R700 VSS.n178 VSS.t24 63.0167
R701 VSS.t31 VSS.n186 63.0167
R702 VSS.n191 VSS.t27 63.0167
R703 VSS.t33 VSS.n199 63.0167
R704 VSS.n205 VSS.t56 63.0167
R705 VSS.t9 VSS.n213 63.0167
R706 VSS.n218 VSS.t10 63.0167
R707 VSS.t8 VSS.n226 63.0167
R708 VSS.t79 VSS.n18 63.0167
R709 VSS.n277 VSS.n276 62.6384
R710 VSS.n149 VSS.n83 53.6672
R711 VSS.n168 VSS.n167 53.6672
R712 VSS.n78 VSS.n70 53.6672
R713 VSS.n182 VSS.n181 53.6672
R714 VSS.n65 VSS.n58 53.6672
R715 VSS.n195 VSS.n194 53.6672
R716 VSS.n53 VSS.n45 53.6672
R717 VSS.n209 VSS.n208 53.6672
R718 VSS.n40 VSS.n33 53.6672
R719 VSS.n222 VSS.n221 53.6672
R720 VSS.n29 VSS.n19 53.6672
R721 VSS.n23 VSS.n20 53.6672
R722 VSS.n232 VSS.n10 50.1672
R723 VSS.n162 VSS.n161 48.4172
R724 VSS.n162 VSS.n75 48.4172
R725 VSS.n173 VSS.n75 48.4172
R726 VSS.n173 VSS.n73 48.4172
R727 VSS.n176 VSS.n73 48.4172
R728 VSS.n176 VSS.n61 48.4172
R729 VSS.n187 VSS.n61 48.4172
R730 VSS.n188 VSS.n187 48.4172
R731 VSS.n189 VSS.n188 48.4172
R732 VSS.n189 VSS.n50 48.4172
R733 VSS.n200 VSS.n50 48.4172
R734 VSS.n200 VSS.n48 48.4172
R735 VSS.n203 VSS.n48 48.4172
R736 VSS.n203 VSS.n36 48.4172
R737 VSS.n214 VSS.n36 48.4172
R738 VSS.n215 VSS.n214 48.4172
R739 VSS.n216 VSS.n215 48.4172
R740 VSS.n216 VSS.n27 48.4172
R741 VSS.n227 VSS.n27 48.4172
R742 VSS.n227 VSS.n25 48.4172
R743 VSS.n248 VSS.n25 48.4172
R744 VSS.n11 VSS.n7 47.035
R745 VSS.n161 VSS.n83 46.6672
R746 VSS.n168 VSS.n75 46.6672
R747 VSS.n73 VSS.n70 46.6672
R748 VSS.n182 VSS.n61 46.6672
R749 VSS.n188 VSS.n58 46.6672
R750 VSS.n195 VSS.n50 46.6672
R751 VSS.n48 VSS.n45 46.6672
R752 VSS.n209 VSS.n36 46.6672
R753 VSS.n215 VSS.n33 46.6672
R754 VSS.n222 VSS.n27 46.6672
R755 VSS.n25 VSS.n19 46.6672
R756 VSS.n242 VSS.n10 43.6832
R757 VSS.n128 VSS.n126 34.1162
R758 VSS.n142 VSS.n140 34.1096
R759 VSS.n134 VSS.n132 34.1096
R760 VSS.n120 VSS.n118 34.1085
R761 VSS.n107 VSS.n105 34.1074
R762 VSS.n113 VSS.n111 34.1063
R763 VSS.n243 VSS.n242 27.7313
R764 VSS.n166 VSS.n83 27.0283
R765 VSS.n169 VSS.n168 27.0283
R766 VSS.n180 VSS.n70 27.0283
R767 VSS.n183 VSS.n182 27.0283
R768 VSS.n193 VSS.n58 27.0283
R769 VSS.n196 VSS.n195 27.0283
R770 VSS.n207 VSS.n45 27.0283
R771 VSS.n210 VSS.n209 27.0283
R772 VSS.n220 VSS.n33 27.0283
R773 VSS.n223 VSS.n222 27.0283
R774 VSS.n252 VSS.n19 27.0283
R775 VSS.n129 VSS.n124 25.6892
R776 VSS.n121 VSS.n116 25.6794
R777 VSS.n103 VSS.n102 25.6774
R778 VSS.n114 VSS.n94 25.6774
R779 VSS.n138 VSS.n92 25.6755
R780 VSS.n135 VSS.n130 25.6559
R781 VSS.n254 VSS.n9 20.0829
R782 VSS.n167 VSS.n166 16.1394
R783 VSS.n169 VSS.n78 16.1394
R784 VSS.n181 VSS.n180 16.1394
R785 VSS.n183 VSS.n65 16.1394
R786 VSS.n194 VSS.n193 16.1394
R787 VSS.n196 VSS.n53 16.1394
R788 VSS.n208 VSS.n207 16.1394
R789 VSS.n210 VSS.n40 16.1394
R790 VSS.n221 VSS.n220 16.1394
R791 VSS.n223 VSS.n29 16.1394
R792 VSS.n252 VSS.n20 16.1394
R793 VSS.n275 VSS.n10 14.8231
R794 VSS.n158 VSS.n149 14.1949
R795 VSS.n254 VSS.n253 14.0041
R796 VSS.n96 VSS.n88 7.83243
R797 VSS.n156 VSS.t59 7.26669
R798 VSS.n281 VSS.t7 7.24741
R799 VSS.n235 VSS.t29 7.23685
R800 VSS.n88 VSS.n0 6.85872
R801 VSS.n135 VSS.n134 6.58153
R802 VSS.n140 VSS.n138 6.56196
R803 VSS.n105 VSS.n103 6.56001
R804 VSS.n114 VSS.n113 6.56001
R805 VSS.n121 VSS.n120 6.55805
R806 VSS.n129 VSS.n128 6.54827
R807 VSS.n273 VSS.n272 6.18898
R808 VSS.n100 VSS.n99 5.95109
R809 VSS.n98 VSS.n97 4.41109
R810 VSS.n284 VSS.n1 4.3205
R811 VSS.n101 VSS.n14 4.01281
R812 VSS.n97 VSS.n96 4.0018
R813 VSS.n271 VSS.n13 3.76189
R814 VSS.n234 VSS.n233 3.57507
R815 VSS.n147 VSS.n146 3.08674
R816 VSS.n230 VSS 2.63091
R817 VSS.n233 VSS.n13 2.60463
R818 VSS.n283 VSS.n282 2.58942
R819 VSS.n237 VSS.n234 2.49507
R820 VSS.n237 VSS.n236 2.49507
R821 VSS.n272 VSS.n5 2.49507
R822 VSS.n280 VSS.n5 2.49507
R823 VSS.t80 VSS.t57 2.39126
R824 VSS.n277 VSS.n9 2.39126
R825 VSS.n95 VSS.n89 2.28848
R826 VSS.n269 VSS.n3 2.22115
R827 VSS.n268 VSS.n267 1.62406
R828 VSS.n99 VSS.n98 1.5405
R829 VSS.n96 VSS.n95 1.52562
R830 VSS.n145 VSS.n14 1.52318
R831 VSS.n170 VSS.n169 1.4287
R832 VSS.n180 VSS.n71 1.4287
R833 VSS.n184 VSS.n183 1.4287
R834 VSS.n193 VSS.n59 1.4287
R835 VSS.n197 VSS.n196 1.4287
R836 VSS.n207 VSS.n46 1.4287
R837 VSS.n211 VSS.n210 1.4287
R838 VSS.n220 VSS.n34 1.4287
R839 VSS.n224 VSS.n223 1.4287
R840 VSS.n252 VSS.n251 1.4287
R841 VSS.n253 VSS.n252 1.3005
R842 VSS.n223 VSS.n28 1.3005
R843 VSS.n220 VSS.n219 1.3005
R844 VSS.n210 VSS.n38 1.3005
R845 VSS.n207 VSS.n206 1.3005
R846 VSS.n196 VSS.n51 1.3005
R847 VSS.n193 VSS.n192 1.3005
R848 VSS.n183 VSS.n63 1.3005
R849 VSS.n180 VSS.n179 1.3005
R850 VSS.n169 VSS.n76 1.3005
R851 VSS.n166 VSS.n84 1.3005
R852 VSS.n166 VSS.n165 1.3005
R853 VSS.n269 VSS.n268 1.06093
R854 VSS.n234 VSS.n229 1.05125
R855 VSS.n236 VSS.n12 1.0355
R856 VSS.n284 VSS.n283 1.01317
R857 VSS.n157 VSS.n84 0.9905
R858 VSS.n272 VSS.n271 0.892674
R859 VSS.n147 VSS.n89 0.798754
R860 VSS.n280 VSS.n279 0.739638
R861 VSS.n273 VSS.n6 0.682364
R862 VSS.n24 VSS.n21 0.653052
R863 VSS.n241 VSS.n12 0.642368
R864 VSS.n274 VSS.n273 0.615063
R865 VSS.n268 VSS.n2 0.596161
R866 VSS.n283 VSS.n2 0.596161
R867 VSS.n248 VSS.n247 0.578278
R868 VSS.t79 VSS.n248 0.578278
R869 VSS.n228 VSS.n227 0.578278
R870 VSS.n227 VSS.t8 0.578278
R871 VSS.n216 VSS.n26 0.578278
R872 VSS.t10 VSS.n216 0.578278
R873 VSS.n214 VSS.n37 0.578278
R874 VSS.n214 VSS.t9 0.578278
R875 VSS.n203 VSS.n202 0.578278
R876 VSS.t56 VSS.n203 0.578278
R877 VSS.n201 VSS.n200 0.578278
R878 VSS.n200 VSS.t33 0.578278
R879 VSS.n189 VSS.n49 0.578278
R880 VSS.t27 VSS.n189 0.578278
R881 VSS.n187 VSS.n62 0.578278
R882 VSS.n187 VSS.t31 0.578278
R883 VSS.n176 VSS.n175 0.578278
R884 VSS.t24 VSS.n176 0.578278
R885 VSS.n174 VSS.n173 0.578278
R886 VSS.n173 VSS.t49 0.578278
R887 VSS.n162 VSS.n74 0.578278
R888 VSS.t30 VSS.n162 0.578278
R889 VSS.n155 VSS.n150 0.564407
R890 VSS.n246 VSS.n245 0.53773
R891 VSS.n86 VSS.n74 0.518
R892 VSS.n150 VSS.n80 0.50094
R893 VSS.n80 VSS.n79 0.50094
R894 VSS.n79 VSS.n67 0.50094
R895 VSS.n67 VSS.n66 0.50094
R896 VSS.n66 VSS.n55 0.50094
R897 VSS.n55 VSS.n54 0.50094
R898 VSS.n54 VSS.n42 0.50094
R899 VSS.n42 VSS.n41 0.50094
R900 VSS.n41 VSS.n30 0.50094
R901 VSS.n30 VSS.n21 0.50094
R902 VSS.n282 VSS.n281 0.49092
R903 VSS.n2 VSS.t76 0.4643
R904 VSS.n2 VSS.t78 0.4643
R905 VSS.n1 VSS.n0 0.459071
R906 VSS.n267 VSS.n266 0.447421
R907 VSS.n230 VSS.n6 0.434866
R908 VSS.n174 VSS.n74 0.431462
R909 VSS.n175 VSS.n174 0.431462
R910 VSS.n175 VSS.n62 0.431462
R911 VSS.n62 VSS.n49 0.431462
R912 VSS.n201 VSS.n49 0.431462
R913 VSS.n202 VSS.n201 0.431462
R914 VSS.n202 VSS.n37 0.431462
R915 VSS.n37 VSS.n26 0.431462
R916 VSS.n228 VSS.n26 0.431462
R917 VSS.n156 VSS.n86 0.409458
R918 VSS.n152 VSS.n151 0.4005
R919 VSS.n152 VSS.n85 0.4005
R920 VSS.n155 VSS.n154 0.4005
R921 VSS.n154 VSS.n153 0.4005
R922 VSS.n170 VSS.n81 0.4005
R923 VSS.n163 VSS.n81 0.4005
R924 VSS.n151 VSS.n82 0.4005
R925 VSS.n164 VSS.n82 0.4005
R926 VSS.n77 VSS.n71 0.4005
R927 VSS.n77 VSS.n72 0.4005
R928 VSS.n171 VSS.n170 0.4005
R929 VSS.n172 VSS.n171 0.4005
R930 VSS.n184 VSS.n68 0.4005
R931 VSS.n177 VSS.n68 0.4005
R932 VSS.n71 VSS.n69 0.4005
R933 VSS.n178 VSS.n69 0.4005
R934 VSS.n64 VSS.n59 0.4005
R935 VSS.n64 VSS.n60 0.4005
R936 VSS.n185 VSS.n184 0.4005
R937 VSS.n186 VSS.n185 0.4005
R938 VSS.n197 VSS.n56 0.4005
R939 VSS.n190 VSS.n56 0.4005
R940 VSS.n59 VSS.n57 0.4005
R941 VSS.n191 VSS.n57 0.4005
R942 VSS.n52 VSS.n46 0.4005
R943 VSS.n52 VSS.n47 0.4005
R944 VSS.n198 VSS.n197 0.4005
R945 VSS.n199 VSS.n198 0.4005
R946 VSS.n211 VSS.n43 0.4005
R947 VSS.n204 VSS.n43 0.4005
R948 VSS.n46 VSS.n44 0.4005
R949 VSS.n205 VSS.n44 0.4005
R950 VSS.n39 VSS.n34 0.4005
R951 VSS.n39 VSS.n35 0.4005
R952 VSS.n212 VSS.n211 0.4005
R953 VSS.n213 VSS.n212 0.4005
R954 VSS.n224 VSS.n31 0.4005
R955 VSS.n217 VSS.n31 0.4005
R956 VSS.n34 VSS.n32 0.4005
R957 VSS.n218 VSS.n32 0.4005
R958 VSS.n251 VSS.n22 0.4005
R959 VSS.n22 VSS.n17 0.4005
R960 VSS.n225 VSS.n224 0.4005
R961 VSS.n226 VSS.n225 0.4005
R962 VSS.n251 VSS.n250 0.4005
R963 VSS.n250 VSS.n18 0.4005
R964 VSS.n158 VSS.n157 0.4005
R965 VSS.n160 VSS.n86 0.4005
R966 VSS.n249 VSS.n24 0.4005
R967 VSS.n159 VSS.n158 0.399253
R968 VSS.n160 VSS.n159 0.399253
R969 VSS.n241 VSS.n229 0.396599
R970 VSS.n247 VSS.n228 0.380594
R971 VSS.n236 VSS.n235 0.348761
R972 VSS.n246 VSS.n24 0.30829
R973 VSS.n270 VSS.n4 0.291269
R974 VSS.n235 VSS.n13 0.239196
R975 VSS.n271 VSS.n270 0.234543
R976 VSS.n266 VSS.n265 0.218565
R977 VSS.n265 VSS.n264 0.217167
R978 VSS.n262 VSS.n2 0.217167
R979 VSS.n263 VSS.n262 0.217167
R980 VSS.n260 VSS.n3 0.217167
R981 VSS.n261 VSS.n260 0.217167
R982 VSS.n282 VSS.n3 0.207891
R983 VSS.n233 VSS.n231 0.2005
R984 VSS.n239 VSS.n237 0.2005
R985 VSS.n239 VSS.n238 0.2005
R986 VSS.n242 VSS.n241 0.2005
R987 VSS.n242 VSS.n9 0.2005
R988 VSS.n258 VSS.n4 0.2005
R989 VSS.n259 VSS.n258 0.2005
R990 VSS.n256 VSS.n5 0.2005
R991 VSS.n256 VSS.n255 0.2005
R992 VSS.n281 VSS.n280 0.176544
R993 VSS.n151 VSS.n150 0.132745
R994 VSS.n170 VSS.n80 0.132745
R995 VSS.n79 VSS.n71 0.132745
R996 VSS.n184 VSS.n67 0.132745
R997 VSS.n66 VSS.n59 0.132745
R998 VSS.n197 VSS.n55 0.132745
R999 VSS.n54 VSS.n46 0.132745
R1000 VSS.n211 VSS.n42 0.132745
R1001 VSS.n41 VSS.n34 0.132745
R1002 VSS.n224 VSS.n30 0.132745
R1003 VSS.n251 VSS.n21 0.132745
R1004 VSS.n151 VSS.n84 0.128704
R1005 VSS.n274 VSS.n12 0.113124
R1006 VSS.n275 VSS.n274 0.111138
R1007 VSS.n276 VSS.n275 0.111138
R1008 VSS.n245 VSS.n244 0.111138
R1009 VSS.n279 VSS.n6 0.105757
R1010 VSS.n279 VSS.n278 0.0967963
R1011 VSS.n278 VSS.n277 0.0967963
R1012 VSS.n270 VSS.n269 0.089904
R1013 VSS.n246 VSS.n229 0.0840962
R1014 VSS.n157 VSS.n156 0.081341
R1015 VSS.n157 VSS.n155 0.0620279
R1016 VSS.n282 VSS.n4 0.0607007
R1017 VSS.n126 VSS.n91 0.0597094
R1018 VSS.n98 VSS.n93 0.0547889
R1019 VSS.n136 VSS.n129 0.0547889
R1020 VSS.n247 VSS.n246 0.0541139
R1021 VSS.n136 VSS.n135 0.0505
R1022 VSS.n138 VSS.n137 0.0505
R1023 VSS.n122 VSS.n121 0.0505
R1024 VSS.n115 VSS.n114 0.0505
R1025 VSS.n103 VSS.n93 0.0505
R1026 VSS.n245 VSS.n230 0.0467676
R1027 VSS.n100 VSS.t20 0.0464575
R1028 VSS.n99 VSS.t71 0.0464575
R1029 VSS.n97 VSS.t1 0.0464575
R1030 VSS.n146 VSS.t67 0.0464575
R1031 VSS.n147 VSS.t3 0.0464575
R1032 VSS.n95 VSS.t23 0.0464575
R1033 VSS.n143 VSS.n142 0.043625
R1034 VSS.n132 VSS.n91 0.043625
R1035 VSS.n118 VSS.n90 0.0422188
R1036 VSS.n108 VSS.n107 0.0408125
R1037 VSS.n111 VSS.n109 0.039529
R1038 VSS.n105 VSS.n104 0.0300775
R1039 VSS.n107 VSS.n106 0.0300775
R1040 VSS.n113 VSS.n112 0.0300775
R1041 VSS.n111 VSS.n110 0.0300775
R1042 VSS.n120 VSS.n119 0.0300775
R1043 VSS.n118 VSS.n117 0.0300775
R1044 VSS.n140 VSS.n139 0.0300775
R1045 VSS.n142 VSS.n141 0.0300775
R1046 VSS.n134 VSS.n133 0.0300775
R1047 VSS.n132 VSS.n131 0.0300775
R1048 VSS.n126 VSS.n125 0.0300775
R1049 VSS.n128 VSS.n127 0.0300775
R1050 VSS.n108 VSS.n101 0.0259594
R1051 VSS.n267 VSS.n14 0.0238731
R1052 VSS.n148 VSS.n147 0.017599
R1053 VSS.n148 VSS.n88 0.017599
R1054 VSS.n99 VSS.n87 0.017099
R1055 VSS.n147 VSS.n87 0.017099
R1056 VSS.n127 VSS.t46 0.01688
R1057 VSS.n127 VSS.t36 0.01688
R1058 VSS.n125 VSS.t54 0.01688
R1059 VSS.n125 VSS.t65 0.01688
R1060 VSS.n106 VSS.t62 0.01688
R1061 VSS.n106 VSS.t47 0.01688
R1062 VSS.n104 VSS.t17 0.01688
R1063 VSS.n104 VSS.t60 0.01688
R1064 VSS.n102 VSS.t52 0.01688
R1065 VSS.n102 VSS.t69 0.01688
R1066 VSS.n110 VSS.t43 0.01688
R1067 VSS.n110 VSS.t14 0.01688
R1068 VSS.n112 VSS.t39 0.01688
R1069 VSS.n112 VSS.t48 0.01688
R1070 VSS.n94 VSS.t41 0.01688
R1071 VSS.n94 VSS.t16 0.01688
R1072 VSS.n117 VSS.t22 0.01688
R1073 VSS.n117 VSS.t55 0.01688
R1074 VSS.n119 VSS.t64 0.01688
R1075 VSS.n119 VSS.t61 0.01688
R1076 VSS.n116 VSS.t12 0.01688
R1077 VSS.n116 VSS.t45 0.01688
R1078 VSS.n141 VSS.t18 0.01688
R1079 VSS.n141 VSS.t37 0.01688
R1080 VSS.n139 VSS.t42 0.01688
R1081 VSS.n139 VSS.t68 0.01688
R1082 VSS.n92 VSS.t21 0.01688
R1083 VSS.n92 VSS.t51 0.01688
R1084 VSS.n131 VSS.t40 0.01688
R1085 VSS.n131 VSS.t53 0.01688
R1086 VSS.n133 VSS.t35 0.01688
R1087 VSS.n133 VSS.t38 0.01688
R1088 VSS.n130 VSS.t63 0.01688
R1089 VSS.n130 VSS.t72 0.01688
R1090 VSS.n124 VSS.t34 0.01688
R1091 VSS.n124 VSS.t70 0.01688
R1092 VSS VSS.n284 0.016025
R1093 VSS.n123 VSS.n89 0.00896236
R1094 VSS.n266 VSS.n1 0.0086575
R1095 VSS.n137 VSS.n123 0.00751474
R1096 VSS.n123 VSS.n122 0.00738071
R1097 VSS.n101 VSS.n100 0.00491176
R1098 VSS.n115 VSS.n93 0.00478891
R1099 VSS.n122 VSS.n115 0.00478891
R1100 VSS.n137 VSS.n136 0.00478891
R1101 VSS.n145 VSS.n144 0.00440625
R1102 VSS VSS.n0 0.003875
R1103 VSS.n144 VSS.n143 0.00371783
R1104 VSS.n144 VSS.n90 0.00341997
R1105 VSS.n146 VSS.n145 0.00294068
R1106 VSS.n109 VSS.n108 0.00252186
R1107 VSS.n109 VSS.n90 0.00252186
R1108 VSS.n143 VSS.n91 0.00252186
R1109 VSS.n159 VSS.t58 0.00187342
R1110 VSS.t2 VSS.n148 0.00150002
R1111 VSS.t2 VSS.n87 0.00100002
R1112 a_3162_2792.n11 a_3162_2792.t41 620.048
R1113 a_3162_2792.n13 a_3162_2792.t37 620.048
R1114 a_3162_2792.t14 a_3162_2792.n2 620.048
R1115 a_3162_2792.t23 a_3162_2792.n67 620.048
R1116 a_3162_2792.n55 a_3162_2792.t6 620.048
R1117 a_3162_2792.n36 a_3162_2792.t31 620.048
R1118 a_3162_2792.t36 a_3162_2792.n33 620.048
R1119 a_3162_2792.t20 a_3162_2792.n48 620.048
R1120 a_3162_2792.t34 a_3162_2792.n36 619.74
R1121 a_3162_2792.n33 a_3162_2792.t38 619.74
R1122 a_3162_2792.t16 a_3162_2792.n29 619.74
R1123 a_3162_2792.t25 a_3162_2792.n24 619.74
R1124 a_3162_2792.n44 a_3162_2792.t9 619.74
R1125 a_3162_2792.n62 a_3162_2792.t18 619.74
R1126 a_3162_2792.t2 a_3162_2792.n56 619.74
R1127 a_3162_2792.t8 a_3162_2792.n25 619.74
R1128 a_3162_2792.n67 a_3162_2792.t39 619.74
R1129 a_3162_2792.t35 a_3162_2792.n2 619.74
R1130 a_3162_2792.n66 a_3162_2792.t43 619.74
R1131 a_3162_2792.n77 a_3162_2792.t40 619.74
R1132 a_3162_2792.n64 a_3162_2792.t10 619.74
R1133 a_3162_2792.n78 a_3162_2792.t4 619.74
R1134 a_3162_2792.t17 a_3162_2792.n13 619.74
R1135 a_3162_2792.t26 a_3162_2792.n11 619.74
R1136 a_3162_2792.t11 a_3162_2792.n1 619.74
R1137 a_3162_2792.t19 a_3162_2792.n7 619.74
R1138 a_3162_2792.n48 a_3162_2792.t27 619.74
R1139 a_3162_2792.n55 a_3162_2792.t13 619.74
R1140 a_3162_2792.n37 a_3162_2792.t3 614.254
R1141 a_3162_2792.n37 a_3162_2792.t34 614.254
R1142 a_3162_2792.n32 a_3162_2792.t3 614.254
R1143 a_3162_2792.t38 a_3162_2792.n32 614.254
R1144 a_3162_2792.n40 a_3162_2792.t32 614.254
R1145 a_3162_2792.n40 a_3162_2792.t16 614.254
R1146 a_3162_2792.t32 a_3162_2792.n39 614.254
R1147 a_3162_2792.n39 a_3162_2792.t25 614.254
R1148 a_3162_2792.n43 a_3162_2792.t28 614.254
R1149 a_3162_2792.t9 a_3162_2792.n43 614.254
R1150 a_3162_2792.n61 a_3162_2792.t28 614.254
R1151 a_3162_2792.t18 a_3162_2792.n61 614.254
R1152 a_3162_2792.t21 a_3162_2792.n57 614.254
R1153 a_3162_2792.n57 a_3162_2792.t2 614.254
R1154 a_3162_2792.n58 a_3162_2792.t21 614.254
R1155 a_3162_2792.n58 a_3162_2792.t8 614.254
R1156 a_3162_2792.n72 a_3162_2792.t39 614.254
R1157 a_3162_2792.t5 a_3162_2792.n72 614.254
R1158 a_3162_2792.n73 a_3162_2792.t5 614.254
R1159 a_3162_2792.n73 a_3162_2792.t35 614.254
R1160 a_3162_2792.t43 a_3162_2792.n65 614.254
R1161 a_3162_2792.n65 a_3162_2792.t12 614.254
R1162 a_3162_2792.n76 a_3162_2792.t12 614.254
R1163 a_3162_2792.t40 a_3162_2792.n76 614.254
R1164 a_3162_2792.t10 a_3162_2792.n22 614.254
R1165 a_3162_2792.n22 a_3162_2792.t22 614.254
R1166 a_3162_2792.t22 a_3162_2792.n21 614.254
R1167 a_3162_2792.n21 a_3162_2792.t4 614.254
R1168 a_3162_2792.n14 a_3162_2792.t33 614.254
R1169 a_3162_2792.n14 a_3162_2792.t17 614.254
R1170 a_3162_2792.n12 a_3162_2792.t26 614.254
R1171 a_3162_2792.t33 a_3162_2792.n12 614.254
R1172 a_3162_2792.t29 a_3162_2792.n17 614.254
R1173 a_3162_2792.n17 a_3162_2792.t11 614.254
R1174 a_3162_2792.n18 a_3162_2792.t19 614.254
R1175 a_3162_2792.n18 a_3162_2792.t29 614.254
R1176 a_3162_2792.t41 a_3162_2792.n10 614.254
R1177 a_3162_2792.n10 a_3162_2792.t7 614.254
R1178 a_3162_2792.t7 a_3162_2792.n9 614.254
R1179 a_3162_2792.t37 a_3162_2792.n9 614.254
R1180 a_3162_2792.t30 a_3162_2792.n68 614.254
R1181 a_3162_2792.n68 a_3162_2792.t14 614.254
R1182 a_3162_2792.n69 a_3162_2792.t23 614.254
R1183 a_3162_2792.n69 a_3162_2792.t30 614.254
R1184 a_3162_2792.t27 a_3162_2792.n47 614.254
R1185 a_3162_2792.n47 a_3162_2792.t24 614.254
R1186 a_3162_2792.n54 a_3162_2792.t24 614.254
R1187 a_3162_2792.t13 a_3162_2792.n54 614.254
R1188 a_3162_2792.n51 a_3162_2792.t6 614.254
R1189 a_3162_2792.n35 a_3162_2792.t42 614.254
R1190 a_3162_2792.t31 a_3162_2792.n35 614.254
R1191 a_3162_2792.t42 a_3162_2792.n34 614.254
R1192 a_3162_2792.n34 a_3162_2792.t36 614.254
R1193 a_3162_2792.n50 a_3162_2792.t20 614.254
R1194 a_3162_2792.t15 a_3162_2792.n50 614.254
R1195 a_3162_2792.n51 a_3162_2792.t15 614.254
R1196 a_3162_2792.n63 a_3162_2792.n23 15.7039
R1197 a_3162_2792.n46 a_3162_2792.n45 15.3876
R1198 a_3162_2792.n46 a_3162_2792.n23 14.6668
R1199 a_3162_2792.n15 a_3162_2792.n9 5.13335
R1200 a_3162_2792.n10 a_3162_2792.n8 5.13335
R1201 a_3162_2792.n35 a_3162_2792.n30 5.02611
R1202 a_3162_2792.n54 a_3162_2792.n53 5.02611
R1203 a_3162_2792.n34 a_3162_2792.n6 5.02611
R1204 a_3162_2792.n38 a_3162_2792.n37 5.02611
R1205 a_3162_2792.n32 a_3162_2792.n31 5.02611
R1206 a_3162_2792.n41 a_3162_2792.n40 5.02611
R1207 a_3162_2792.n39 a_3162_2792.n26 5.02611
R1208 a_3162_2792.n43 a_3162_2792.n42 5.02611
R1209 a_3162_2792.n61 a_3162_2792.n60 5.02611
R1210 a_3162_2792.n57 a_3162_2792.n28 5.02611
R1211 a_3162_2792.n59 a_3162_2792.n58 5.02611
R1212 a_3162_2792.n50 a_3162_2792.n49 5.02611
R1213 a_3162_2792.n70 a_3162_2792.n69 5.02611
R1214 a_3162_2792.n68 a_3162_2792.n4 5.02611
R1215 a_3162_2792.n74 a_3162_2792.n73 5.02611
R1216 a_3162_2792.n72 a_3162_2792.n71 5.02611
R1217 a_3162_2792.n76 a_3162_2792.n75 5.02611
R1218 a_3162_2792.n65 a_3162_2792.n5 5.02611
R1219 a_3162_2792.n21 a_3162_2792.n3 5.02611
R1220 a_3162_2792.n22 a_3162_2792.n20 5.02611
R1221 a_3162_2792.n12 a_3162_2792.n8 5.02611
R1222 a_3162_2792.n15 a_3162_2792.n14 5.02611
R1223 a_3162_2792.n19 a_3162_2792.n18 5.02611
R1224 a_3162_2792.n17 a_3162_2792.n16 5.02611
R1225 a_3162_2792.n47 a_3162_2792.n27 5.02611
R1226 a_3162_2792.n52 a_3162_2792.n51 5.02611
R1227 a_3162_2792.n64 a_3162_2792.n63 2.8286
R1228 a_3162_2792.n79 a_3162_2792.n0 1.12638
R1229 a_3162_2792.n0 a_3162_2792.t1 1.04563
R1230 a_3162_2792.t0 a_3162_2792.n79 0.96115
R1231 a_3162_2792.n70 a_3162_2792.n6 0.437096
R1232 a_3162_2792.n30 a_3162_2792.n4 0.437096
R1233 a_3162_2792.n63 a_3162_2792.n62 0.321929
R1234 a_3162_2792.n45 a_3162_2792.n44 0.321929
R1235 a_3162_2792.n79 a_3162_2792.n78 0.321929
R1236 a_3162_2792.n64 a_3162_2792.n7 0.308818
R1237 a_3162_2792.n11 a_3162_2792.n7 0.308818
R1238 a_3162_2792.n13 a_3162_2792.n1 0.308818
R1239 a_3162_2792.n78 a_3162_2792.n1 0.308818
R1240 a_3162_2792.n78 a_3162_2792.n77 0.308818
R1241 a_3162_2792.n77 a_3162_2792.n2 0.308818
R1242 a_3162_2792.n67 a_3162_2792.n66 0.308818
R1243 a_3162_2792.n66 a_3162_2792.n64 0.308818
R1244 a_3162_2792.n56 a_3162_2792.n55 0.308818
R1245 a_3162_2792.n56 a_3162_2792.n44 0.308818
R1246 a_3162_2792.n44 a_3162_2792.n29 0.308818
R1247 a_3162_2792.n36 a_3162_2792.n29 0.308818
R1248 a_3162_2792.n33 a_3162_2792.n24 0.308818
R1249 a_3162_2792.n62 a_3162_2792.n24 0.308818
R1250 a_3162_2792.n62 a_3162_2792.n25 0.308818
R1251 a_3162_2792.n48 a_3162_2792.n25 0.308818
R1252 a_3162_2792.n45 a_3162_2792.n0 0.157817
R1253 a_3162_2792.n49 a_3162_2792.n23 0.130713
R1254 a_3162_2792.n52 a_3162_2792.n46 0.130713
R1255 a_3162_2792.n19 a_3162_2792.n8 0.107734
R1256 a_3162_2792.n20 a_3162_2792.n19 0.107734
R1257 a_3162_2792.n20 a_3162_2792.n5 0.107734
R1258 a_3162_2792.n71 a_3162_2792.n5 0.107734
R1259 a_3162_2792.n71 a_3162_2792.n70 0.107734
R1260 a_3162_2792.n31 a_3162_2792.n6 0.107734
R1261 a_3162_2792.n31 a_3162_2792.n26 0.107734
R1262 a_3162_2792.n60 a_3162_2792.n26 0.107734
R1263 a_3162_2792.n60 a_3162_2792.n59 0.107734
R1264 a_3162_2792.n59 a_3162_2792.n27 0.107734
R1265 a_3162_2792.n49 a_3162_2792.n27 0.107734
R1266 a_3162_2792.n16 a_3162_2792.n15 0.107734
R1267 a_3162_2792.n16 a_3162_2792.n3 0.107734
R1268 a_3162_2792.n75 a_3162_2792.n3 0.107734
R1269 a_3162_2792.n75 a_3162_2792.n74 0.107734
R1270 a_3162_2792.n74 a_3162_2792.n4 0.107734
R1271 a_3162_2792.n38 a_3162_2792.n30 0.107734
R1272 a_3162_2792.n41 a_3162_2792.n38 0.107734
R1273 a_3162_2792.n42 a_3162_2792.n41 0.107734
R1274 a_3162_2792.n42 a_3162_2792.n28 0.107734
R1275 a_3162_2792.n53 a_3162_2792.n28 0.107734
R1276 a_3162_2792.n53 a_3162_2792.n52 0.107734
R1277 D4 D4.t0 9.40368
R1278 x1.MINUS x1.MINUS.t2 50.8861
R1279 x1.MINUS.n0 x1.MINUS.t0 10.548
R1280 x1.MINUS.n0 x1.MINUS.t1 9.3904
R1281 x1.MINUS x1.MINUS.n0 0.642147
R1282 D8 D8.t0 9.40368
R1283 D7 D7.t0 9.40368
R1284 D1 D1.t0 9.40368
R1285 a_2442_2792.n0 a_2442_2792.t3 39.1381
R1286 a_2442_2792.n1 a_2442_2792.t0 36.2918
R1287 a_2442_2792.n0 a_2442_2792.t2 3.29486
R1288 a_2442_2792.n1 a_2442_2792.n0 0.643925
R1289 a_2442_2792.t1 a_2442_2792.n1 0.608291
R1290 a_2576_5968.t0 a_2576_5968.n0 3.08975
R1291 a_2576_5968.n0 a_2576_5968.t2 0.551973
R1292 a_2576_5968.n0 a_2576_5968.t1 0.545657
R1293 D11 D11.t0 9.40368
R1294 D0 D0.t0 9.40368
R1295 D3 D3.t0 9.40368
R1296 D10 D10.t0 9.40368
R1297 D2 D2.t0 9.40368
R1298 D9 D9.t0 9.40368
R1299 D6 D6.t0 9.40368
R1300 D5 D5.t0 9.40368
C0 D3 D4 0.04296f
C1 D6 a_5085_9832# 0.01074f
C2 D7 D6 0.04296f
C3 a_10065_9832# a_9069_9832# 0.02769f
C4 x1.MINUS x1.ADJ 0
C5 D8 a_3093_9832# 0.01073f
C6 VDD a_579_8278# 0.04908f
C7 D5 D4 0.04296f
C8 D7 D8 0.04296f
C9 D11 D10 0.04296f
C10 a_7077_9832# VDD 0.00899f
C11 a_9069_9832# a_8073_9832# 0.02515f
C12 a_11061_9832# VDD 0.01075f
C13 OUT a_5085_9832# 0
C14 a_2097_9832# a_579_8278# 0
C15 x1.ADJ a_3093_9832# 0.00485f
C16 OUT VDD 0.35912p
C17 a_579_8278# a_1101_9832# 0.04073f
C18 a_7077_9832# D4 0.01074f
C19 a_4089_9832# OUT 0
C20 a_6081_9832# D5 0.01074f
C21 x1.MINUS VDD 0.55678f
C22 x1.ADJ a_5085_9832# 0.00556f
C23 D3 a_8073_9832# 0.01074f
C24 D9 D8 0.04296f
C25 x1.ADJ VDD 0.10745p
C26 a_7077_9832# a_6081_9832# 0.02559f
C27 a_4089_9832# x1.ADJ 0.00556f
C28 x1.ADJ a_2097_9832# 0.00495f
C29 a_10065_9832# a_11061_9832# 0.02501f
C30 a_6081_9832# OUT 0
C31 D1 D2 0.04296f
C32 a_3093_9832# VDD 0.00806f
C33 OUT a_10065_9832# 0
C34 OUT x1.PLUS 0
C35 a_4089_9832# a_3093_9832# 0.02562f
C36 OUT a_9069_9832# 0
C37 a_6081_9832# x1.ADJ 0.00556f
C38 a_2097_9832# a_3093_9832# 0.02561f
C39 a_5085_9832# VDD 0.00899f
C40 a_7077_9832# a_8073_9832# 0.02555f
C41 x1.MINUS x1.PLUS 0.42578f
C42 a_4089_9832# a_5085_9832# 0.02558f
C43 a_4089_9832# D7 0.01074f
C44 a_10065_9832# x1.ADJ 0.00527f
C45 x1.PLUS x1.ADJ 0.01905f
C46 OUT a_8073_9832# 0
C47 a_4089_9832# VDD 0.00899f
C48 D5 D6 0.04296f
C49 x1.ADJ a_9069_9832# 0.00527f
C50 a_2097_9832# VDD 0.00461f
C51 VDD a_1101_9832# 0.00402f
C52 D0 a_11061_9832# 0.01675f
C53 x1.ADJ a_8073_9832# 0.00556f
C54 D11 a_579_8278# 0.01756f
C55 a_6081_9832# a_5085_9832# 0.02558f
C56 a_2097_9832# a_1101_9832# 0.02673f
C57 D10 a_1101_9832# 0.01077f
C58 D9 a_2097_9832# 0.01073f
C59 a_6081_9832# VDD 0.00899f
C60 D1 a_10065_9832# 0.01059f
C61 D9 D10 0.04296f
C62 D2 a_9069_9832# 0.01059f
C63 a_10065_9832# VDD 0.00899f
C64 x1.PLUS VDD 0.65789f
C65 a_9069_9832# VDD 0.00899f
C66 a_7077_9832# OUT 0
C67 OUT a_11061_9832# 0
C68 D3 D2 0.04296f
C69 a_8073_9832# VDD 0.00899f
C70 x1.ADJ a_579_8278# 0
C71 a_7077_9832# x1.ADJ 0.00556f
C72 a_11061_9832# x1.ADJ 0.0113f
C73 OUT x1.ADJ 58.5278f
C74 D1 D0 0.04296f
C75 OUT VSS 0.50973p
C76 D0 VSS 0.76613f
C77 D1 VSS 0.71867f
C78 D2 VSS 0.71867f
C79 D3 VSS 0.71867f
C80 D4 VSS 0.71867f
C81 D5 VSS 0.71867f
C82 D6 VSS 0.71867f
C83 D7 VSS 0.71867f
C84 D8 VSS 0.71867f
C85 D9 VSS 0.71867f
C86 D10 VSS 0.72562f
C87 D11 VSS 0.81129f
C88 VDD VSS 1.00675p
C89 x1.ADJ VSS 13.08234f
C90 x1.PLUS VSS 5.89767f
C91 x1.MINUS VSS 4.93227f
C92 a_11061_9832# VSS 1.47836f
C93 a_10065_9832# VSS 1.33657f
C94 a_9069_9832# VSS 1.33136f
C95 a_8073_9832# VSS 1.31747f
C96 a_7077_9832# VSS 1.31709f
C97 a_6081_9832# VSS 1.31719f
C98 a_5085_9832# VSS 1.3172f
C99 a_4089_9832# VSS 1.31717f
C100 a_3093_9832# VSS 1.31693f
C101 a_2097_9832# VSS 1.31844f
C102 a_1101_9832# VSS 1.34282f
C103 a_579_8278# VSS 2.6074f
C104 a_2576_5968.t1 VSS 1.48083f
C105 a_2576_5968.t2 VSS 1.47213f
C106 a_2576_5968.n0 VSS 6.7289f
C107 a_2576_5968.t0 VSS 2.81814f
C108 a_2442_2792.t2 VSS 1.11687f
C109 a_2442_2792.t3 VSS 0.48774f
C110 a_2442_2792.n0 VSS 1.69797f
C111 a_2442_2792.t0 VSS 0.43386f
C112 a_2442_2792.n1 VSS 1.14289f
C113 a_2442_2792.t1 VSS 0.62068f
C114 x1.MINUS.t2 VSS 1.16926f
C115 x1.MINUS.t0 VSS 0.4579f
C116 x1.MINUS.t1 VSS 0.12155f
C117 x1.MINUS.n0 VSS 1.37625f
C118 a_3162_2792.t1 VSS 0.16263f
C119 a_3162_2792.n0 VSS 0.31945f
C120 a_3162_2792.n1 VSS 0.44188f
C121 a_3162_2792.t4 VSS 0.87386f
C122 a_3162_2792.n2 VSS 0.88152f
C123 a_3162_2792.t12 VSS 0.87002f
C124 a_3162_2792.n3 VSS 0.03661f
C125 a_3162_2792.n4 VSS 0.08305f
C126 a_3162_2792.t39 VSS 0.87386f
C127 a_3162_2792.n5 VSS 0.03661f
C128 a_3162_2792.n6 VSS 0.08305f
C129 a_3162_2792.n7 VSS 0.44188f
C130 a_3162_2792.n8 VSS 0.06784f
C131 a_3162_2792.t19 VSS 0.87386f
C132 a_3162_2792.n9 VSS 0.87908f
C133 a_3162_2792.t7 VSS 0.87002f
C134 a_3162_2792.n10 VSS 0.87908f
C135 a_3162_2792.t41 VSS 0.87407f
C136 a_3162_2792.n11 VSS 0.88152f
C137 a_3162_2792.t26 VSS 0.87386f
C138 a_3162_2792.n12 VSS 0.87841f
C139 a_3162_2792.t33 VSS 0.87002f
C140 a_3162_2792.t37 VSS 0.87407f
C141 a_3162_2792.n13 VSS 0.88152f
C142 a_3162_2792.t17 VSS 0.87386f
C143 a_3162_2792.n14 VSS 0.87841f
C144 a_3162_2792.n15 VSS 0.06797f
C145 a_3162_2792.n16 VSS 0.03661f
C146 a_3162_2792.t11 VSS 0.87386f
C147 a_3162_2792.n17 VSS 0.87841f
C148 a_3162_2792.t29 VSS 0.87002f
C149 a_3162_2792.n18 VSS 0.87841f
C150 a_3162_2792.n19 VSS 0.03661f
C151 a_3162_2792.n20 VSS 0.03661f
C152 a_3162_2792.n21 VSS 0.87841f
C153 a_3162_2792.t22 VSS 0.87002f
C154 a_3162_2792.n22 VSS 0.87841f
C155 a_3162_2792.t10 VSS 0.87386f
C156 a_3162_2792.n23 VSS 1.85749f
C157 a_3162_2792.n24 VSS 0.44188f
C158 a_3162_2792.n25 VSS 0.44188f
C159 a_3162_2792.t28 VSS 0.87002f
C160 a_3162_2792.n26 VSS 0.03661f
C161 a_3162_2792.n27 VSS 0.03661f
C162 a_3162_2792.t8 VSS 0.87386f
C163 a_3162_2792.n28 VSS 0.03661f
C164 a_3162_2792.n29 VSS 0.44188f
C165 a_3162_2792.n30 VSS 0.08305f
C166 a_3162_2792.t3 VSS 0.87002f
C167 a_3162_2792.n31 VSS 0.03661f
C168 a_3162_2792.n32 VSS 0.87841f
C169 a_3162_2792.t38 VSS 0.87386f
C170 a_3162_2792.n33 VSS 0.88152f
C171 a_3162_2792.t36 VSS 0.87407f
C172 a_3162_2792.n34 VSS 0.87841f
C173 a_3162_2792.t42 VSS 0.87002f
C174 a_3162_2792.n35 VSS 0.87841f
C175 a_3162_2792.t31 VSS 0.87407f
C176 a_3162_2792.n36 VSS 0.88152f
C177 a_3162_2792.t34 VSS 0.87386f
C178 a_3162_2792.n37 VSS 0.87841f
C179 a_3162_2792.n38 VSS 0.03661f
C180 a_3162_2792.t25 VSS 0.87386f
C181 a_3162_2792.n39 VSS 0.87841f
C182 a_3162_2792.t32 VSS 0.87002f
C183 a_3162_2792.t16 VSS 0.87386f
C184 a_3162_2792.n40 VSS 0.87841f
C185 a_3162_2792.n41 VSS 0.03661f
C186 a_3162_2792.n42 VSS 0.03661f
C187 a_3162_2792.n43 VSS 0.87841f
C188 a_3162_2792.t9 VSS 0.87386f
C189 a_3162_2792.n44 VSS 0.44188f
C190 a_3162_2792.t6 VSS 0.87407f
C191 a_3162_2792.t24 VSS 0.87002f
C192 a_3162_2792.n45 VSS 0.94324f
C193 a_3162_2792.n46 VSS 1.84049f
C194 a_3162_2792.n47 VSS 0.87841f
C195 a_3162_2792.t27 VSS 0.87386f
C196 a_3162_2792.n48 VSS 0.88152f
C197 a_3162_2792.t20 VSS 0.87407f
C198 a_3162_2792.n49 VSS 0.03985f
C199 a_3162_2792.n50 VSS 0.87841f
C200 a_3162_2792.t15 VSS 0.87002f
C201 a_3162_2792.n51 VSS 0.87841f
C202 a_3162_2792.n52 VSS 0.03985f
C203 a_3162_2792.n53 VSS 0.03661f
C204 a_3162_2792.n54 VSS 0.87841f
C205 a_3162_2792.t13 VSS 0.87386f
C206 a_3162_2792.n55 VSS 0.88152f
C207 a_3162_2792.n56 VSS 0.44188f
C208 a_3162_2792.t2 VSS 0.87386f
C209 a_3162_2792.n57 VSS 0.87841f
C210 a_3162_2792.t21 VSS 0.87002f
C211 a_3162_2792.n58 VSS 0.87841f
C212 a_3162_2792.n59 VSS 0.03661f
C213 a_3162_2792.n60 VSS 0.03661f
C214 a_3162_2792.n61 VSS 0.87841f
C215 a_3162_2792.t18 VSS 0.87386f
C216 a_3162_2792.n62 VSS 0.44188f
C217 a_3162_2792.n63 VSS 0.96415f
C218 a_3162_2792.n64 VSS 0.53838f
C219 a_3162_2792.n65 VSS 0.87841f
C220 a_3162_2792.t43 VSS 0.87386f
C221 a_3162_2792.n66 VSS 0.44188f
C222 a_3162_2792.n67 VSS 0.88152f
C223 a_3162_2792.t23 VSS 0.87407f
C224 a_3162_2792.t14 VSS 0.87407f
C225 a_3162_2792.n68 VSS 0.87841f
C226 a_3162_2792.t30 VSS 0.87002f
C227 a_3162_2792.n69 VSS 0.87841f
C228 a_3162_2792.n70 VSS 0.08305f
C229 a_3162_2792.n71 VSS 0.03661f
C230 a_3162_2792.n72 VSS 0.87841f
C231 a_3162_2792.t5 VSS 0.87002f
C232 a_3162_2792.t35 VSS 0.87386f
C233 a_3162_2792.n73 VSS 0.87841f
C234 a_3162_2792.n74 VSS 0.03661f
C235 a_3162_2792.n75 VSS 0.03661f
C236 a_3162_2792.n76 VSS 0.87841f
C237 a_3162_2792.t40 VSS 0.87386f
C238 a_3162_2792.n77 VSS 0.44188f
C239 a_3162_2792.n78 VSS 0.44188f
C240 a_3162_2792.n79 VSS 0.36061f
C241 a_3162_2792.t0 VSS 0.24707f
C242 x1.PLUS.t2 VSS 0.65419f
C243 x1.PLUS.n0 VSS 1.51411f
C244 x1.PLUS.t1 VSS 0.48742f
C245 x1.PLUS.n1 VSS 1.48847f
C246 x1.PLUS.t0 VSS 0.10848f
C247 VDD.t1 VSS 1.00837f
C248 VDD.n0 VSS 6.02013f
C249 VDD.t34 VSS 1.00837f
C250 VDD.n1 VSS 6.48282f
C251 VDD.n2 VSS 2.55874f
C252 VDD.t20 VSS 1.00837f
C253 VDD.n3 VSS 10.3773f
C254 VDD.t0 VSS 78.0634f
C255 VDD.t4 VSS 58.3844f
C256 VDD.n4 VSS 4.68757f
C257 VDD.t38 VSS 1.00837f
C258 VDD.n5 VSS 2.63903f
C259 VDD.n6 VSS 7.51976f
C260 VDD.t11 VSS 0.42617f
C261 VDD.t3 VSS 0.42617f
C262 VDD.n7 VSS 1.49672f
C263 VDD.n8 VSS 4.89144f
C264 VDD.n9 VSS 5.23913f
C265 VDD.t7 VSS 0.42617f
C266 VDD.t46 VSS 0.42617f
C267 VDD.n10 VSS 1.49684f
C268 VDD.t47 VSS 1.00837f
C269 VDD.n11 VSS 5.32741f
C270 VDD.t13 VSS 0.14096f
C271 VDD.n12 VSS 0.3587f
C272 VDD.t28 VSS 0.14096f
C273 VDD.n13 VSS 0.35267f
C274 VDD.n14 VSS 0.21534f
C275 VDD.n15 VSS 0.12211f
C276 VDD.n16 VSS 0.0609f
C277 VDD.n17 VSS 0.17078f
C278 VDD.n18 VSS 0.71302f
C279 VDD.t27 VSS 0.57071f
C280 VDD.n19 VSS 0.47662f
C281 VDD.n20 VSS 0.0609f
C282 VDD.n21 VSS 0.10864f
C283 VDD.n22 VSS 0.04904f
C284 VDD.n23 VSS 0.60075f
C285 VDD.n24 VSS 0.02152f
C286 VDD.t50 VSS 0.90053f
C287 VDD.t12 VSS 0.74441f
C288 VDD.n25 VSS 20.2555f
C289 VDD.n26 VSS 0.11134f
C290 VDD.n27 VSS 0.17078f
C291 VDD.n28 VSS 0.27904f
C292 VDD.n29 VSS 0.34802f
C293 VDD.n30 VSS 0.25696f
C294 VDD.t49 VSS 0.03573f
C295 VDD.n31 VSS 0.26132f
C296 VDD.n32 VSS 0.2907f
C297 VDD.n33 VSS 1.10372f
C298 VDD.n34 VSS 0.10864f
C299 VDD.n35 VSS 0.14449f
C300 VDD.n36 VSS 0.45436f
C301 VDD.t51 VSS 0.94546f
C302 VDD.n37 VSS 0.26208f
C303 VDD.n38 VSS 0.09158f
C304 VDD.n39 VSS 0.059f
C305 VDD.n40 VSS 0.03872f
C306 VDD.n41 VSS 0.08736f
C307 VDD.n42 VSS 0.27166f
C308 VDD.n43 VSS 2.73803f
C309 VDD.n44 VSS 2.41719f
C310 VDD.n45 VSS 12.0148f
C311 VDD.t2 VSS 0.42617f
C312 VDD.t15 VSS 0.42617f
C313 VDD.n46 VSS 1.49674f
C314 VDD.t36 VSS 0.42617f
C315 VDD.t8 VSS 0.42617f
C316 VDD.n47 VSS 1.49675f
C317 VDD.t6 VSS 0.42617f
C318 VDD.t26 VSS 0.42617f
C319 VDD.n48 VSS 0.85233f
C320 VDD.n49 VSS 1.00955f
C321 VDD.t25 VSS 0.42617f
C322 VDD.t41 VSS 0.42617f
C323 VDD.n50 VSS 0.85233f
C324 VDD.n51 VSS 0.52161f
C325 VDD.n52 VSS 0.74737f
C326 VDD.t18 VSS 0.42617f
C327 VDD.t31 VSS 0.42617f
C328 VDD.n53 VSS 1.49672f
C329 VDD.t37 VSS 0.42617f
C330 VDD.t44 VSS 0.42617f
C331 VDD.n54 VSS 0.85233f
C332 VDD.n55 VSS 0.88188f
C333 VDD.t10 VSS 0.42617f
C334 VDD.t17 VSS 0.42617f
C335 VDD.n56 VSS 0.85233f
C336 VDD.n57 VSS 0.52164f
C337 VDD.n58 VSS 0.58429f
C338 VDD.n59 VSS 5.35337f
C339 VDD.n60 VSS 4.45326f
C340 VDD.n61 VSS 0.58426f
C341 VDD.t39 VSS 0.42617f
C342 VDD.t48 VSS 0.42617f
C343 VDD.n62 VSS 0.85233f
C344 VDD.n63 VSS 0.52161f
C345 VDD.t22 VSS 0.42617f
C346 VDD.t33 VSS 0.42617f
C347 VDD.n64 VSS 0.85233f
C348 VDD.n65 VSS 0.81323f
C349 VDD.n66 VSS 10.1797f
C350 VDD.n67 VSS 9.3727f
C351 VDD.n68 VSS 10.4395f
C352 VDD.t14 VSS 0.42617f
C353 VDD.t19 VSS 0.42617f
C354 VDD.n69 VSS 0.85233f
C355 VDD.n70 VSS 0.85556f
C356 VDD.t42 VSS 0.42617f
C357 VDD.t29 VSS 0.42617f
C358 VDD.n71 VSS 0.85233f
C359 VDD.n72 VSS 0.52166f
C360 VDD.n73 VSS 0.58413f
C361 VDD.n74 VSS 4.23753f
C362 VDD.t30 VSS 0.42617f
C363 VDD.t35 VSS 0.42617f
C364 VDD.n75 VSS 1.49677f
C365 VDD.t43 VSS 0.42617f
C366 VDD.t5 VSS 0.42617f
C367 VDD.n76 VSS 0.85233f
C368 VDD.n77 VSS 0.85556f
C369 VDD.t16 VSS 0.42617f
C370 VDD.t24 VSS 0.42617f
C371 VDD.n78 VSS 0.85233f
C372 VDD.n79 VSS 0.52164f
C373 VDD.n80 VSS 0.58422f
C374 VDD.n81 VSS 3.45166f
C375 VDD.n82 VSS 5.42433f
C376 VDD.n83 VSS 0.58429f
C377 VDD.t45 VSS 0.42617f
C378 VDD.t40 VSS 0.42617f
C379 VDD.n84 VSS 0.85233f
C380 VDD.n85 VSS 0.52161f
C381 VDD.t32 VSS 0.42617f
C382 VDD.t23 VSS 0.42617f
C383 VDD.n86 VSS 0.85233f
C384 VDD.n87 VSS 0.81323f
C385 VDD.n88 VSS 11.7013f
C386 VDD.n89 VSS 2.58977f
C387 VDD.t21 VSS 1.00837f
C388 VDD.n90 VSS 4.95597f
C389 VDD.n91 VSS 8.0135f
C390 VDD.n92 VSS 3.60709f
C391 VDD.t9 VSS 77.235f
C392 VDD.n93 VSS 3.60709f
C393 VDD.n94 VSS 6.68422f
C394 VDD.n95 VSS 7.96035f
C395 VDD.n96 VSS 3.08542f
C396 VDD.n97 VSS 15.0807f
C397 OUT.n0 VSS 50.6208f
C398 OUT.t56 VSS 0.64634f
C399 OUT.t59 VSS 0.64634f
C400 OUT.n1 VSS 2.27605f
C401 OUT.n2 VSS 0.76517f
C402 OUT.n3 VSS 0.01528f
C403 OUT.t0 VSS 0.64634f
C404 OUT.t68 VSS 0.64634f
C405 OUT.n4 VSS 1.32831f
C406 OUT.n5 VSS 0.01019f
C407 OUT.t52 VSS 0.64634f
C408 OUT.t50 VSS 0.64634f
C409 OUT.n6 VSS 1.36083f
C410 OUT.t78 VSS 0.64634f
C411 OUT.t48 VSS 0.64634f
C412 OUT.n7 VSS 2.27603f
C413 OUT.n8 VSS 0.76519f
C414 OUT.t1 VSS 0.64634f
C415 OUT.t61 VSS 0.64634f
C416 OUT.n9 VSS 1.29268f
C417 OUT.n10 VSS 0.76622f
C418 OUT.n11 VSS 1.51892f
C419 OUT.n12 VSS 0.02037f
C420 OUT.t67 VSS 0.64634f
C421 OUT.t75 VSS 0.64634f
C422 OUT.n13 VSS 1.32831f
C423 OUT.t79 VSS 0.64634f
C424 OUT.t54 VSS 0.64634f
C425 OUT.n14 VSS 1.29268f
C426 OUT.n15 VSS 0.76623f
C427 OUT.n16 VSS 1.55154f
C428 OUT.t38 VSS 0.64634f
C429 OUT.t5 VSS 0.64634f
C430 OUT.n17 VSS 1.43962f
C431 OUT.t45 VSS 0.64634f
C432 OUT.t11 VSS 0.64634f
C433 OUT.n18 VSS 2.27608f
C434 OUT.t8 VSS 1.83064f
C435 OUT.n19 VSS 1.94351f
C436 OUT.t25 VSS 1.52934f
C437 OUT.n20 VSS 1.42439f
C438 OUT.t36 VSS 3.1693f
C439 OUT.n21 VSS 0.7668f
C440 OUT.t69 VSS 0.64634f
C441 OUT.t70 VSS 0.64634f
C442 OUT.n22 VSS 2.27595f
C443 OUT.n23 VSS 0.76524f
C444 OUT.t44 VSS 0.64634f
C445 OUT.t16 VSS 0.64634f
C446 OUT.n24 VSS 1.40832f
C447 OUT.n25 VSS 1.47135f
C448 OUT.t40 VSS 0.64634f
C449 OUT.t24 VSS 0.64634f
C450 OUT.n26 VSS 1.29268f
C451 OUT.n27 VSS 0.76625f
C452 OUT.t21 VSS 0.64634f
C453 OUT.t4 VSS 0.64634f
C454 OUT.n28 VSS 2.27603f
C455 OUT.n29 VSS 0.76512f
C456 OUT.n30 VSS 0.01019f
C457 OUT.n31 VSS 0.10172p
C458 OUT.t65 VSS 0.64634f
C459 OUT.t62 VSS 0.64634f
C460 OUT.n32 VSS 2.27603f
C461 OUT.n33 VSS 0.76519f
C462 OUT.t72 VSS 0.64634f
C463 OUT.t58 VSS 0.64634f
C464 OUT.n34 VSS 1.29268f
C465 OUT.n35 VSS 0.76624f
C466 OUT.t80 VSS 0.64634f
C467 OUT.t60 VSS 0.64634f
C468 OUT.n36 VSS 1.29268f
C469 OUT.n37 VSS 1.46835f
C470 OUT.n38 VSS 0.01528f
C471 OUT.t6 VSS 0.64634f
C472 OUT.t37 VSS 0.64634f
C473 OUT.n39 VSS 1.29268f
C474 OUT.t10 VSS 0.64634f
C475 OUT.t30 VSS 0.64634f
C476 OUT.n40 VSS 2.27597f
C477 OUT.t33 VSS 0.64634f
C478 OUT.t27 VSS 0.64634f
C479 OUT.n41 VSS 1.29268f
C480 OUT.n42 VSS 1.40731f
C481 OUT.t34 VSS 0.64634f
C482 OUT.t31 VSS 0.64634f
C483 OUT.n43 VSS 1.29268f
C484 OUT.n44 VSS 0.76629f
C485 OUT.t14 VSS 0.64634f
C486 OUT.t28 VSS 0.64634f
C487 OUT.n45 VSS 2.276f
C488 OUT.n46 VSS 0.76514f
C489 OUT.t42 VSS 1.61869f
C490 OUT.n47 VSS 2.156f
C491 OUT.t18 VSS 1.52934f
C492 OUT.n48 VSS 1.42456f
C493 OUT.t41 VSS 3.16922f
C494 OUT.n49 VSS 0.76686f
C495 OUT.t12 VSS 0.64634f
C496 OUT.t26 VSS 0.64634f
C497 OUT.n50 VSS 1.46812f
C498 OUT.n51 VSS 1.41136f
C499 OUT.t19 VSS 0.64634f
C500 OUT.t23 VSS 0.64634f
C501 OUT.n52 VSS 1.29268f
C502 OUT.n53 VSS 0.76621f
C503 OUT.t35 VSS 0.64634f
C504 OUT.t15 VSS 0.64634f
C505 OUT.n54 VSS 2.276f
C506 OUT.n55 VSS 0.76514f
C507 OUT.n56 VSS 0.01019f
C508 OUT.t81 VSS 1.81528f
C509 OUT.n57 VSS 1.95913f
C510 OUT.t55 VSS 1.63828f
C511 OUT.n58 VSS 1.31553f
C512 OUT.t77 VSS 3.16925f
C513 OUT.n59 VSS 0.76684f
C514 OUT.t84 VSS 1.5174f
C515 OUT.t39 VSS 0.64634f
C516 OUT.t29 VSS 0.64634f
C517 OUT.n60 VSS 1.29268f
C518 OUT.n61 VSS 1.42331f
C519 OUT.t9 VSS 0.64634f
C520 OUT.t20 VSS 0.64634f
C521 OUT.n62 VSS 1.29268f
C522 OUT.n63 VSS 0.76629f
C523 OUT.t17 VSS 0.64634f
C524 OUT.t32 VSS 0.64634f
C525 OUT.n64 VSS 2.27595f
C526 OUT.n65 VSS 0.76518f
C527 OUT.n66 VSS 50.1943f
C528 OUT.n67 VSS 0.01019f
C529 OUT.n68 VSS 0.76516f
C530 OUT.t43 VSS 0.64634f
C531 OUT.t13 VSS 0.64634f
C532 OUT.n69 VSS 1.29268f
C533 OUT.n70 VSS 0.76634f
C534 OUT.n71 VSS 1.58725f
C535 OUT.n72 VSS 0.13455f
C536 OUT.t57 VSS 0.64634f
C537 OUT.t64 VSS 0.64634f
C538 OUT.n73 VSS 1.29268f
C539 OUT.n74 VSS 0.76625f
C540 OUT.t83 VSS 0.64634f
C541 OUT.t53 VSS 0.64634f
C542 OUT.n75 VSS 1.29268f
C543 OUT.n76 VSS 1.43636f
C544 OUT.n77 VSS 0.16158f
C545 OUT.n78 VSS 0.20093f
C546 OUT.t46 VSS 0.64634f
C547 OUT.t2 VSS 0.64634f
C548 OUT.n79 VSS 1.29268f
C549 OUT.n80 VSS 1.40731f
C550 OUT.t66 VSS 0.64634f
C551 OUT.t76 VSS 0.64634f
C552 OUT.n81 VSS 1.29268f
C553 OUT.n82 VSS 0.76625f
C554 OUT.t3 VSS 0.64634f
C555 OUT.t51 VSS 0.64634f
C556 OUT.n83 VSS 2.27595f
C557 OUT.n84 VSS 0.76524f
C558 OUT.n85 VSS 0.01019f
C559 OUT.t63 VSS 1.63828f
C560 OUT.n86 VSS 2.13659f
C561 OUT.t73 VSS 1.63828f
C562 OUT.n87 VSS 1.31771f
C563 OUT.t71 VSS 3.16868f
C564 OUT.n88 VSS 0.777f
C565 OUT.n89 VSS 0.01528f
C566 OUT.n90 VSS 0.76509f
C567 OUT.t22 VSS 0.64634f
C568 OUT.t7 VSS 0.64634f
C569 OUT.n91 VSS 1.29268f
C570 OUT.n92 VSS 0.76621f
C571 OUT.n93 VSS 1.43995f
C572 OUT.n94 VSS 0.01019f
C573 OUT.n95 VSS 1.55154f
C574 OUT.t82 VSS 0.64634f
C575 OUT.t47 VSS 0.64634f
C576 OUT.n96 VSS 1.29268f
C577 OUT.n97 VSS 0.76623f
C578 OUT.t49 VSS 0.64634f
C579 OUT.t74 VSS 0.64634f
C580 OUT.n98 VSS 2.27605f
C581 OUT.n99 VSS 0.76517f
C582 OUT.n100 VSS 50.5134f
C583 x1.ADJ.n0 VSS 0.11837f
C584 x1.ADJ.n1 VSS 0.22101f
C585 x1.ADJ.n2 VSS 3.6619f
C586 x1.ADJ.n3 VSS 0.88445f
C587 x1.ADJ.n4 VSS 1.78693f
C588 x1.ADJ.t27 VSS 1.7629f
C589 x1.ADJ.n5 VSS 0.07419f
C590 x1.ADJ.n6 VSS 0.16828f
C591 x1.ADJ.t40 VSS 1.77067f
C592 x1.ADJ.n7 VSS 0.07419f
C593 x1.ADJ.n8 VSS 0.16828f
C594 x1.ADJ.n9 VSS 0.88539f
C595 x1.ADJ.n10 VSS 0.07419f
C596 x1.ADJ.t45 VSS 1.77106f
C597 x1.ADJ.n11 VSS 0.08581f
C598 x1.ADJ.n12 VSS 0.89584f
C599 x1.ADJ.t6 VSS 1.7629f
C600 x1.ADJ.n13 VSS 1.77991f
C601 x1.ADJ.t37 VSS 1.77067f
C602 x1.ADJ.n14 VSS 1.78981f
C603 x1.ADJ.n15 VSS 0.89773f
C604 x1.ADJ.t43 VSS 1.77067f
C605 x1.ADJ.t22 VSS 1.77067f
C606 x1.ADJ.t8 VSS 1.77067f
C607 x1.ADJ.n16 VSS 1.77991f
C608 x1.ADJ.t35 VSS 1.7629f
C609 x1.ADJ.n17 VSS 1.77991f
C610 x1.ADJ.n18 VSS 0.07419f
C611 x1.ADJ.n19 VSS 0.07419f
C612 x1.ADJ.n20 VSS 1.77991f
C613 x1.ADJ.t11 VSS 1.7629f
C614 x1.ADJ.t28 VSS 1.77067f
C615 x1.ADJ.n21 VSS 1.77991f
C616 x1.ADJ.n22 VSS 0.07419f
C617 x1.ADJ.n23 VSS 0.07419f
C618 x1.ADJ.n24 VSS 1.77991f
C619 x1.ADJ.t20 VSS 1.77067f
C620 x1.ADJ.n25 VSS 1.78693f
C621 x1.ADJ.t30 VSS 1.7711f
C622 x1.ADJ.n26 VSS 1.77991f
C623 x1.ADJ.t13 VSS 1.7629f
C624 x1.ADJ.n27 VSS 1.77991f
C625 x1.ADJ.n28 VSS 0.08581f
C626 x1.ADJ.n29 VSS 3.7736f
C627 x1.ADJ.n30 VSS 0.89773f
C628 x1.ADJ.n31 VSS 0.89773f
C629 x1.ADJ.t38 VSS 1.7629f
C630 x1.ADJ.n32 VSS 0.07419f
C631 x1.ADJ.n33 VSS 0.13103f
C632 x1.ADJ.t21 VSS 1.77067f
C633 x1.ADJ.n34 VSS 0.07419f
C634 x1.ADJ.n35 VSS 0.89584f
C635 x1.ADJ.n36 VSS 0.16828f
C636 x1.ADJ.t12 VSS 1.7629f
C637 x1.ADJ.n37 VSS 0.07419f
C638 x1.ADJ.n38 VSS 1.77991f
C639 x1.ADJ.t44 VSS 1.77067f
C640 x1.ADJ.n39 VSS 1.78981f
C641 x1.ADJ.t18 VSS 1.77106f
C642 x1.ADJ.n40 VSS 1.77991f
C643 x1.ADJ.t31 VSS 1.7629f
C644 x1.ADJ.n41 VSS 1.77991f
C645 x1.ADJ.t4 VSS 1.7711f
C646 x1.ADJ.n42 VSS 1.78693f
C647 x1.ADJ.t29 VSS 1.77067f
C648 x1.ADJ.n43 VSS 1.77991f
C649 x1.ADJ.n44 VSS 0.07419f
C650 x1.ADJ.t36 VSS 1.77067f
C651 x1.ADJ.n45 VSS 1.77991f
C652 x1.ADJ.t3 VSS 1.7629f
C653 x1.ADJ.t19 VSS 1.77067f
C654 x1.ADJ.n46 VSS 1.77991f
C655 x1.ADJ.n47 VSS 0.07419f
C656 x1.ADJ.n48 VSS 0.07419f
C657 x1.ADJ.n49 VSS 1.77991f
C658 x1.ADJ.t15 VSS 1.77067f
C659 x1.ADJ.n50 VSS 0.92668f
C660 x1.ADJ.t24 VSS 1.7711f
C661 x1.ADJ.t26 VSS 1.7629f
C662 x1.ADJ.n51 VSS 1.77991f
C663 x1.ADJ.t16 VSS 1.77067f
C664 x1.ADJ.n52 VSS 1.78981f
C665 x1.ADJ.t39 VSS 1.77106f
C666 x1.ADJ.n53 VSS 1.78112f
C667 x1.ADJ.t10 VSS 1.7629f
C668 x1.ADJ.n54 VSS 1.78113f
C669 x1.ADJ.n55 VSS 0.1313f
C670 x1.ADJ.n56 VSS 1.77991f
C671 x1.ADJ.t41 VSS 1.77067f
C672 x1.ADJ.n57 VSS 1.78693f
C673 x1.ADJ.n58 VSS 0.89584f
C674 x1.ADJ.t7 VSS 1.77067f
C675 x1.ADJ.n59 VSS 1.77991f
C676 x1.ADJ.t34 VSS 1.7629f
C677 x1.ADJ.n60 VSS 1.77991f
C678 x1.ADJ.n61 VSS 0.07419f
C679 x1.ADJ.n62 VSS 0.07419f
C680 x1.ADJ.n63 VSS 1.77991f
C681 x1.ADJ.t33 VSS 1.77067f
C682 x1.ADJ.n64 VSS 1.09506f
C683 x1.ADJ.n65 VSS 1.95263f
C684 x1.ADJ.n66 VSS 0.01248f
C685 x1.ADJ.n67 VSS 1.77991f
C686 x1.ADJ.t17 VSS 1.77067f
C687 x1.ADJ.n68 VSS 0.89758f
C688 x1.ADJ.n69 VSS 1.78981f
C689 x1.ADJ.t5 VSS 1.77106f
C690 x1.ADJ.t32 VSS 1.7711f
C691 x1.ADJ.n70 VSS 1.77991f
C692 x1.ADJ.t14 VSS 1.7629f
C693 x1.ADJ.n71 VSS 1.77991f
C694 x1.ADJ.n72 VSS 0.16828f
C695 x1.ADJ.n73 VSS 0.07419f
C696 x1.ADJ.n74 VSS 1.77991f
C697 x1.ADJ.t9 VSS 1.7629f
C698 x1.ADJ.t25 VSS 1.77067f
C699 x1.ADJ.n75 VSS 1.77991f
C700 x1.ADJ.n76 VSS 0.07419f
C701 x1.ADJ.n77 VSS 0.07419f
C702 x1.ADJ.n78 VSS 1.77991f
C703 x1.ADJ.t42 VSS 1.77067f
C704 x1.ADJ.n79 VSS 0.89572f
C705 x1.ADJ.n80 VSS 0.01151f
C706 x1.ADJ.n81 VSS 0.1704f
C707 x1.ADJ.n82 VSS 1.88927f
C708 x1.ADJ.n83 VSS 0.16583f
C709 x1.ADJ.t0 VSS 0.28804f
C710 x1.ADJ.n84 VSS 0.1522f
C711 x1.ADJ.t1 VSS 0.38096f
C712 x1.ADJ.n85 VSS 0.41248f
C713 x1.ADJ.n86 VSS 0.26011f
C714 x1.ADJ.t23 VSS 0.28871f
C715 x1.ADJ.n87 VSS 0.19674f
C716 x1.ADJ.t2 VSS 0.03385f
.ends

