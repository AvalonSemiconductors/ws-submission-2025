VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aef2
  CLASS BLOCK ;
  FOREIGN aef2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 236.000 BY 188.000 ;
  OBS
      LAYER Metal5 ;
        RECT 86.000 181.500 97.000 182.000 ;
        RECT 81.000 181.000 102.000 181.500 ;
        RECT 77.500 180.500 105.500 181.000 ;
        RECT 74.500 180.000 108.500 180.500 ;
        RECT 72.000 179.500 111.000 180.000 ;
        RECT 70.000 179.000 113.000 179.500 ;
        RECT 68.000 178.500 83.500 179.000 ;
        RECT 99.500 178.500 115.000 179.000 ;
        RECT 66.500 178.000 79.500 178.500 ;
        RECT 103.500 178.000 116.500 178.500 ;
        RECT 65.000 177.500 76.500 178.000 ;
        RECT 107.000 177.500 118.000 178.000 ;
        RECT 63.500 177.000 74.000 177.500 ;
        RECT 109.500 177.000 119.500 177.500 ;
        RECT 62.000 176.500 71.500 177.000 ;
        RECT 111.500 176.500 121.000 177.000 ;
        RECT 60.500 176.000 69.500 176.500 ;
        RECT 113.500 176.000 122.500 176.500 ;
        RECT 59.500 175.500 68.000 176.000 ;
        RECT 113.500 175.500 123.500 176.000 ;
        RECT 58.000 175.000 66.000 175.500 ;
        RECT 113.500 175.000 125.000 175.500 ;
        RECT 57.000 174.500 64.500 175.000 ;
        RECT 111.500 174.500 126.000 175.000 ;
        RECT 56.000 174.000 63.000 174.500 ;
        RECT 109.500 174.000 127.000 174.500 ;
        RECT 54.500 173.500 62.000 174.000 ;
        RECT 107.500 173.500 128.500 174.000 ;
        RECT 53.500 173.000 60.500 173.500 ;
        RECT 105.500 173.000 129.500 173.500 ;
        RECT 52.500 172.500 59.500 173.000 ;
        RECT 104.000 172.500 130.500 173.000 ;
        RECT 51.500 172.000 58.000 172.500 ;
        RECT 102.000 172.000 131.500 172.500 ;
        RECT 50.500 171.500 57.000 172.000 ;
        RECT 100.500 171.500 132.500 172.000 ;
        RECT 49.500 171.000 56.000 171.500 ;
        RECT 98.500 171.000 133.000 171.500 ;
        RECT 49.000 170.500 55.000 171.000 ;
        RECT 97.000 170.500 134.000 171.000 ;
        RECT 48.000 170.000 54.000 170.500 ;
        RECT 95.500 170.000 135.000 170.500 ;
        RECT 47.000 169.500 53.000 170.000 ;
        RECT 94.500 169.500 136.000 170.000 ;
        RECT 46.500 169.000 52.000 169.500 ;
        RECT 93.000 169.000 136.500 169.500 ;
        RECT 211.500 169.000 212.500 169.500 ;
        RECT 45.500 168.500 51.000 169.000 ;
        RECT 91.500 168.500 137.500 169.000 ;
        RECT 210.500 168.500 213.500 169.000 ;
        RECT 44.500 168.000 50.000 168.500 ;
        RECT 90.000 168.000 138.500 168.500 ;
        RECT 209.500 168.000 214.000 168.500 ;
        RECT 44.000 167.500 49.500 168.000 ;
        RECT 89.000 167.500 130.500 168.000 ;
        RECT 134.000 167.500 139.000 168.000 ;
        RECT 209.000 167.500 214.500 168.000 ;
        RECT 43.000 167.000 48.500 167.500 ;
        RECT 87.500 167.000 128.500 167.500 ;
        RECT 134.500 167.000 140.000 167.500 ;
        RECT 208.500 167.000 214.500 167.500 ;
        RECT 42.500 166.500 47.500 167.000 ;
        RECT 86.500 166.500 126.500 167.000 ;
        RECT 135.500 166.500 140.500 167.000 ;
        RECT 208.000 166.500 215.000 167.000 ;
        RECT 41.500 166.000 47.000 166.500 ;
        RECT 85.000 166.000 124.500 166.500 ;
        RECT 136.500 166.000 141.500 166.500 ;
        RECT 207.500 166.000 215.000 166.500 ;
        RECT 41.000 165.500 46.000 166.000 ;
        RECT 84.000 165.500 123.000 166.000 ;
        RECT 137.000 165.500 142.000 166.000 ;
        RECT 207.000 165.500 211.000 166.000 ;
        RECT 40.500 165.000 45.500 165.500 ;
        RECT 83.000 165.000 121.000 165.500 ;
        RECT 138.000 165.000 142.500 165.500 ;
        RECT 206.000 165.000 210.500 165.500 ;
        RECT 212.000 165.000 215.000 166.000 ;
        RECT 39.500 164.500 44.500 165.000 ;
        RECT 82.000 164.500 119.000 165.000 ;
        RECT 138.500 164.500 143.500 165.000 ;
        RECT 205.500 164.500 210.000 165.000 ;
        RECT 39.000 164.000 44.000 164.500 ;
        RECT 81.000 164.000 117.500 164.500 ;
        RECT 139.500 164.000 144.000 164.500 ;
        RECT 205.000 164.000 209.500 164.500 ;
        RECT 38.500 163.500 43.000 164.000 ;
        RECT 80.000 163.500 116.000 164.000 ;
        RECT 140.000 163.500 144.500 164.000 ;
        RECT 204.500 163.500 209.000 164.000 ;
        RECT 37.500 163.000 42.500 163.500 ;
        RECT 79.000 163.000 114.500 163.500 ;
        RECT 140.500 163.000 145.500 163.500 ;
        RECT 203.500 163.000 208.000 163.500 ;
        RECT 37.000 162.500 41.500 163.000 ;
        RECT 78.000 162.500 113.000 163.000 ;
        RECT 141.500 162.500 146.000 163.000 ;
        RECT 203.000 162.500 207.500 163.000 ;
        RECT 212.500 162.500 215.000 165.000 ;
        RECT 36.500 162.000 41.000 162.500 ;
        RECT 77.000 162.000 111.500 162.500 ;
        RECT 142.000 162.000 146.500 162.500 ;
        RECT 202.500 162.000 207.000 162.500 ;
        RECT 36.000 161.500 40.500 162.000 ;
        RECT 76.000 161.500 110.500 162.000 ;
        RECT 142.500 161.500 147.000 162.000 ;
        RECT 201.500 161.500 206.500 162.000 ;
        RECT 35.000 161.000 39.500 161.500 ;
        RECT 75.000 161.000 109.000 161.500 ;
        RECT 143.500 161.000 148.000 161.500 ;
        RECT 201.000 161.000 205.500 161.500 ;
        RECT 34.500 160.500 39.000 161.000 ;
        RECT 74.000 160.500 107.500 161.000 ;
        RECT 144.000 160.500 148.500 161.000 ;
        RECT 200.500 160.500 205.000 161.000 ;
        RECT 34.000 160.000 38.500 160.500 ;
        RECT 73.500 160.000 106.500 160.500 ;
        RECT 144.500 160.000 149.000 160.500 ;
        RECT 199.500 160.000 204.500 160.500 ;
        RECT 33.500 159.500 38.000 160.000 ;
        RECT 72.500 159.500 105.000 160.000 ;
        RECT 145.000 159.500 149.500 160.000 ;
        RECT 199.000 159.500 204.000 160.000 ;
        RECT 33.000 159.000 37.000 159.500 ;
        RECT 71.500 159.000 104.000 159.500 ;
        RECT 146.000 159.000 150.000 159.500 ;
        RECT 198.500 159.000 203.000 159.500 ;
        RECT 32.500 158.500 36.500 159.000 ;
        RECT 71.000 158.500 102.500 159.000 ;
        RECT 146.500 158.500 150.500 159.000 ;
        RECT 197.500 158.500 202.500 159.000 ;
        RECT 32.000 158.000 36.000 158.500 ;
        RECT 70.000 158.000 101.500 158.500 ;
        RECT 147.000 158.000 151.000 158.500 ;
        RECT 197.000 158.000 202.000 158.500 ;
        RECT 212.500 158.000 215.500 162.500 ;
        RECT 31.500 157.500 35.500 158.000 ;
        RECT 69.000 157.500 100.500 158.000 ;
        RECT 147.500 157.500 151.500 158.000 ;
        RECT 196.000 157.500 201.000 158.000 ;
        RECT 31.000 157.000 35.000 157.500 ;
        RECT 68.500 157.000 99.500 157.500 ;
        RECT 148.000 157.000 152.000 157.500 ;
        RECT 195.500 157.000 200.500 157.500 ;
        RECT 30.500 156.500 34.500 157.000 ;
        RECT 67.500 156.500 98.500 157.000 ;
        RECT 148.500 156.500 152.500 157.000 ;
        RECT 194.500 156.500 199.500 157.000 ;
        RECT 30.000 156.000 34.000 156.500 ;
        RECT 67.000 156.000 97.000 156.500 ;
        RECT 149.000 156.000 153.000 156.500 ;
        RECT 193.500 156.000 199.000 156.500 ;
        RECT 29.500 155.500 33.500 156.000 ;
        RECT 66.000 155.500 96.000 156.000 ;
        RECT 149.500 155.500 153.500 156.000 ;
        RECT 193.000 155.500 198.000 156.000 ;
        RECT 29.000 155.000 33.000 155.500 ;
        RECT 65.500 155.000 95.000 155.500 ;
        RECT 150.000 155.000 154.000 155.500 ;
        RECT 192.000 155.000 197.500 155.500 ;
        RECT 212.500 155.000 215.000 158.000 ;
        RECT 28.500 154.500 32.500 155.000 ;
        RECT 64.500 154.500 94.000 155.000 ;
        RECT 151.000 154.500 154.500 155.000 ;
        RECT 191.000 154.500 196.500 155.000 ;
        RECT 28.000 154.000 32.000 154.500 ;
        RECT 64.000 154.000 93.500 154.500 ;
        RECT 151.500 154.000 155.000 154.500 ;
        RECT 190.000 154.000 196.000 154.500 ;
        RECT 27.500 153.500 31.500 154.000 ;
        RECT 63.500 153.500 92.500 154.000 ;
        RECT 151.500 153.500 155.500 154.000 ;
        RECT 189.000 153.500 195.000 154.000 ;
        RECT 27.000 153.000 31.000 153.500 ;
        RECT 62.500 153.000 91.500 153.500 ;
        RECT 152.000 153.000 156.000 153.500 ;
        RECT 188.000 153.000 194.000 153.500 ;
        RECT 26.500 152.500 30.500 153.000 ;
        RECT 62.000 152.500 90.500 153.000 ;
        RECT 152.500 152.500 156.500 153.000 ;
        RECT 187.000 152.500 193.500 153.000 ;
        RECT 26.000 152.000 30.000 152.500 ;
        RECT 61.000 152.000 89.500 152.500 ;
        RECT 153.000 152.000 157.000 152.500 ;
        RECT 186.000 152.000 192.500 152.500 ;
        RECT 25.500 151.500 29.500 152.000 ;
        RECT 60.500 151.500 88.500 152.000 ;
        RECT 153.500 151.500 157.500 152.000 ;
        RECT 185.000 151.500 191.500 152.000 ;
        RECT 212.000 151.500 215.000 155.000 ;
        RECT 25.000 151.000 29.000 151.500 ;
        RECT 60.000 151.000 88.000 151.500 ;
        RECT 154.000 151.000 158.000 151.500 ;
        RECT 183.500 151.000 190.500 151.500 ;
        RECT 25.000 150.500 28.500 151.000 ;
        RECT 59.500 150.500 87.000 151.000 ;
        RECT 154.500 150.500 158.000 151.000 ;
        RECT 182.500 150.500 189.500 151.000 ;
        RECT 212.000 150.500 214.500 151.500 ;
        RECT 24.500 150.000 28.000 150.500 ;
        RECT 58.500 150.000 86.000 150.500 ;
        RECT 155.000 150.000 158.500 150.500 ;
        RECT 181.000 150.000 188.500 150.500 ;
        RECT 24.000 149.500 27.500 150.000 ;
        RECT 58.000 149.500 85.500 150.000 ;
        RECT 155.500 149.500 159.000 150.000 ;
        RECT 180.000 149.500 187.500 150.000 ;
        RECT 23.500 149.000 27.000 149.500 ;
        RECT 57.500 149.000 84.500 149.500 ;
        RECT 156.000 149.000 159.500 149.500 ;
        RECT 179.000 149.000 186.000 149.500 ;
        RECT 23.000 148.500 27.000 149.000 ;
        RECT 57.000 148.500 83.500 149.000 ;
        RECT 156.000 148.500 160.000 149.000 ;
        RECT 177.500 148.500 185.000 149.000 ;
        RECT 23.000 148.000 26.500 148.500 ;
        RECT 56.500 148.000 83.000 148.500 ;
        RECT 156.500 148.000 160.000 148.500 ;
        RECT 176.500 148.000 183.500 148.500 ;
        RECT 211.500 148.000 214.500 150.500 ;
        RECT 22.500 147.500 26.000 148.000 ;
        RECT 56.000 147.500 82.000 148.000 ;
        RECT 157.000 147.500 160.500 148.000 ;
        RECT 175.500 147.500 182.500 148.000 ;
        RECT 22.000 147.000 25.500 147.500 ;
        RECT 55.000 147.000 81.500 147.500 ;
        RECT 157.500 147.000 161.000 147.500 ;
        RECT 174.500 147.000 181.500 147.500 ;
        RECT 211.500 147.000 214.000 148.000 ;
        RECT 21.500 146.000 25.000 147.000 ;
        RECT 54.500 146.500 80.500 147.000 ;
        RECT 158.000 146.500 161.500 147.000 ;
        RECT 173.000 146.500 180.000 147.000 ;
        RECT 54.000 146.000 80.000 146.500 ;
        RECT 158.000 146.000 162.000 146.500 ;
        RECT 172.000 146.000 179.000 146.500 ;
        RECT 21.000 145.500 24.500 146.000 ;
        RECT 53.500 145.500 79.000 146.000 ;
        RECT 158.500 145.500 162.000 146.000 ;
        RECT 171.500 145.500 178.000 146.000 ;
        RECT 20.500 145.000 24.000 145.500 ;
        RECT 53.000 145.000 78.500 145.500 ;
        RECT 159.000 145.000 162.500 145.500 ;
        RECT 170.500 145.000 176.500 145.500 ;
        RECT 211.000 145.000 214.000 147.000 ;
        RECT 20.000 144.000 23.500 145.000 ;
        RECT 52.500 144.500 77.500 145.000 ;
        RECT 52.000 144.000 77.000 144.500 ;
        RECT 159.500 144.000 163.000 145.000 ;
        RECT 169.500 144.500 175.500 145.000 ;
        RECT 211.000 144.500 213.500 145.000 ;
        RECT 168.500 144.000 174.500 144.500 ;
        RECT 19.500 143.500 23.000 144.000 ;
        RECT 51.500 143.500 76.000 144.000 ;
        RECT 160.000 143.500 163.500 144.000 ;
        RECT 167.500 143.500 173.500 144.000 ;
        RECT 19.000 142.500 22.500 143.500 ;
        RECT 51.000 143.000 75.500 143.500 ;
        RECT 160.500 143.000 164.000 143.500 ;
        RECT 166.500 143.000 172.500 143.500 ;
        RECT 50.500 142.500 75.000 143.000 ;
        RECT 161.000 142.500 164.000 143.000 ;
        RECT 166.000 142.500 171.500 143.000 ;
        RECT 210.500 142.500 213.500 144.500 ;
        RECT 18.500 142.000 22.000 142.500 ;
        RECT 50.000 142.000 74.000 142.500 ;
        RECT 161.000 142.000 170.500 142.500 ;
        RECT 210.500 142.000 213.000 142.500 ;
        RECT 18.000 141.500 21.500 142.000 ;
        RECT 49.500 141.500 73.500 142.000 ;
        RECT 161.500 141.500 170.000 142.000 ;
        RECT 18.000 141.000 21.000 141.500 ;
        RECT 49.000 141.000 73.000 141.500 ;
        RECT 162.000 141.000 169.000 141.500 ;
        RECT 17.500 140.500 21.000 141.000 ;
        RECT 48.500 140.500 72.000 141.000 ;
        RECT 162.000 140.500 168.000 141.000 ;
        RECT 210.000 140.500 213.000 142.000 ;
        RECT 17.500 140.000 20.500 140.500 ;
        RECT 48.000 140.000 71.500 140.500 ;
        RECT 162.500 140.000 167.000 140.500 ;
        RECT 210.000 140.000 212.500 140.500 ;
        RECT 17.000 139.500 20.500 140.000 ;
        RECT 47.500 139.500 71.000 140.000 ;
        RECT 163.000 139.500 166.500 140.000 ;
        RECT 16.500 139.000 20.000 139.500 ;
        RECT 47.000 139.000 70.500 139.500 ;
        RECT 163.000 139.000 165.500 139.500 ;
        RECT 16.500 138.500 19.500 139.000 ;
        RECT 46.500 138.500 70.000 139.000 ;
        RECT 163.500 138.500 165.500 139.000 ;
        RECT 16.000 138.000 19.500 138.500 ;
        RECT 46.000 138.000 69.000 138.500 ;
        RECT 163.500 138.000 166.000 138.500 ;
        RECT 209.500 138.000 212.500 140.000 ;
        RECT 16.000 137.500 19.000 138.000 ;
        RECT 45.500 137.500 68.500 138.000 ;
        RECT 164.000 137.500 166.000 138.000 ;
        RECT 15.500 137.000 18.500 137.500 ;
        RECT 45.000 137.000 68.000 137.500 ;
        RECT 15.000 136.500 18.500 137.000 ;
        RECT 44.500 136.500 67.500 137.000 ;
        RECT 164.500 136.500 166.500 137.500 ;
        RECT 209.000 136.500 212.000 138.000 ;
        RECT 15.000 136.000 18.000 136.500 ;
        RECT 44.000 136.000 67.000 136.500 ;
        RECT 14.500 135.500 18.000 136.000 ;
        RECT 43.500 135.500 66.000 136.000 ;
        RECT 165.000 135.500 167.000 136.500 ;
        RECT 209.000 136.000 211.500 136.500 ;
        RECT 14.500 135.000 17.500 135.500 ;
        RECT 43.500 135.000 65.500 135.500 ;
        RECT 165.500 135.000 167.500 135.500 ;
        RECT 14.000 134.500 17.500 135.000 ;
        RECT 43.000 134.500 65.000 135.000 ;
        RECT 165.500 134.500 168.000 135.000 ;
        RECT 14.000 134.000 17.000 134.500 ;
        RECT 42.500 134.000 64.500 134.500 ;
        RECT 142.000 134.000 154.000 134.500 ;
        RECT 13.500 133.500 17.000 134.000 ;
        RECT 42.000 133.500 64.000 134.000 ;
        RECT 84.000 133.500 85.000 134.000 ;
        RECT 139.000 133.500 157.500 134.000 ;
        RECT 166.000 133.500 168.000 134.500 ;
        RECT 208.500 134.500 211.500 136.000 ;
        RECT 208.500 134.000 211.000 134.500 ;
        RECT 13.500 133.000 16.500 133.500 ;
        RECT 41.500 133.000 63.500 133.500 ;
        RECT 84.000 133.000 85.500 133.500 ;
        RECT 136.500 133.000 159.500 133.500 ;
        RECT 13.000 132.500 16.500 133.000 ;
        RECT 41.000 132.500 63.000 133.000 ;
        RECT 13.000 132.000 16.000 132.500 ;
        RECT 12.500 131.500 16.000 132.000 ;
        RECT 40.500 132.000 62.500 132.500 ;
        RECT 83.500 132.000 86.000 133.000 ;
        RECT 134.500 132.500 143.000 133.000 ;
        RECT 153.500 132.500 162.000 133.000 ;
        RECT 166.500 132.500 168.500 133.500 ;
        RECT 208.000 132.500 211.000 134.000 ;
        RECT 229.000 133.500 230.500 134.000 ;
        RECT 228.000 133.000 231.500 133.500 ;
        RECT 227.000 132.500 232.000 133.000 ;
        RECT 133.000 132.000 139.500 132.500 ;
        RECT 157.000 132.000 163.500 132.500 ;
        RECT 40.500 131.500 62.000 132.000 ;
        RECT 12.500 130.500 15.500 131.500 ;
        RECT 40.000 131.000 61.500 131.500 ;
        RECT 83.000 131.000 86.500 132.000 ;
        RECT 131.500 131.500 137.000 132.000 ;
        RECT 159.500 131.500 165.000 132.000 ;
        RECT 167.000 131.500 169.000 132.500 ;
        RECT 130.000 131.000 135.000 131.500 ;
        RECT 161.000 131.000 169.500 131.500 ;
        RECT 39.500 130.500 61.000 131.000 ;
        RECT 82.500 130.500 87.000 131.000 ;
        RECT 128.500 130.500 133.500 131.000 ;
        RECT 163.000 130.500 169.500 131.000 ;
        RECT 207.500 131.000 210.500 132.500 ;
        RECT 226.000 132.000 232.000 132.500 ;
        RECT 225.000 131.500 232.500 132.000 ;
        RECT 224.500 131.000 232.500 131.500 ;
        RECT 207.500 130.500 210.000 131.000 ;
        RECT 223.500 130.500 232.500 131.000 ;
        RECT 12.000 129.500 15.000 130.500 ;
        RECT 39.000 130.000 60.500 130.500 ;
        RECT 82.500 130.000 87.500 130.500 ;
        RECT 127.500 130.000 132.000 130.500 ;
        RECT 164.500 130.000 170.000 130.500 ;
        RECT 38.500 129.500 60.000 130.000 ;
        RECT 82.000 129.500 87.500 130.000 ;
        RECT 126.500 129.500 130.500 130.000 ;
        RECT 166.000 129.500 171.000 130.000 ;
        RECT 11.500 128.500 14.500 129.500 ;
        RECT 38.500 129.000 59.500 129.500 ;
        RECT 38.000 128.500 59.000 129.000 ;
        RECT 82.000 128.500 88.000 129.500 ;
        RECT 125.500 129.000 129.500 129.500 ;
        RECT 167.000 129.000 172.000 129.500 ;
        RECT 207.000 129.000 210.000 130.500 ;
        RECT 222.500 130.000 228.500 130.500 ;
        RECT 221.500 129.500 227.500 130.000 ;
        RECT 221.000 129.000 226.500 129.500 ;
        RECT 124.500 128.500 128.000 129.000 ;
        RECT 168.000 128.500 173.000 129.000 ;
        RECT 11.000 127.000 14.000 128.500 ;
        RECT 37.500 128.000 58.500 128.500 ;
        RECT 37.000 127.500 58.000 128.000 ;
        RECT 81.500 127.500 88.500 128.500 ;
        RECT 123.500 128.000 127.000 128.500 ;
        RECT 169.000 128.000 174.000 128.500 ;
        RECT 122.500 127.500 126.000 128.000 ;
        RECT 170.000 127.500 175.000 128.000 ;
        RECT 206.500 127.500 209.500 129.000 ;
        RECT 220.000 128.500 225.500 129.000 ;
        RECT 219.000 128.000 225.000 128.500 ;
        RECT 229.500 128.000 232.500 130.500 ;
        RECT 218.000 127.500 224.000 128.000 ;
        RECT 37.000 127.000 57.500 127.500 ;
        RECT 81.500 127.000 89.000 127.500 ;
        RECT 122.000 127.000 125.000 127.500 ;
        RECT 171.000 127.000 175.500 127.500 ;
        RECT 10.500 126.000 13.500 127.000 ;
        RECT 36.500 126.500 57.000 127.000 ;
        RECT 36.000 126.000 56.500 126.500 ;
        RECT 81.000 126.000 89.500 127.000 ;
        RECT 121.000 126.500 124.000 127.000 ;
        RECT 172.000 126.500 176.500 127.000 ;
        RECT 120.500 126.000 123.500 126.500 ;
        RECT 173.000 126.000 177.000 126.500 ;
        RECT 206.000 126.000 209.000 127.500 ;
        RECT 217.000 127.000 223.000 127.500 ;
        RECT 215.500 126.500 222.000 127.000 ;
        RECT 229.500 126.500 232.000 128.000 ;
        RECT 214.500 126.000 221.000 126.500 ;
        RECT 10.000 124.500 13.000 126.000 ;
        RECT 35.500 125.500 56.000 126.000 ;
        RECT 35.500 125.000 55.500 125.500 ;
        RECT 80.500 125.000 90.000 126.000 ;
        RECT 119.500 125.500 122.500 126.000 ;
        RECT 174.000 125.500 178.000 126.000 ;
        RECT 119.000 125.000 121.500 125.500 ;
        RECT 174.500 125.000 178.500 125.500 ;
        RECT 35.000 124.500 55.000 125.000 ;
        RECT 80.500 124.500 90.500 125.000 ;
        RECT 118.000 124.500 121.000 125.000 ;
        RECT 175.500 124.500 179.000 125.000 ;
        RECT 205.500 124.500 208.500 126.000 ;
        RECT 213.500 125.500 220.000 126.000 ;
        RECT 212.000 125.000 219.000 125.500 ;
        RECT 211.000 124.500 218.000 125.000 ;
        RECT 9.500 123.500 12.500 124.500 ;
        RECT 34.500 124.000 54.500 124.500 ;
        RECT 80.000 124.000 91.000 124.500 ;
        RECT 117.500 124.000 120.000 124.500 ;
        RECT 176.000 124.000 180.000 124.500 ;
        RECT 205.000 124.000 208.500 124.500 ;
        RECT 209.500 124.000 217.000 124.500 ;
        RECT 34.500 123.500 54.000 124.000 ;
        RECT 79.500 123.500 92.500 124.000 ;
        RECT 117.000 123.500 119.500 124.000 ;
        RECT 177.000 123.500 180.500 124.000 ;
        RECT 205.000 123.500 216.000 124.000 ;
        RECT 229.000 123.500 232.000 126.500 ;
        RECT 9.500 123.000 12.000 123.500 ;
        RECT 34.000 123.000 53.500 123.500 ;
        RECT 79.000 123.000 93.500 123.500 ;
        RECT 116.000 123.000 119.000 123.500 ;
        RECT 177.500 123.000 181.000 123.500 ;
        RECT 204.500 123.000 215.000 123.500 ;
        RECT 229.000 123.000 231.500 123.500 ;
        RECT 9.000 122.000 12.000 123.000 ;
        RECT 33.500 122.500 53.000 123.000 ;
        RECT 78.000 122.500 95.000 123.000 ;
        RECT 115.500 122.500 118.000 123.000 ;
        RECT 178.000 122.500 181.500 123.000 ;
        RECT 202.000 122.500 213.500 123.000 ;
        RECT 33.000 122.000 53.000 122.500 ;
        RECT 77.500 122.000 96.500 122.500 ;
        RECT 115.000 122.000 117.500 122.500 ;
        RECT 178.500 122.000 182.000 122.500 ;
        RECT 200.000 122.000 212.000 122.500 ;
        RECT 9.000 121.500 11.500 122.000 ;
        RECT 33.000 121.500 52.500 122.000 ;
        RECT 76.500 121.500 97.500 122.000 ;
        RECT 114.500 121.500 117.000 122.000 ;
        RECT 179.500 121.500 182.500 122.000 ;
        RECT 198.000 121.500 210.500 122.000 ;
        RECT 8.500 120.500 11.500 121.500 ;
        RECT 32.500 121.000 52.000 121.500 ;
        RECT 75.500 121.000 99.000 121.500 ;
        RECT 114.000 121.000 116.500 121.500 ;
        RECT 180.000 121.000 183.500 121.500 ;
        RECT 196.000 121.000 209.000 121.500 ;
        RECT 32.000 120.500 51.500 121.000 ;
        RECT 74.500 120.500 100.000 121.000 ;
        RECT 113.500 120.500 116.000 121.000 ;
        RECT 180.500 120.500 184.000 121.000 ;
        RECT 194.500 120.500 207.500 121.000 ;
        RECT 228.500 120.500 231.500 123.000 ;
        RECT 8.500 120.000 11.000 120.500 ;
        RECT 32.000 120.000 51.000 120.500 ;
        RECT 73.500 120.000 100.500 120.500 ;
        RECT 113.000 120.000 115.000 120.500 ;
        RECT 181.000 120.000 184.500 120.500 ;
        RECT 192.500 120.000 205.500 120.500 ;
        RECT 228.500 120.000 231.000 120.500 ;
        RECT 8.000 118.500 11.000 120.000 ;
        RECT 31.500 119.500 50.500 120.000 ;
        RECT 73.000 119.500 101.000 120.000 ;
        RECT 112.500 119.500 114.500 120.000 ;
        RECT 181.500 119.500 185.000 120.000 ;
        RECT 191.000 119.500 203.000 120.000 ;
        RECT 31.000 118.500 50.000 119.500 ;
        RECT 72.000 119.000 100.500 119.500 ;
        RECT 112.000 119.000 114.000 119.500 ;
        RECT 182.000 119.000 185.500 119.500 ;
        RECT 189.500 119.000 201.000 119.500 ;
        RECT 71.500 118.500 99.500 119.000 ;
        RECT 111.500 118.500 113.500 119.000 ;
        RECT 182.500 118.500 185.500 119.000 ;
        RECT 188.000 118.500 198.500 119.000 ;
        RECT 7.500 117.000 10.500 118.500 ;
        RECT 30.500 118.000 49.500 118.500 ;
        RECT 70.500 118.000 99.000 118.500 ;
        RECT 111.000 118.000 113.000 118.500 ;
        RECT 183.000 118.000 196.500 118.500 ;
        RECT 228.000 118.000 231.000 120.000 ;
        RECT 30.000 117.500 49.000 118.000 ;
        RECT 70.500 117.500 98.000 118.000 ;
        RECT 110.500 117.500 112.500 118.000 ;
        RECT 183.500 117.500 194.500 118.000 ;
        RECT 228.000 117.500 230.500 118.000 ;
        RECT 30.000 117.000 48.500 117.500 ;
        RECT 71.000 117.000 97.500 117.500 ;
        RECT 110.000 117.000 112.000 117.500 ;
        RECT 184.000 117.000 192.500 117.500 ;
        RECT 7.500 116.500 10.000 117.000 ;
        RECT 7.000 115.000 10.000 116.500 ;
        RECT 29.500 116.000 48.000 117.000 ;
        RECT 71.500 116.500 96.500 117.000 ;
        RECT 109.500 116.500 111.500 117.000 ;
        RECT 184.500 116.500 190.500 117.000 ;
        RECT 73.000 116.000 95.500 116.500 ;
        RECT 109.000 116.000 111.500 116.500 ;
        RECT 185.000 116.000 189.000 116.500 ;
        RECT 227.500 116.000 230.500 117.500 ;
        RECT 29.000 115.500 47.500 116.000 ;
        RECT 74.000 115.500 94.500 116.000 ;
        RECT 109.000 115.500 111.000 116.000 ;
        RECT 185.500 115.500 188.000 116.000 ;
        RECT 227.500 115.500 230.000 116.000 ;
        RECT 28.500 115.000 47.000 115.500 ;
        RECT 75.000 115.000 93.500 115.500 ;
        RECT 108.500 115.000 110.500 115.500 ;
        RECT 186.000 115.000 188.000 115.500 ;
        RECT 7.000 114.500 9.500 115.000 ;
        RECT 28.500 114.500 46.500 115.000 ;
        RECT 76.500 114.500 93.000 115.000 ;
        RECT 108.000 114.500 110.000 115.000 ;
        RECT 186.000 114.500 188.500 115.000 ;
        RECT 6.500 113.000 9.500 114.500 ;
        RECT 28.000 114.000 46.500 114.500 ;
        RECT 78.000 114.000 92.000 114.500 ;
        RECT 27.500 113.500 46.000 114.000 ;
        RECT 79.000 113.500 91.500 114.000 ;
        RECT 107.500 113.500 109.500 114.500 ;
        RECT 186.500 114.000 188.500 114.500 ;
        RECT 227.000 114.000 230.000 115.500 ;
        RECT 187.000 113.500 189.000 114.000 ;
        RECT 227.000 113.500 229.500 114.000 ;
        RECT 27.500 113.000 45.500 113.500 ;
        RECT 80.000 113.000 91.000 113.500 ;
        RECT 107.000 113.000 109.000 113.500 ;
        RECT 6.500 112.000 9.000 113.000 ;
        RECT 27.000 112.000 45.000 113.000 ;
        RECT 81.000 112.500 91.000 113.000 ;
        RECT 106.500 112.500 108.500 113.000 ;
        RECT 187.500 112.500 189.500 113.500 ;
        RECT 81.000 112.000 90.500 112.500 ;
        RECT 6.000 110.500 9.000 112.000 ;
        RECT 26.500 111.500 44.500 112.000 ;
        RECT 26.000 111.000 44.000 111.500 ;
        RECT 81.500 111.000 90.500 112.000 ;
        RECT 106.000 111.500 108.000 112.500 ;
        RECT 188.000 112.000 190.000 112.500 ;
        RECT 226.500 112.000 229.500 113.500 ;
        RECT 188.500 111.500 190.500 112.000 ;
        RECT 105.500 111.000 107.500 111.500 ;
        RECT 189.000 111.000 190.500 111.500 ;
        RECT 26.000 110.500 43.500 111.000 ;
        RECT 82.000 110.500 90.000 111.000 ;
        RECT 6.000 109.500 8.500 110.500 ;
        RECT 25.500 110.000 43.500 110.500 ;
        RECT 82.500 110.000 90.000 110.500 ;
        RECT 105.000 110.000 107.000 111.000 ;
        RECT 189.000 110.500 191.000 111.000 ;
        RECT 226.000 110.500 229.000 112.000 ;
        RECT 25.500 109.500 43.000 110.000 ;
        RECT 82.500 109.500 89.500 110.000 ;
        RECT 5.500 107.500 8.500 109.500 ;
        RECT 25.000 108.500 42.500 109.500 ;
        RECT 83.000 108.500 89.500 109.500 ;
        RECT 104.500 109.500 106.500 110.000 ;
        RECT 189.500 109.500 191.500 110.500 ;
        RECT 226.000 110.000 228.500 110.500 ;
        RECT 104.500 109.000 106.000 109.500 ;
        RECT 190.000 109.000 192.000 109.500 ;
        RECT 104.000 108.500 106.000 109.000 ;
        RECT 190.500 108.500 192.000 109.000 ;
        RECT 225.500 108.500 228.500 110.000 ;
        RECT 24.500 108.000 42.000 108.500 ;
        RECT 5.500 106.000 8.000 107.500 ;
        RECT 24.000 107.000 41.500 108.000 ;
        RECT 83.500 107.500 89.000 108.500 ;
        RECT 104.000 108.000 105.500 108.500 ;
        RECT 190.500 108.000 192.500 108.500 ;
        RECT 103.500 107.500 105.500 108.000 ;
        RECT 191.000 107.500 192.500 108.000 ;
        RECT 84.000 107.000 88.500 107.500 ;
        RECT 103.500 107.000 105.000 107.500 ;
        RECT 191.000 107.000 193.000 107.500 ;
        RECT 225.000 107.000 228.000 108.500 ;
        RECT 23.500 106.500 41.000 107.000 ;
        RECT 23.500 106.000 40.500 106.500 ;
        RECT 84.500 106.000 88.500 107.000 ;
        RECT 103.000 106.500 105.000 107.000 ;
        RECT 5.000 103.500 8.000 106.000 ;
        RECT 23.000 105.500 40.500 106.000 ;
        RECT 23.000 105.000 40.000 105.500 ;
        RECT 85.000 105.000 88.000 106.000 ;
        RECT 102.500 105.500 104.500 106.500 ;
        RECT 191.500 106.000 193.500 107.000 ;
        RECT 192.000 105.500 193.500 106.000 ;
        RECT 224.500 105.500 227.500 107.000 ;
        RECT 102.500 105.000 104.000 105.500 ;
        RECT 192.000 105.000 194.000 105.500 ;
        RECT 22.500 104.000 39.500 105.000 ;
        RECT 59.500 104.500 60.500 105.000 ;
        RECT 85.500 104.500 87.500 105.000 ;
        RECT 22.000 103.500 39.000 104.000 ;
        RECT 59.000 103.500 61.000 104.500 ;
        RECT 86.000 104.000 87.500 104.500 ;
        RECT 102.000 104.500 104.000 105.000 ;
        RECT 192.500 104.500 194.000 105.000 ;
        RECT 224.000 104.500 227.000 105.500 ;
        RECT 102.000 104.000 103.500 104.500 ;
        RECT 192.500 104.000 194.500 104.500 ;
        RECT 86.500 103.500 87.000 104.000 ;
        RECT 101.500 103.500 103.500 104.000 ;
        RECT 193.000 103.500 194.500 104.000 ;
        RECT 5.000 100.500 7.500 103.500 ;
        RECT 22.000 103.000 38.500 103.500 ;
        RECT 21.500 102.500 38.500 103.000 ;
        RECT 58.500 102.500 61.500 103.500 ;
        RECT 101.500 103.000 103.000 103.500 ;
        RECT 193.000 103.000 195.000 103.500 ;
        RECT 223.500 103.000 226.500 104.500 ;
        RECT 101.000 102.500 103.000 103.000 ;
        RECT 21.500 102.000 38.000 102.500 ;
        RECT 58.000 102.000 62.000 102.500 ;
        RECT 21.000 101.000 37.500 102.000 ;
        RECT 57.500 101.500 62.000 102.000 ;
        RECT 101.000 101.500 102.500 102.500 ;
        RECT 193.500 102.000 195.000 103.000 ;
        RECT 223.000 102.000 226.000 103.000 ;
        RECT 193.500 101.500 195.500 102.000 ;
        RECT 4.500 89.500 7.500 100.500 ;
        RECT 20.500 100.000 37.000 101.000 ;
        RECT 57.500 100.500 62.500 101.500 ;
        RECT 57.000 100.000 62.500 100.500 ;
        RECT 100.500 101.000 102.500 101.500 ;
        RECT 194.000 101.000 195.500 101.500 ;
        RECT 222.500 101.500 226.000 102.000 ;
        RECT 100.500 100.000 102.000 101.000 ;
        RECT 194.000 100.500 196.000 101.000 ;
        RECT 222.500 100.500 225.500 101.500 ;
        RECT 20.000 99.500 36.500 100.000 ;
        RECT 57.000 99.500 63.000 100.000 ;
        RECT 20.000 99.000 36.000 99.500 ;
        RECT 19.500 98.500 36.000 99.000 ;
        RECT 56.500 99.000 63.000 99.500 ;
        RECT 100.000 99.500 102.000 100.000 ;
        RECT 194.500 99.500 196.000 100.500 ;
        RECT 222.000 99.500 225.000 100.500 ;
        RECT 56.500 98.500 63.500 99.000 ;
        RECT 100.000 98.500 101.500 99.500 ;
        RECT 194.500 99.000 196.500 99.500 ;
        RECT 19.500 98.000 35.500 98.500 ;
        RECT 56.000 98.000 64.000 98.500 ;
        RECT 99.500 98.000 101.500 98.500 ;
        RECT 19.000 97.500 35.500 98.000 ;
        RECT 55.000 97.500 64.500 98.000 ;
        RECT 19.000 97.000 35.000 97.500 ;
        RECT 54.000 97.000 65.500 97.500 ;
        RECT 18.500 96.500 35.000 97.000 ;
        RECT 53.000 96.500 66.500 97.000 ;
        RECT 99.500 96.500 101.000 98.000 ;
        RECT 195.000 97.500 196.500 99.000 ;
        RECT 221.500 99.000 225.000 99.500 ;
        RECT 221.500 98.000 224.500 99.000 ;
        RECT 195.000 97.000 197.000 97.500 ;
        RECT 221.000 97.000 224.000 98.000 ;
        RECT 18.500 96.000 34.500 96.500 ;
        RECT 51.500 96.000 68.000 96.500 ;
        RECT 99.000 96.000 101.000 96.500 ;
        RECT 18.000 95.000 34.000 96.000 ;
        RECT 51.000 95.500 69.000 96.000 ;
        RECT 50.000 95.000 69.500 95.500 ;
        RECT 17.500 94.000 33.500 95.000 ;
        RECT 49.000 94.000 70.500 95.000 ;
        RECT 99.000 94.500 100.500 96.000 ;
        RECT 195.500 95.500 197.000 97.000 ;
        RECT 220.500 96.000 223.500 97.000 ;
        RECT 195.500 95.000 197.500 95.500 ;
        RECT 220.000 95.000 223.000 96.000 ;
        RECT 98.500 94.000 100.500 94.500 ;
        RECT 17.000 93.000 33.000 94.000 ;
        RECT 50.000 93.500 70.000 94.000 ;
        RECT 51.000 93.000 69.000 93.500 ;
        RECT 16.500 92.000 32.500 93.000 ;
        RECT 52.000 92.500 68.000 93.000 ;
        RECT 53.000 92.000 67.000 92.500 ;
        RECT 16.000 91.000 32.000 92.000 ;
        RECT 54.000 91.500 66.000 92.000 ;
        RECT 98.500 91.500 100.000 94.000 ;
        RECT 196.000 93.500 197.500 95.000 ;
        RECT 219.500 94.500 223.000 95.000 ;
        RECT 219.500 94.000 222.500 94.500 ;
        RECT 219.000 93.500 222.500 94.000 ;
        RECT 196.000 92.500 198.000 93.500 ;
        RECT 219.000 93.000 222.000 93.500 ;
        RECT 55.000 91.000 65.000 91.500 ;
        RECT 98.000 91.000 100.000 91.500 ;
        RECT 15.500 90.500 31.500 91.000 ;
        RECT 56.000 90.500 64.000 91.000 ;
        RECT 15.500 90.000 31.000 90.500 ;
        RECT 56.000 90.000 63.500 90.500 ;
        RECT 5.000 87.000 7.500 89.500 ;
        RECT 15.000 89.500 31.000 90.000 ;
        RECT 15.000 88.500 30.500 89.500 ;
        RECT 56.500 89.000 63.000 90.000 ;
        RECT 14.500 87.500 30.000 88.500 ;
        RECT 57.000 88.000 62.500 89.000 ;
        RECT 5.000 84.000 8.000 87.000 ;
        RECT 14.000 86.500 29.500 87.500 ;
        RECT 57.500 87.000 62.000 88.000 ;
        RECT 58.000 86.500 62.000 87.000 ;
        RECT 98.000 86.500 99.500 91.000 ;
        RECT 196.500 90.000 198.000 92.500 ;
        RECT 218.500 92.500 222.000 93.000 ;
        RECT 218.500 92.000 221.500 92.500 ;
        RECT 218.000 91.500 221.500 92.000 ;
        RECT 218.000 91.000 221.000 91.500 ;
        RECT 217.500 90.500 221.000 91.000 ;
        RECT 217.500 90.000 220.500 90.500 ;
        RECT 196.500 89.000 198.500 90.000 ;
        RECT 217.000 89.500 220.500 90.000 ;
        RECT 217.000 89.000 220.000 89.500 ;
        RECT 13.500 85.500 29.000 86.500 ;
        RECT 58.000 86.000 61.500 86.500 ;
        RECT 13.500 85.000 28.500 85.500 ;
        RECT 58.500 85.000 61.000 86.000 ;
        RECT 13.000 84.000 28.500 85.000 ;
        RECT 59.000 84.000 60.500 85.000 ;
        RECT 5.500 83.000 8.000 84.000 ;
        RECT 12.500 83.000 28.000 84.000 ;
        RECT 59.500 83.500 60.000 84.000 ;
        RECT 5.500 80.500 8.500 83.000 ;
        RECT 12.000 82.000 27.500 83.000 ;
        RECT 12.000 81.500 27.000 82.000 ;
        RECT 97.500 81.500 99.500 86.500 ;
        RECT 197.000 81.500 198.500 89.000 ;
        RECT 216.500 88.500 220.000 89.000 ;
        RECT 216.500 88.000 219.500 88.500 ;
        RECT 216.000 87.500 219.000 88.000 ;
        RECT 215.500 87.000 219.000 87.500 ;
        RECT 215.500 86.500 218.500 87.000 ;
        RECT 215.000 86.000 218.500 86.500 ;
        RECT 224.000 86.000 225.500 86.500 ;
        RECT 215.000 85.500 218.000 86.000 ;
        RECT 222.500 85.500 226.500 86.000 ;
        RECT 214.500 85.000 218.000 85.500 ;
        RECT 221.000 85.000 227.000 85.500 ;
        RECT 214.000 84.500 218.000 85.000 ;
        RECT 219.000 84.500 227.500 85.000 ;
        RECT 214.000 84.000 227.500 84.500 ;
        RECT 213.500 83.000 227.500 84.000 ;
        RECT 212.500 82.500 222.000 83.000 ;
        RECT 208.500 82.000 220.500 82.500 ;
        RECT 224.500 82.000 227.500 83.000 ;
        RECT 202.000 81.500 219.000 82.000 ;
        RECT 11.500 81.000 27.000 81.500 ;
        RECT 11.500 80.500 26.500 81.000 ;
        RECT 6.000 79.500 8.500 80.500 ;
        RECT 11.000 80.000 26.500 80.500 ;
        RECT 84.000 80.000 84.500 80.500 ;
        RECT 6.000 78.000 9.000 79.500 ;
        RECT 11.000 79.000 26.000 80.000 ;
        RECT 84.000 79.500 85.000 80.000 ;
        RECT 10.500 78.500 26.000 79.000 ;
        RECT 83.500 79.000 85.000 79.500 ;
        RECT 83.500 78.500 85.500 79.000 ;
        RECT 10.500 78.000 25.500 78.500 ;
        RECT 6.500 77.000 9.000 78.000 ;
        RECT 10.000 77.500 25.500 78.000 ;
        RECT 83.000 78.000 85.500 78.500 ;
        RECT 83.000 77.500 86.000 78.000 ;
        RECT 10.000 77.000 25.000 77.500 ;
        RECT 6.500 76.500 25.000 77.000 ;
        RECT 82.500 77.000 86.000 77.500 ;
        RECT 98.000 77.500 99.500 81.500 ;
        RECT 181.500 81.000 217.500 81.500 ;
        RECT 176.000 80.500 215.500 81.000 ;
        RECT 224.000 80.500 227.000 82.000 ;
        RECT 173.000 80.000 213.000 80.500 ;
        RECT 170.500 79.500 207.000 80.000 ;
        RECT 168.000 79.000 199.000 79.500 ;
        RECT 223.500 79.000 226.500 80.500 ;
        RECT 166.500 78.500 181.500 79.000 ;
        RECT 165.000 78.000 176.000 78.500 ;
        RECT 223.000 78.000 226.000 79.000 ;
        RECT 163.500 77.500 173.500 78.000 ;
        RECT 222.500 77.500 226.000 78.000 ;
        RECT 82.500 76.500 86.500 77.000 ;
        RECT 98.000 76.500 100.000 77.500 ;
        RECT 162.000 77.000 171.000 77.500 ;
        RECT 160.500 76.500 169.000 77.000 ;
        RECT 222.500 76.500 225.500 77.500 ;
        RECT 6.500 75.500 24.500 76.500 ;
        RECT 82.000 76.000 87.000 76.500 ;
        RECT 81.500 75.500 88.000 76.000 ;
        RECT 7.000 75.000 24.500 75.500 ;
        RECT 80.500 75.000 89.000 75.500 ;
        RECT 7.000 74.000 24.000 75.000 ;
        RECT 79.500 74.500 90.000 75.000 ;
        RECT 98.500 74.500 100.000 76.500 ;
        RECT 159.500 76.000 167.000 76.500 ;
        RECT 158.000 75.500 165.500 76.000 ;
        RECT 222.000 75.500 225.000 76.500 ;
        RECT 157.000 75.000 164.000 75.500 ;
        RECT 221.500 75.000 225.000 75.500 ;
        RECT 156.000 74.500 162.500 75.000 ;
        RECT 221.500 74.500 224.500 75.000 ;
        RECT 78.500 74.000 91.000 74.500 ;
        RECT 98.500 74.000 100.500 74.500 ;
        RECT 155.000 74.000 161.000 74.500 ;
        RECT 221.000 74.000 224.500 74.500 ;
        RECT 7.000 73.500 23.500 74.000 ;
        RECT 78.000 73.500 90.500 74.000 ;
        RECT 7.500 73.000 23.500 73.500 ;
        RECT 78.500 73.000 90.000 73.500 ;
        RECT 7.500 71.500 23.000 73.000 ;
        RECT 79.500 72.500 89.000 73.000 ;
        RECT 99.000 72.500 100.500 74.000 ;
        RECT 154.000 73.500 159.500 74.000 ;
        RECT 221.000 73.500 224.000 74.000 ;
        RECT 153.000 73.000 158.500 73.500 ;
        RECT 220.500 73.000 224.000 73.500 ;
        RECT 152.000 72.500 157.000 73.000 ;
        RECT 220.500 72.500 223.500 73.000 ;
        RECT 81.000 72.000 88.000 72.500 ;
        RECT 99.000 72.000 101.000 72.500 ;
        RECT 151.000 72.000 156.000 72.500 ;
        RECT 220.000 72.000 223.500 72.500 ;
        RECT 82.000 71.500 87.000 72.000 ;
        RECT 8.000 70.000 22.500 71.500 ;
        RECT 82.500 70.500 86.500 71.500 ;
        RECT 99.500 70.500 101.000 72.000 ;
        RECT 150.000 71.500 155.000 72.000 ;
        RECT 220.000 71.500 223.000 72.000 ;
        RECT 149.000 71.000 154.000 71.500 ;
        RECT 219.500 71.000 223.000 71.500 ;
        RECT 148.000 70.500 152.500 71.000 ;
        RECT 219.500 70.500 222.500 71.000 ;
        RECT 57.000 70.000 57.500 70.500 ;
        RECT 8.500 69.000 22.000 70.000 ;
        RECT 57.000 69.500 58.000 70.000 ;
        RECT 83.000 69.500 86.000 70.500 ;
        RECT 99.500 70.000 101.500 70.500 ;
        RECT 147.500 70.000 151.500 70.500 ;
        RECT 219.000 70.000 222.500 70.500 ;
        RECT 8.500 68.500 21.500 69.000 ;
        RECT 56.500 68.500 58.500 69.500 ;
        RECT 83.500 68.500 85.500 69.500 ;
        RECT 100.000 69.000 101.500 70.000 ;
        RECT 146.500 69.500 150.500 70.000 ;
        RECT 219.000 69.500 222.000 70.000 ;
        RECT 145.500 69.000 149.500 69.500 ;
        RECT 218.500 69.000 222.000 69.500 ;
        RECT 100.000 68.500 102.000 69.000 ;
        RECT 144.500 68.500 149.000 69.000 ;
        RECT 218.500 68.500 221.500 69.000 ;
        RECT 9.000 67.500 21.500 68.500 ;
        RECT 56.000 67.500 59.000 68.500 ;
        RECT 84.000 68.000 85.500 68.500 ;
        RECT 84.500 67.500 85.000 68.000 ;
        RECT 100.500 67.500 102.000 68.500 ;
        RECT 143.500 68.000 148.000 68.500 ;
        RECT 218.000 68.000 221.500 68.500 ;
        RECT 143.000 67.500 147.000 68.000 ;
        RECT 217.500 67.500 221.000 68.000 ;
        RECT 9.000 67.000 21.000 67.500 ;
        RECT 9.500 66.000 21.000 67.000 ;
        RECT 55.500 66.500 59.500 67.500 ;
        RECT 100.500 67.000 102.500 67.500 ;
        RECT 142.000 67.000 146.000 67.500 ;
        RECT 217.500 67.000 220.500 67.500 ;
        RECT 55.000 66.000 60.000 66.500 ;
        RECT 101.000 66.000 102.500 67.000 ;
        RECT 141.000 66.500 145.500 67.000 ;
        RECT 217.000 66.500 220.500 67.000 ;
        RECT 140.500 66.000 144.500 66.500 ;
        RECT 217.000 66.000 220.000 66.500 ;
        RECT 9.500 65.500 20.500 66.000 ;
        RECT 54.500 65.500 60.500 66.000 ;
        RECT 101.000 65.500 103.000 66.000 ;
        RECT 139.500 65.500 144.000 66.000 ;
        RECT 216.500 65.500 220.000 66.000 ;
        RECT 10.000 65.000 20.500 65.500 ;
        RECT 53.500 65.000 61.500 65.500 ;
        RECT 101.500 65.000 103.000 65.500 ;
        RECT 138.500 65.000 143.000 65.500 ;
        RECT 216.000 65.000 219.500 65.500 ;
        RECT 10.000 64.000 20.000 65.000 ;
        RECT 52.500 64.500 62.500 65.000 ;
        RECT 101.500 64.500 103.500 65.000 ;
        RECT 138.000 64.500 142.000 65.000 ;
        RECT 216.000 64.500 219.000 65.000 ;
        RECT 51.500 64.000 63.500 64.500 ;
        RECT 102.000 64.000 103.500 64.500 ;
        RECT 137.000 64.000 141.500 64.500 ;
        RECT 215.500 64.000 219.000 64.500 ;
        RECT 10.500 63.500 20.000 64.000 ;
        RECT 10.500 62.500 19.500 63.500 ;
        RECT 50.500 63.000 64.000 64.000 ;
        RECT 102.000 63.500 104.000 64.000 ;
        RECT 136.500 63.500 140.500 64.000 ;
        RECT 215.000 63.500 218.500 64.000 ;
        RECT 51.500 62.500 63.500 63.000 ;
        RECT 102.500 62.500 104.000 63.500 ;
        RECT 135.500 63.000 140.000 63.500 ;
        RECT 215.000 63.000 218.000 63.500 ;
        RECT 134.500 62.500 139.000 63.000 ;
        RECT 214.500 62.500 218.000 63.000 ;
        RECT 11.000 62.000 19.500 62.500 ;
        RECT 52.500 62.000 62.500 62.500 ;
        RECT 102.500 62.000 104.500 62.500 ;
        RECT 134.000 62.000 138.000 62.500 ;
        RECT 214.000 62.000 217.500 62.500 ;
        RECT 11.000 61.500 19.000 62.000 ;
        RECT 53.500 61.500 61.500 62.000 ;
        RECT 103.000 61.500 104.500 62.000 ;
        RECT 133.000 61.500 137.500 62.000 ;
        RECT 11.500 60.500 19.000 61.500 ;
        RECT 54.500 61.000 60.500 61.500 ;
        RECT 103.000 61.000 105.000 61.500 ;
        RECT 132.500 61.000 136.500 61.500 ;
        RECT 213.500 61.000 217.000 62.000 ;
        RECT 55.000 60.500 60.000 61.000 ;
        RECT 103.500 60.500 105.500 61.000 ;
        RECT 131.500 60.500 136.000 61.000 ;
        RECT 213.000 60.500 216.500 61.000 ;
        RECT 12.000 59.000 18.500 60.500 ;
        RECT 55.500 59.500 59.500 60.500 ;
        RECT 104.000 60.000 105.500 60.500 ;
        RECT 131.000 60.000 135.000 60.500 ;
        RECT 212.500 60.000 216.000 60.500 ;
        RECT 104.000 59.500 106.000 60.000 ;
        RECT 130.000 59.500 134.500 60.000 ;
        RECT 212.000 59.500 215.500 60.000 ;
        RECT 12.500 58.000 18.000 59.000 ;
        RECT 56.000 58.500 59.000 59.500 ;
        RECT 104.500 59.000 106.000 59.500 ;
        RECT 129.500 59.000 133.500 59.500 ;
        RECT 211.500 59.000 215.500 59.500 ;
        RECT 104.500 58.500 106.500 59.000 ;
        RECT 128.500 58.500 132.500 59.000 ;
        RECT 211.500 58.500 215.000 59.000 ;
        RECT 13.000 57.500 18.000 58.000 ;
        RECT 56.500 57.500 58.500 58.500 ;
        RECT 105.000 58.000 106.500 58.500 ;
        RECT 128.000 58.000 132.000 58.500 ;
        RECT 211.000 58.000 214.500 58.500 ;
        RECT 105.000 57.500 107.000 58.000 ;
        RECT 127.000 57.500 131.000 58.000 ;
        RECT 210.500 57.500 214.000 58.000 ;
        RECT 13.000 57.000 17.500 57.500 ;
        RECT 13.500 56.000 17.500 57.000 ;
        RECT 57.000 57.000 58.000 57.500 ;
        RECT 105.500 57.000 107.500 57.500 ;
        RECT 126.500 57.000 130.500 57.500 ;
        RECT 210.000 57.000 213.500 57.500 ;
        RECT 57.000 56.500 57.500 57.000 ;
        RECT 106.000 56.500 107.500 57.000 ;
        RECT 125.500 56.500 129.500 57.000 ;
        RECT 209.500 56.500 213.500 57.000 ;
        RECT 106.000 56.000 108.000 56.500 ;
        RECT 125.000 56.000 129.000 56.500 ;
        RECT 209.000 56.000 213.000 56.500 ;
        RECT 14.000 55.000 17.500 56.000 ;
        RECT 14.500 54.500 17.500 55.000 ;
        RECT 106.500 55.500 108.500 56.000 ;
        RECT 124.000 55.500 128.000 56.000 ;
        RECT 208.500 55.500 212.500 56.000 ;
        RECT 106.500 54.500 109.000 55.500 ;
        RECT 123.500 55.000 127.000 55.500 ;
        RECT 208.000 55.000 212.000 55.500 ;
        RECT 123.000 54.500 126.500 55.000 ;
        RECT 208.000 54.500 211.500 55.000 ;
        RECT 14.500 54.000 18.000 54.500 ;
        RECT 106.000 54.000 109.500 54.500 ;
        RECT 122.000 54.000 126.000 54.500 ;
        RECT 207.500 54.000 211.000 54.500 ;
        RECT 15.000 53.500 18.000 54.000 ;
        RECT 105.500 53.500 110.000 54.000 ;
        RECT 121.500 53.500 125.000 54.000 ;
        RECT 207.000 53.500 210.500 54.000 ;
        RECT 15.000 53.000 18.500 53.500 ;
        RECT 15.500 52.500 18.500 53.000 ;
        RECT 105.000 53.000 110.500 53.500 ;
        RECT 120.500 53.000 124.500 53.500 ;
        RECT 206.500 53.000 210.000 53.500 ;
        RECT 105.000 52.500 107.500 53.000 ;
        RECT 108.500 52.500 110.500 53.000 ;
        RECT 120.000 52.500 123.500 53.000 ;
        RECT 206.000 52.500 210.000 53.000 ;
        RECT 16.000 52.000 19.000 52.500 ;
        RECT 104.500 52.000 107.000 52.500 ;
        RECT 109.000 52.000 111.000 52.500 ;
        RECT 119.000 52.000 123.000 52.500 ;
        RECT 205.500 52.000 209.500 52.500 ;
        RECT 16.000 51.500 19.500 52.000 ;
        RECT 104.000 51.500 106.500 52.000 ;
        RECT 109.500 51.500 111.500 52.000 ;
        RECT 118.500 51.500 122.000 52.000 ;
        RECT 205.000 51.500 209.000 52.000 ;
        RECT 16.500 51.000 19.500 51.500 ;
        RECT 103.500 51.000 106.000 51.500 ;
        RECT 110.000 51.000 112.000 51.500 ;
        RECT 118.000 51.000 121.500 51.500 ;
        RECT 204.500 51.000 208.500 51.500 ;
        RECT 16.500 50.500 20.000 51.000 ;
        RECT 103.000 50.500 105.500 51.000 ;
        RECT 110.500 50.500 112.500 51.000 ;
        RECT 117.000 50.500 120.500 51.000 ;
        RECT 204.000 50.500 208.000 51.000 ;
        RECT 17.000 50.000 20.000 50.500 ;
        RECT 102.500 50.000 105.000 50.500 ;
        RECT 111.000 50.000 113.000 50.500 ;
        RECT 116.500 50.000 120.000 50.500 ;
        RECT 203.000 50.000 207.500 50.500 ;
        RECT 17.000 49.500 20.500 50.000 ;
        RECT 102.000 49.500 105.000 50.000 ;
        RECT 111.500 49.500 113.500 50.000 ;
        RECT 115.500 49.500 119.000 50.000 ;
        RECT 202.500 49.500 207.000 50.000 ;
        RECT 17.500 49.000 21.000 49.500 ;
        RECT 101.500 49.000 104.500 49.500 ;
        RECT 111.500 49.000 114.000 49.500 ;
        RECT 115.000 49.000 118.500 49.500 ;
        RECT 202.000 49.000 206.500 49.500 ;
        RECT 18.000 48.500 21.000 49.000 ;
        RECT 101.000 48.500 104.000 49.000 ;
        RECT 112.000 48.500 117.500 49.000 ;
        RECT 201.500 48.500 206.000 49.000 ;
        RECT 18.000 48.000 21.500 48.500 ;
        RECT 101.000 48.000 103.500 48.500 ;
        RECT 112.500 48.000 117.000 48.500 ;
        RECT 201.000 48.000 205.000 48.500 ;
        RECT 18.500 47.500 22.000 48.000 ;
        RECT 100.500 47.500 103.000 48.000 ;
        RECT 112.500 47.500 116.000 48.000 ;
        RECT 200.500 47.500 204.500 48.000 ;
        RECT 19.000 47.000 22.000 47.500 ;
        RECT 100.000 47.000 102.500 47.500 ;
        RECT 112.000 47.000 115.500 47.500 ;
        RECT 200.000 47.000 204.000 47.500 ;
        RECT 19.000 46.500 22.500 47.000 ;
        RECT 99.500 46.500 102.000 47.000 ;
        RECT 111.500 46.500 114.500 47.000 ;
        RECT 199.500 46.500 203.500 47.000 ;
        RECT 19.500 46.000 23.000 46.500 ;
        RECT 99.000 46.000 101.500 46.500 ;
        RECT 110.500 46.000 114.000 46.500 ;
        RECT 198.500 46.000 203.000 46.500 ;
        RECT 20.000 45.500 23.000 46.000 ;
        RECT 98.500 45.500 101.000 46.000 ;
        RECT 110.000 45.500 113.000 46.000 ;
        RECT 198.000 45.500 202.500 46.000 ;
        RECT 20.000 45.000 23.500 45.500 ;
        RECT 98.000 45.000 100.500 45.500 ;
        RECT 109.000 45.000 112.500 45.500 ;
        RECT 197.500 45.000 202.000 45.500 ;
        RECT 20.500 44.500 24.000 45.000 ;
        RECT 97.500 44.500 100.000 45.000 ;
        RECT 108.500 44.500 111.500 45.000 ;
        RECT 197.000 44.500 201.500 45.000 ;
        RECT 21.000 43.500 24.500 44.500 ;
        RECT 97.000 44.000 99.500 44.500 ;
        RECT 107.500 44.000 111.000 44.500 ;
        RECT 196.000 44.000 200.500 44.500 ;
        RECT 96.500 43.500 99.500 44.000 ;
        RECT 107.000 43.500 110.000 44.000 ;
        RECT 195.500 43.500 200.000 44.000 ;
        RECT 21.500 43.000 25.000 43.500 ;
        RECT 96.000 43.000 99.000 43.500 ;
        RECT 106.500 43.000 109.500 43.500 ;
        RECT 195.000 43.000 199.500 43.500 ;
        RECT 22.000 42.500 25.500 43.000 ;
        RECT 96.000 42.500 98.500 43.000 ;
        RECT 105.500 42.500 108.500 43.000 ;
        RECT 194.000 42.500 199.000 43.000 ;
        RECT 22.500 42.000 26.000 42.500 ;
        RECT 95.500 42.000 98.000 42.500 ;
        RECT 105.000 42.000 108.000 42.500 ;
        RECT 193.500 42.000 198.000 42.500 ;
        RECT 22.500 41.500 26.500 42.000 ;
        RECT 95.000 41.500 97.500 42.000 ;
        RECT 104.000 41.500 107.000 42.000 ;
        RECT 193.000 41.500 197.500 42.000 ;
        RECT 23.000 41.000 26.500 41.500 ;
        RECT 94.500 41.000 97.000 41.500 ;
        RECT 103.500 41.000 106.500 41.500 ;
        RECT 192.000 41.000 197.000 41.500 ;
        RECT 23.500 40.500 27.000 41.000 ;
        RECT 94.000 40.500 96.500 41.000 ;
        RECT 102.500 40.500 105.500 41.000 ;
        RECT 191.500 40.500 196.000 41.000 ;
        RECT 24.000 40.000 27.500 40.500 ;
        RECT 93.500 40.000 96.000 40.500 ;
        RECT 101.500 40.000 105.000 40.500 ;
        RECT 190.500 40.000 195.500 40.500 ;
        RECT 24.500 39.500 28.000 40.000 ;
        RECT 93.000 39.500 95.500 40.000 ;
        RECT 101.000 39.500 104.000 40.000 ;
        RECT 190.000 39.500 195.000 40.000 ;
        RECT 24.500 39.000 28.500 39.500 ;
        RECT 92.500 39.000 95.000 39.500 ;
        RECT 100.000 39.000 103.500 39.500 ;
        RECT 189.000 39.000 194.000 39.500 ;
        RECT 25.000 38.500 29.000 39.000 ;
        RECT 92.000 38.500 94.500 39.000 ;
        RECT 99.500 38.500 102.500 39.000 ;
        RECT 188.500 38.500 193.500 39.000 ;
        RECT 25.500 38.000 29.500 38.500 ;
        RECT 91.500 38.000 94.000 38.500 ;
        RECT 98.500 38.000 102.000 38.500 ;
        RECT 187.500 38.000 192.500 38.500 ;
        RECT 26.000 37.500 30.000 38.000 ;
        RECT 91.000 37.500 93.500 38.000 ;
        RECT 98.000 37.500 101.000 38.000 ;
        RECT 187.000 37.500 192.000 38.000 ;
        RECT 26.500 37.000 30.500 37.500 ;
        RECT 90.500 37.000 93.000 37.500 ;
        RECT 97.000 37.000 100.000 37.500 ;
        RECT 186.000 37.000 191.000 37.500 ;
        RECT 27.000 36.500 31.000 37.000 ;
        RECT 27.500 36.000 31.000 36.500 ;
        RECT 90.000 36.500 92.500 37.000 ;
        RECT 96.500 36.500 99.500 37.000 ;
        RECT 185.000 36.500 190.500 37.000 ;
        RECT 90.000 36.000 92.000 36.500 ;
        RECT 95.500 36.000 99.000 36.500 ;
        RECT 184.500 36.000 189.500 36.500 ;
        RECT 28.000 35.500 31.500 36.000 ;
        RECT 89.500 35.500 92.000 36.000 ;
        RECT 94.500 35.500 98.000 36.000 ;
        RECT 183.500 35.500 189.000 36.000 ;
        RECT 28.500 35.000 32.000 35.500 ;
        RECT 89.000 35.000 91.500 35.500 ;
        RECT 94.000 35.000 97.500 35.500 ;
        RECT 182.500 35.000 188.000 35.500 ;
        RECT 29.000 34.500 32.500 35.000 ;
        RECT 88.500 34.500 91.000 35.000 ;
        RECT 93.000 34.500 96.500 35.000 ;
        RECT 182.000 34.500 187.500 35.000 ;
        RECT 29.500 34.000 33.000 34.500 ;
        RECT 88.000 34.000 90.500 34.500 ;
        RECT 92.000 34.000 96.000 34.500 ;
        RECT 181.000 34.000 186.500 34.500 ;
        RECT 30.000 33.500 34.000 34.000 ;
        RECT 87.500 33.500 90.500 34.000 ;
        RECT 91.500 33.500 95.000 34.000 ;
        RECT 180.000 33.500 185.500 34.000 ;
        RECT 30.500 33.000 34.500 33.500 ;
        RECT 87.000 33.000 94.500 33.500 ;
        RECT 179.500 33.000 185.000 33.500 ;
        RECT 30.500 32.500 35.000 33.000 ;
        RECT 86.500 32.500 93.500 33.000 ;
        RECT 178.500 32.500 184.000 33.000 ;
        RECT 31.500 32.000 35.500 32.500 ;
        RECT 86.000 32.000 93.000 32.500 ;
        RECT 177.500 32.000 183.000 32.500 ;
        RECT 32.000 31.500 36.000 32.000 ;
        RECT 85.500 31.500 92.000 32.000 ;
        RECT 176.500 31.500 182.500 32.000 ;
        RECT 32.500 31.000 36.500 31.500 ;
        RECT 85.000 31.000 91.500 31.500 ;
        RECT 175.500 31.000 181.500 31.500 ;
        RECT 33.000 30.500 37.000 31.000 ;
        RECT 84.500 30.500 90.500 31.000 ;
        RECT 174.500 30.500 180.500 31.000 ;
        RECT 33.500 30.000 37.500 30.500 ;
        RECT 84.000 30.000 90.000 30.500 ;
        RECT 173.500 30.000 179.500 30.500 ;
        RECT 34.000 29.500 38.500 30.000 ;
        RECT 83.500 29.500 89.000 30.000 ;
        RECT 172.500 29.500 178.500 30.000 ;
        RECT 34.500 29.000 39.000 29.500 ;
        RECT 83.000 29.000 88.000 29.500 ;
        RECT 171.500 29.000 177.500 29.500 ;
        RECT 35.000 28.500 39.500 29.000 ;
        RECT 82.500 28.500 87.500 29.000 ;
        RECT 170.500 28.500 177.000 29.000 ;
        RECT 35.500 28.000 40.000 28.500 ;
        RECT 82.000 28.000 86.500 28.500 ;
        RECT 169.500 28.000 176.000 28.500 ;
        RECT 36.500 27.500 41.000 28.000 ;
        RECT 81.500 27.500 85.500 28.000 ;
        RECT 168.500 27.500 175.000 28.000 ;
        RECT 37.000 27.000 41.500 27.500 ;
        RECT 80.500 27.000 85.000 27.500 ;
        RECT 167.000 27.000 174.000 27.500 ;
        RECT 37.500 26.500 42.500 27.000 ;
        RECT 79.500 26.500 84.000 27.000 ;
        RECT 166.000 26.500 172.500 27.000 ;
        RECT 38.000 26.000 43.000 26.500 ;
        RECT 78.500 26.000 83.000 26.500 ;
        RECT 165.000 26.000 171.500 26.500 ;
        RECT 39.000 25.500 43.500 26.000 ;
        RECT 77.500 25.500 82.500 26.000 ;
        RECT 163.500 25.500 170.500 26.000 ;
        RECT 39.500 25.000 44.500 25.500 ;
        RECT 77.000 25.000 81.500 25.500 ;
        RECT 162.500 25.000 169.500 25.500 ;
        RECT 40.000 24.500 45.000 25.000 ;
        RECT 76.000 24.500 80.500 25.000 ;
        RECT 161.500 24.500 168.500 25.000 ;
        RECT 41.000 24.000 46.000 24.500 ;
        RECT 75.000 24.000 79.500 24.500 ;
        RECT 160.000 24.000 167.500 24.500 ;
        RECT 41.500 23.500 46.500 24.000 ;
        RECT 74.000 23.500 78.500 24.000 ;
        RECT 159.000 23.500 166.000 24.000 ;
        RECT 42.500 23.000 47.500 23.500 ;
        RECT 73.000 23.000 78.000 23.500 ;
        RECT 157.500 23.000 165.000 23.500 ;
        RECT 43.000 22.500 48.500 23.000 ;
        RECT 72.000 22.500 77.000 23.000 ;
        RECT 156.500 22.500 164.000 23.000 ;
        RECT 44.000 22.000 49.000 22.500 ;
        RECT 71.500 22.000 76.000 22.500 ;
        RECT 155.000 22.000 162.500 22.500 ;
        RECT 44.500 21.500 50.000 22.000 ;
        RECT 70.500 21.500 75.000 22.000 ;
        RECT 153.500 21.500 161.500 22.000 ;
        RECT 45.500 21.000 51.000 21.500 ;
        RECT 69.500 21.000 74.000 21.500 ;
        RECT 152.000 21.000 160.000 21.500 ;
        RECT 46.000 20.500 52.000 21.000 ;
        RECT 68.500 20.500 73.000 21.000 ;
        RECT 151.000 20.500 159.000 21.000 ;
        RECT 47.000 20.000 53.000 20.500 ;
        RECT 67.500 20.000 72.000 20.500 ;
        RECT 149.500 20.000 157.500 20.500 ;
        RECT 48.000 19.500 53.500 20.000 ;
        RECT 66.500 19.500 71.000 20.000 ;
        RECT 148.000 19.500 156.000 20.000 ;
        RECT 48.500 19.000 55.000 19.500 ;
        RECT 65.500 19.000 70.000 19.500 ;
        RECT 146.500 19.000 155.000 19.500 ;
        RECT 49.500 18.500 56.000 19.000 ;
        RECT 64.500 18.500 69.500 19.000 ;
        RECT 145.000 18.500 153.500 19.000 ;
        RECT 50.500 18.000 57.000 18.500 ;
        RECT 63.500 18.000 68.500 18.500 ;
        RECT 143.000 18.000 152.000 18.500 ;
        RECT 51.500 17.500 58.000 18.000 ;
        RECT 62.500 17.500 67.500 18.000 ;
        RECT 141.500 17.500 150.500 18.000 ;
        RECT 52.500 17.000 59.500 17.500 ;
        RECT 61.500 17.000 66.500 17.500 ;
        RECT 140.000 17.000 149.000 17.500 ;
        RECT 53.500 16.500 65.500 17.000 ;
        RECT 138.000 16.500 147.500 17.000 ;
        RECT 54.500 16.000 64.000 16.500 ;
        RECT 136.500 16.000 146.000 16.500 ;
        RECT 55.500 15.500 63.000 16.000 ;
        RECT 134.500 15.500 144.500 16.000 ;
        RECT 55.500 15.000 62.000 15.500 ;
        RECT 133.000 15.000 143.000 15.500 ;
        RECT 54.500 14.500 61.000 15.000 ;
        RECT 131.000 14.500 141.500 15.000 ;
        RECT 53.000 14.000 60.000 14.500 ;
        RECT 128.500 14.000 139.500 14.500 ;
        RECT 52.000 13.500 59.000 14.000 ;
        RECT 126.500 13.500 138.000 14.000 ;
        RECT 51.000 13.000 58.000 13.500 ;
        RECT 124.000 13.000 136.000 13.500 ;
        RECT 50.000 12.500 57.000 13.000 ;
        RECT 121.500 12.500 134.500 13.000 ;
        RECT 48.500 12.000 55.500 12.500 ;
        RECT 118.500 12.000 132.500 12.500 ;
        RECT 47.500 11.500 54.500 12.000 ;
        RECT 115.500 11.500 130.500 12.000 ;
        RECT 46.000 11.000 53.500 11.500 ;
        RECT 110.500 11.000 128.500 11.500 ;
        RECT 45.000 10.500 52.000 11.000 ;
        RECT 102.000 10.500 126.000 11.000 ;
        RECT 43.500 10.000 51.000 10.500 ;
        RECT 89.000 10.000 123.500 10.500 ;
        RECT 42.500 9.500 50.000 10.000 ;
        RECT 66.500 9.500 121.000 10.000 ;
        RECT 41.000 9.000 49.000 9.500 ;
        RECT 61.500 9.000 118.000 9.500 ;
        RECT 39.500 8.500 47.500 9.000 ;
        RECT 58.000 8.500 114.000 9.000 ;
        RECT 38.000 8.000 46.500 8.500 ;
        RECT 54.500 8.000 108.500 8.500 ;
        RECT 36.500 7.500 45.000 8.000 ;
        RECT 51.500 7.500 96.000 8.000 ;
        RECT 35.500 7.000 43.500 7.500 ;
        RECT 48.500 7.000 71.500 7.500 ;
        RECT 35.000 6.500 42.500 7.000 ;
        RECT 46.000 6.500 64.500 7.000 ;
        RECT 34.500 6.000 42.500 6.500 ;
        RECT 43.500 6.000 60.000 6.500 ;
        RECT 34.500 5.500 56.500 6.000 ;
        RECT 34.500 5.000 53.500 5.500 ;
        RECT 34.500 4.500 50.500 5.000 ;
        RECT 34.500 4.000 48.000 4.500 ;
        RECT 34.500 3.500 45.500 4.000 ;
        RECT 35.000 3.000 43.000 3.500 ;
        RECT 35.500 2.500 40.500 3.000 ;
        RECT 36.000 2.000 38.000 2.500 ;
  END
END aef2
END LIBRARY

