* NGSPICE file created from test_counter.ext - technology: gf180mcuD
.subckt test_counter VDD VSS clk counter[0] counter[10] counter[11] counter[1] counter[2]
+ counter[3] counter[4] counter[5] counter[6] counter[7] counter[8] counter[9] rst
XFILLER_5_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_66_ net10 _31_ net11 _33_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_49_ _12_ _16_ _17_ _23_ _24_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_12_Left_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput7 net7 counter[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Left_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_65_ net10 _31_ _32_ _09_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_48_ net13 net14 net4 _23_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput10 net10 counter[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput8 net8 counter[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_12_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_81_ _11_ net1 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_47_ net14 _20_ net4 _22_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_64_ net10 _31_ _14_ _32_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_8_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput11 net11 counter[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput9 net9 counter[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_80_ _10_ net15 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_63_ net2 _30_ _31_ _08_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_46_ net14 _20_ _21_ _01_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput12 net12 counter[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_12_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_62_ net8 net9 _15_ _31_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_4_Left_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_45_ net14 _20_ _14_ _21_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput13 net13 counter[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_12_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_61_ net8 _15_ net9 _30_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_44_ net2 _19_ _20_ _00_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput14 net14 counter[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_60_ _29_ _07_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_43_ _12_ _13_ _16_ _17_ _20_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_42_ net12 _18_ net13 _19_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_41_ _16_ _17_ _18_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_11_Left_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_40_ net8 net9 net10 net11 _17_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Left_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 clk net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput2 rst net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_79_ _09_ net15 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_0_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_78_ _08_ net15 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_77_ _07_ net15 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_9_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout15 net1 net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_76_ _06_ net15 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_59_ net8 _15_ _28_ _29_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_10_Left_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_75_ _05_ net15 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_4_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_58_ net8 _15_ net2 _28_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_74_ _04_ net15 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_57_ net2 _15_ _27_ _06_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_56_ net3 net6 net7 _27_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_73_ _03_ net1 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_39_ net3 net6 net7 _16_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_2_Left_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_72_ _02_ net15 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_55_ net3 net6 _26_ _05_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_38_ net3 net6 net7 _15_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_54_ net3 net6 _14_ _26_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_71_ _01_ net15 net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_37_ net2 _14_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_8_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_70_ _00_ net15 net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_53_ net3 net2 _04_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_36_ net13 _13_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_52_ net5 _24_ _25_ _03_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_35_ net12 _12_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_6_Left_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_9_Left_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_51_ net5 _24_ _14_ _25_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_50_ net2 _22_ _24_ _02_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Left_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_8_Left_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput3 net3 counter[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XTAP_TAPCELL_ROW_12_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_69_ net12 _18_ _34_ _11_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput4 net4 counter[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_12_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_68_ net12 _18_ _14_ _34_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_5_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput5 net5 counter[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_12_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_67_ net2 _18_ _33_ _10_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput6 net6 counter[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_6_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

