magic
tech gf180mcuD
magscale 1 10
timestamp 1763231934
<< pwell >>
rect -344 -566 344 566
<< mvpsubdiff >>
rect -312 462 312 534
rect -312 418 -240 462
rect -312 23 -299 418
rect -253 23 -240 418
rect 240 418 312 462
rect -312 -462 -240 23
rect 240 -418 253 418
rect 299 -418 312 418
rect 240 -462 312 -418
rect -312 -534 312 -462
<< mvpsubdiffcont >>
rect -299 23 -253 418
rect 253 -418 299 418
<< polysilicon >>
rect -100 309 100 322
rect -100 263 -87 309
rect 87 263 100 309
rect -100 200 100 263
rect -100 -263 100 -200
rect -100 -309 -87 -263
rect 87 -309 100 -263
rect -100 -322 100 -309
<< polycontact >>
rect -87 263 87 309
rect -87 -309 87 -263
<< mvnhighres >>
rect -100 -200 100 200
<< metal1 >>
rect -299 418 -253 521
rect 253 418 299 521
rect -98 263 -87 309
rect 87 263 98 309
rect -299 12 -253 23
rect -98 -309 -87 -263
rect 87 -309 98 -263
rect 253 -521 299 -418
<< properties >>
string FIXED_BBOX -276 -498 276 498
string gencell ppolyf_u_1k_6p0
string library gf180mcu
string parameters w 1.0 l 2.0 m 1 nx 1 wmin 1.000 lmin 1.000 class resistor rho 1000 val 2.0k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
