VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aef2
  CLASS BLOCK ;
  FOREIGN aef2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 247.500 BY 235.500 ;
  OBS
      LAYER Metal5 ;
        RECT 231.500 229.000 232.500 229.500 ;
        RECT 231.000 228.000 232.500 229.000 ;
        RECT 230.500 227.500 232.500 228.000 ;
        RECT 230.000 227.000 232.500 227.500 ;
        RECT 230.000 226.500 233.000 227.000 ;
        RECT 229.500 226.000 233.000 226.500 ;
        RECT 229.000 225.500 233.000 226.000 ;
        RECT 228.500 224.500 233.000 225.500 ;
        RECT 228.000 224.000 233.000 224.500 ;
        RECT 227.500 223.500 233.500 224.000 ;
        RECT 227.000 223.000 233.500 223.500 ;
        RECT 226.500 222.500 233.500 223.000 ;
        RECT 226.000 222.000 233.500 222.500 ;
        RECT 225.500 221.000 233.500 222.000 ;
        RECT 225.000 220.500 234.000 221.000 ;
        RECT 224.500 220.000 234.000 220.500 ;
        RECT 223.500 219.500 234.000 220.000 ;
        RECT 223.000 219.000 234.000 219.500 ;
        RECT 222.500 218.500 234.000 219.000 ;
        RECT 222.000 218.000 234.000 218.500 ;
        RECT 221.500 217.500 234.000 218.000 ;
        RECT 220.500 217.000 234.000 217.500 ;
        RECT 220.000 216.500 234.500 217.000 ;
        RECT 219.500 216.000 234.500 216.500 ;
        RECT 218.500 215.500 234.500 216.000 ;
        RECT 218.000 215.000 234.500 215.500 ;
        RECT 217.000 214.500 234.500 215.000 ;
        RECT 216.500 214.000 234.500 214.500 ;
        RECT 215.500 213.500 234.500 214.000 ;
        RECT 214.500 213.000 234.500 213.500 ;
        RECT 213.500 212.500 235.000 213.000 ;
        RECT 213.000 212.000 235.000 212.500 ;
        RECT 212.000 211.500 235.000 212.000 ;
        RECT 211.000 211.000 235.000 211.500 ;
        RECT 210.000 210.500 235.000 211.000 ;
        RECT 208.500 210.000 235.000 210.500 ;
        RECT 207.500 209.500 235.000 210.000 ;
        RECT 206.500 209.000 235.000 209.500 ;
        RECT 205.500 208.500 235.000 209.000 ;
        RECT 204.000 208.000 235.000 208.500 ;
        RECT 203.000 207.500 235.000 208.000 ;
        RECT 201.500 207.000 235.000 207.500 ;
        RECT 200.500 206.500 235.500 207.000 ;
        RECT 199.000 206.000 235.500 206.500 ;
        RECT 198.000 205.500 235.500 206.000 ;
        RECT 196.500 205.000 235.500 205.500 ;
        RECT 195.500 204.500 235.500 205.000 ;
        RECT 194.500 204.000 235.500 204.500 ;
        RECT 193.000 203.500 235.500 204.000 ;
        RECT 192.000 203.000 235.500 203.500 ;
        RECT 190.500 202.500 235.500 203.000 ;
        RECT 189.500 202.000 235.500 202.500 ;
        RECT 188.500 201.500 235.500 202.000 ;
        RECT 187.500 201.000 235.500 201.500 ;
        RECT 186.500 200.500 235.500 201.000 ;
        RECT 185.500 200.000 235.500 200.500 ;
        RECT 184.500 199.500 235.500 200.000 ;
        RECT 183.500 199.000 235.500 199.500 ;
        RECT 182.500 198.500 235.500 199.000 ;
        RECT 182.000 198.000 235.500 198.500 ;
        RECT 181.000 197.500 235.500 198.000 ;
        RECT 180.000 197.000 235.500 197.500 ;
        RECT 179.500 196.500 235.500 197.000 ;
        RECT 178.500 196.000 235.500 196.500 ;
        RECT 177.500 195.500 235.500 196.000 ;
        RECT 177.000 195.000 235.500 195.500 ;
        RECT 176.500 194.500 235.500 195.000 ;
        RECT 175.500 194.000 235.500 194.500 ;
        RECT 175.000 193.500 235.500 194.000 ;
        RECT 174.000 193.000 235.500 193.500 ;
        RECT 173.500 192.500 235.500 193.000 ;
        RECT 173.000 192.000 235.500 192.500 ;
        RECT 172.000 191.500 235.500 192.000 ;
        RECT 171.500 191.000 235.500 191.500 ;
        RECT 171.000 190.500 235.500 191.000 ;
        RECT 170.500 190.000 235.500 190.500 ;
        RECT 169.500 189.500 235.500 190.000 ;
        RECT 169.000 189.000 235.500 189.500 ;
        RECT 168.500 188.500 235.500 189.000 ;
        RECT 87.000 188.000 104.500 188.500 ;
        RECT 168.000 188.000 235.500 188.500 ;
        RECT 83.000 187.500 108.500 188.000 ;
        RECT 167.500 187.500 235.500 188.000 ;
        RECT 80.000 187.000 111.500 187.500 ;
        RECT 167.000 187.000 235.000 187.500 ;
        RECT 77.000 186.500 114.000 187.000 ;
        RECT 166.500 186.500 235.000 187.000 ;
        RECT 75.000 186.000 116.000 186.500 ;
        RECT 166.000 186.000 235.000 186.500 ;
        RECT 73.000 185.500 118.000 186.000 ;
        RECT 165.500 185.500 235.000 186.000 ;
        RECT 71.000 185.000 120.000 185.500 ;
        RECT 165.000 185.000 235.000 185.500 ;
        RECT 69.500 184.500 119.500 185.000 ;
        RECT 164.500 184.500 235.000 185.000 ;
        RECT 68.000 184.000 117.000 184.500 ;
        RECT 164.000 184.000 235.000 184.500 ;
        RECT 66.500 183.500 115.000 184.000 ;
        RECT 163.500 183.500 235.000 184.000 ;
        RECT 65.000 183.000 113.000 183.500 ;
        RECT 163.000 183.000 235.000 183.500 ;
        RECT 64.000 182.500 111.500 183.000 ;
        RECT 162.500 182.500 235.000 183.000 ;
        RECT 62.500 182.000 109.500 182.500 ;
        RECT 162.000 182.000 235.000 182.500 ;
        RECT 61.000 181.500 107.500 182.000 ;
        RECT 162.000 181.500 234.500 182.000 ;
        RECT 60.000 181.000 106.000 181.500 ;
        RECT 161.500 181.000 234.500 181.500 ;
        RECT 59.000 180.500 104.500 181.000 ;
        RECT 161.000 180.500 234.500 181.000 ;
        RECT 58.000 180.000 102.500 180.500 ;
        RECT 160.500 180.000 234.500 180.500 ;
        RECT 57.000 179.500 101.000 180.000 ;
        RECT 160.000 179.500 234.500 180.000 ;
        RECT 56.000 179.000 99.500 179.500 ;
        RECT 55.000 178.500 98.000 179.000 ;
        RECT 159.500 178.500 234.500 179.500 ;
        RECT 54.000 178.000 97.000 178.500 ;
        RECT 159.000 178.000 234.000 178.500 ;
        RECT 53.000 177.500 95.500 178.000 ;
        RECT 158.500 177.500 234.000 178.000 ;
        RECT 52.000 177.000 94.000 177.500 ;
        RECT 158.000 177.000 234.000 177.500 ;
        RECT 51.000 176.500 93.000 177.000 ;
        RECT 137.000 176.500 140.000 177.000 ;
        RECT 50.500 176.000 91.500 176.500 ;
        RECT 135.000 176.000 141.000 176.500 ;
        RECT 157.500 176.000 234.000 177.000 ;
        RECT 49.500 175.500 90.500 176.000 ;
        RECT 132.500 175.500 141.500 176.000 ;
        RECT 157.000 175.500 234.000 176.000 ;
        RECT 48.500 175.000 89.000 175.500 ;
        RECT 130.500 175.000 142.500 175.500 ;
        RECT 156.500 175.000 234.000 175.500 ;
        RECT 48.000 174.500 88.000 175.000 ;
        RECT 129.000 174.500 143.000 175.000 ;
        RECT 47.000 174.000 87.000 174.500 ;
        RECT 127.000 174.000 144.000 174.500 ;
        RECT 156.000 174.000 233.500 175.000 ;
        RECT 46.500 173.500 86.000 174.000 ;
        RECT 125.000 173.500 144.500 174.000 ;
        RECT 155.500 173.500 233.500 174.000 ;
        RECT 45.500 173.000 85.000 173.500 ;
        RECT 123.500 173.000 145.500 173.500 ;
        RECT 45.000 172.500 84.000 173.000 ;
        RECT 122.000 172.500 146.000 173.000 ;
        RECT 155.000 172.500 233.500 173.500 ;
        RECT 44.500 172.000 83.000 172.500 ;
        RECT 120.500 172.000 147.000 172.500 ;
        RECT 154.500 172.000 233.000 172.500 ;
        RECT 43.500 171.500 81.500 172.000 ;
        RECT 119.000 171.500 147.500 172.000 ;
        RECT 43.000 171.000 81.000 171.500 ;
        RECT 117.500 171.000 148.500 171.500 ;
        RECT 154.000 171.000 233.000 172.000 ;
        RECT 42.000 170.500 80.000 171.000 ;
        RECT 116.000 170.500 149.000 171.000 ;
        RECT 153.500 170.500 233.000 171.000 ;
        RECT 41.500 170.000 79.000 170.500 ;
        RECT 115.000 170.000 149.500 170.500 ;
        RECT 154.000 170.000 233.000 170.500 ;
        RECT 41.000 169.500 78.000 170.000 ;
        RECT 113.500 169.500 150.000 170.000 ;
        RECT 154.500 169.500 232.500 170.000 ;
        RECT 40.500 169.000 77.000 169.500 ;
        RECT 112.000 169.000 151.000 169.500 ;
        RECT 155.500 169.000 232.500 169.500 ;
        RECT 39.500 168.500 76.000 169.000 ;
        RECT 111.000 168.500 151.500 169.000 ;
        RECT 156.000 168.500 232.500 169.000 ;
        RECT 39.000 168.000 75.500 168.500 ;
        RECT 109.500 168.000 152.000 168.500 ;
        RECT 156.500 168.000 232.500 168.500 ;
        RECT 38.500 167.500 74.500 168.000 ;
        RECT 108.500 167.500 152.500 168.000 ;
        RECT 157.000 167.500 232.000 168.000 ;
        RECT 38.000 167.000 73.500 167.500 ;
        RECT 107.500 167.000 153.500 167.500 ;
        RECT 157.500 167.000 232.000 167.500 ;
        RECT 37.500 166.500 73.000 167.000 ;
        RECT 106.000 166.500 154.000 167.000 ;
        RECT 158.000 166.500 232.000 167.000 ;
        RECT 37.000 166.000 72.000 166.500 ;
        RECT 105.000 166.000 154.500 166.500 ;
        RECT 158.500 166.000 232.000 166.500 ;
        RECT 36.000 165.500 71.500 166.000 ;
        RECT 104.000 165.500 155.000 166.000 ;
        RECT 159.000 165.500 231.500 166.000 ;
        RECT 242.000 165.500 242.500 166.000 ;
        RECT 35.500 165.000 70.500 165.500 ;
        RECT 103.000 165.000 155.500 165.500 ;
        RECT 159.500 165.000 231.500 165.500 ;
        RECT 241.500 165.000 242.500 165.500 ;
        RECT 35.000 164.500 70.000 165.000 ;
        RECT 102.000 164.500 156.000 165.000 ;
        RECT 160.000 164.500 231.500 165.000 ;
        RECT 241.000 164.500 242.500 165.000 ;
        RECT 34.500 164.000 69.000 164.500 ;
        RECT 100.500 164.000 156.500 164.500 ;
        RECT 160.500 164.000 231.500 164.500 ;
        RECT 240.000 164.000 242.500 164.500 ;
        RECT 34.000 163.500 68.500 164.000 ;
        RECT 100.000 163.500 157.000 164.000 ;
        RECT 161.000 163.500 231.000 164.000 ;
        RECT 239.500 163.500 242.500 164.000 ;
        RECT 33.500 163.000 67.500 163.500 ;
        RECT 99.000 163.000 157.500 163.500 ;
        RECT 161.500 163.000 231.000 163.500 ;
        RECT 238.500 163.000 242.500 163.500 ;
        RECT 33.000 162.500 67.000 163.000 ;
        RECT 98.000 162.500 158.000 163.000 ;
        RECT 162.000 162.500 230.500 163.000 ;
        RECT 238.000 162.500 242.500 163.000 ;
        RECT 32.500 162.000 66.000 162.500 ;
        RECT 97.000 162.000 158.500 162.500 ;
        RECT 162.000 162.000 228.500 162.500 ;
        RECT 237.000 162.000 242.500 162.500 ;
        RECT 32.000 161.500 65.500 162.000 ;
        RECT 96.000 161.500 159.000 162.000 ;
        RECT 162.500 161.500 226.000 162.000 ;
        RECT 236.000 161.500 242.500 162.000 ;
        RECT 31.500 161.000 65.000 161.500 ;
        RECT 95.000 161.000 159.500 161.500 ;
        RECT 163.000 161.000 223.500 161.500 ;
        RECT 235.000 161.000 242.500 161.500 ;
        RECT 31.000 160.500 64.000 161.000 ;
        RECT 94.000 160.500 160.000 161.000 ;
        RECT 163.500 160.500 221.500 161.000 ;
        RECT 234.000 160.500 242.500 161.000 ;
        RECT 30.500 160.000 63.500 160.500 ;
        RECT 93.000 160.000 160.500 160.500 ;
        RECT 164.000 160.000 219.500 160.500 ;
        RECT 232.500 160.000 242.500 160.500 ;
        RECT 30.000 159.500 63.000 160.000 ;
        RECT 92.500 159.500 161.000 160.000 ;
        RECT 164.500 159.500 218.000 160.000 ;
        RECT 231.000 159.500 242.500 160.000 ;
        RECT 29.500 159.000 62.500 159.500 ;
        RECT 91.500 159.000 161.500 159.500 ;
        RECT 164.500 159.000 216.000 159.500 ;
        RECT 229.000 159.000 242.500 159.500 ;
        RECT 29.500 158.500 61.500 159.000 ;
        RECT 90.500 158.500 162.000 159.000 ;
        RECT 165.000 158.500 214.500 159.000 ;
        RECT 226.500 158.500 243.000 159.000 ;
        RECT 29.000 158.000 61.000 158.500 ;
        RECT 89.500 158.000 162.500 158.500 ;
        RECT 165.500 158.000 213.000 158.500 ;
        RECT 224.000 158.000 243.000 158.500 ;
        RECT 28.500 157.500 60.500 158.000 ;
        RECT 89.000 157.500 162.500 158.000 ;
        RECT 166.000 157.500 211.000 158.000 ;
        RECT 222.000 157.500 243.000 158.000 ;
        RECT 28.000 157.000 60.000 157.500 ;
        RECT 88.000 157.000 163.000 157.500 ;
        RECT 166.500 157.000 209.500 157.500 ;
        RECT 219.500 157.000 243.000 157.500 ;
        RECT 27.500 156.500 59.000 157.000 ;
        RECT 87.500 156.500 163.500 157.000 ;
        RECT 166.500 156.500 208.000 157.000 ;
        RECT 217.500 156.500 243.000 157.000 ;
        RECT 27.000 156.000 58.500 156.500 ;
        RECT 86.500 156.000 164.000 156.500 ;
        RECT 167.000 156.000 207.000 156.500 ;
        RECT 215.500 156.000 243.000 156.500 ;
        RECT 27.000 155.500 58.000 156.000 ;
        RECT 85.500 155.500 164.500 156.000 ;
        RECT 167.500 155.500 205.500 156.000 ;
        RECT 214.000 155.500 243.000 156.000 ;
        RECT 26.500 155.000 57.500 155.500 ;
        RECT 85.000 155.000 165.000 155.500 ;
        RECT 26.000 154.500 57.000 155.000 ;
        RECT 84.000 154.500 165.000 155.000 ;
        RECT 168.000 155.000 204.500 155.500 ;
        RECT 212.000 155.000 243.000 155.500 ;
        RECT 168.000 154.500 203.500 155.000 ;
        RECT 210.500 154.500 243.000 155.000 ;
        RECT 25.500 154.000 56.500 154.500 ;
        RECT 83.500 154.000 165.500 154.500 ;
        RECT 168.500 154.000 202.000 154.500 ;
        RECT 209.000 154.000 243.000 154.500 ;
        RECT 25.000 153.500 56.000 154.000 ;
        RECT 82.500 153.500 166.000 154.000 ;
        RECT 169.000 153.500 201.000 154.000 ;
        RECT 207.500 153.500 243.000 154.000 ;
        RECT 25.000 153.000 55.000 153.500 ;
        RECT 82.000 153.000 166.500 153.500 ;
        RECT 169.000 153.000 200.000 153.500 ;
        RECT 206.000 153.000 243.000 153.500 ;
        RECT 24.500 152.500 54.500 153.000 ;
        RECT 81.000 152.500 166.500 153.000 ;
        RECT 169.500 152.500 199.000 153.000 ;
        RECT 205.000 152.500 243.000 153.000 ;
        RECT 24.000 152.000 54.000 152.500 ;
        RECT 80.500 152.000 167.000 152.500 ;
        RECT 170.000 152.000 198.000 152.500 ;
        RECT 203.500 152.000 243.000 152.500 ;
        RECT 23.500 151.500 53.500 152.000 ;
        RECT 80.000 151.500 167.500 152.000 ;
        RECT 170.000 151.500 197.000 152.000 ;
        RECT 202.500 151.500 243.000 152.000 ;
        RECT 23.500 151.000 53.000 151.500 ;
        RECT 79.000 151.000 168.000 151.500 ;
        RECT 170.500 151.000 196.500 151.500 ;
        RECT 201.500 151.000 243.000 151.500 ;
        RECT 23.000 150.500 52.500 151.000 ;
        RECT 78.500 150.500 168.000 151.000 ;
        RECT 171.000 150.500 195.500 151.000 ;
        RECT 200.500 150.500 243.000 151.000 ;
        RECT 22.500 150.000 52.000 150.500 ;
        RECT 78.000 150.000 168.500 150.500 ;
        RECT 171.000 150.000 194.500 150.500 ;
        RECT 199.500 150.000 242.500 150.500 ;
        RECT 22.500 149.500 51.500 150.000 ;
        RECT 77.000 149.500 169.000 150.000 ;
        RECT 171.500 149.500 194.000 150.000 ;
        RECT 198.500 149.500 242.500 150.000 ;
        RECT 22.000 149.000 51.000 149.500 ;
        RECT 76.500 149.000 169.000 149.500 ;
        RECT 172.000 149.000 193.000 149.500 ;
        RECT 197.500 149.000 242.500 149.500 ;
        RECT 21.500 148.500 50.500 149.000 ;
        RECT 76.000 148.500 169.500 149.000 ;
        RECT 172.000 148.500 192.500 149.000 ;
        RECT 196.500 148.500 242.500 149.000 ;
        RECT 21.500 148.000 50.000 148.500 ;
        RECT 75.000 148.000 170.000 148.500 ;
        RECT 172.500 148.000 191.500 148.500 ;
        RECT 195.500 148.000 242.500 148.500 ;
        RECT 21.000 147.500 49.500 148.000 ;
        RECT 74.500 147.500 170.000 148.000 ;
        RECT 173.000 147.500 191.000 148.000 ;
        RECT 195.000 147.500 242.500 148.000 ;
        RECT 20.500 147.000 49.000 147.500 ;
        RECT 74.000 147.000 170.500 147.500 ;
        RECT 173.000 147.000 190.500 147.500 ;
        RECT 194.000 147.000 242.500 147.500 ;
        RECT 20.500 146.500 48.500 147.000 ;
        RECT 73.500 146.500 171.000 147.000 ;
        RECT 20.000 146.000 48.000 146.500 ;
        RECT 72.500 146.000 171.000 146.500 ;
        RECT 173.500 146.500 189.500 147.000 ;
        RECT 193.500 146.500 242.500 147.000 ;
        RECT 173.500 146.000 189.000 146.500 ;
        RECT 192.500 146.000 242.500 146.500 ;
        RECT 19.500 145.000 47.500 146.000 ;
        RECT 72.000 145.500 171.500 146.000 ;
        RECT 174.000 145.500 188.500 146.000 ;
        RECT 192.000 145.500 242.500 146.000 ;
        RECT 71.500 145.000 171.500 145.500 ;
        RECT 174.500 145.000 188.000 145.500 ;
        RECT 191.000 145.000 242.500 145.500 ;
        RECT 19.000 144.500 47.000 145.000 ;
        RECT 71.000 144.500 172.000 145.000 ;
        RECT 174.500 144.500 187.000 145.000 ;
        RECT 190.500 144.500 242.500 145.000 ;
        RECT 19.000 144.000 46.500 144.500 ;
        RECT 70.500 144.000 172.500 144.500 ;
        RECT 18.500 143.500 46.000 144.000 ;
        RECT 70.000 143.500 172.500 144.000 ;
        RECT 175.000 144.000 186.500 144.500 ;
        RECT 190.000 144.000 242.500 144.500 ;
        RECT 175.000 143.500 186.000 144.000 ;
        RECT 189.000 143.500 242.500 144.000 ;
        RECT 18.500 143.000 45.500 143.500 ;
        RECT 69.000 143.000 173.000 143.500 ;
        RECT 175.500 143.000 185.500 143.500 ;
        RECT 188.500 143.000 242.500 143.500 ;
        RECT 18.000 142.500 45.000 143.000 ;
        RECT 68.500 142.500 173.000 143.000 ;
        RECT 176.000 142.500 185.000 143.000 ;
        RECT 188.000 142.500 242.500 143.000 ;
        RECT 17.500 142.000 44.500 142.500 ;
        RECT 68.000 142.000 173.500 142.500 ;
        RECT 176.000 142.000 184.500 142.500 ;
        RECT 187.500 142.000 242.500 142.500 ;
        RECT 17.500 141.500 44.000 142.000 ;
        RECT 67.500 141.500 148.000 142.000 ;
        RECT 162.000 141.500 173.500 142.000 ;
        RECT 176.500 141.500 184.000 142.000 ;
        RECT 186.500 141.500 242.500 142.000 ;
        RECT 17.000 140.500 43.500 141.500 ;
        RECT 67.000 141.000 145.000 141.500 ;
        RECT 165.000 141.000 174.000 141.500 ;
        RECT 176.500 141.000 183.500 141.500 ;
        RECT 186.000 141.000 242.500 141.500 ;
        RECT 66.500 140.500 87.500 141.000 ;
        RECT 89.000 140.500 142.500 141.000 ;
        RECT 167.500 140.500 174.000 141.000 ;
        RECT 177.000 140.500 183.000 141.000 ;
        RECT 185.500 140.500 242.500 141.000 ;
        RECT 16.500 140.000 43.000 140.500 ;
        RECT 66.000 140.000 87.500 140.500 ;
        RECT 89.500 140.000 140.500 140.500 ;
        RECT 169.500 140.000 174.500 140.500 ;
        RECT 177.000 140.000 182.500 140.500 ;
        RECT 185.000 140.000 242.000 140.500 ;
        RECT 16.500 139.500 42.500 140.000 ;
        RECT 65.500 139.500 87.000 140.000 ;
        RECT 89.500 139.500 139.000 140.000 ;
        RECT 148.000 139.500 162.000 140.000 ;
        RECT 171.000 139.500 174.500 140.000 ;
        RECT 177.500 139.500 182.000 140.000 ;
        RECT 184.500 139.500 242.000 140.000 ;
        RECT 16.000 139.000 42.000 139.500 ;
        RECT 65.000 139.000 87.000 139.500 ;
        RECT 90.000 139.000 137.500 139.500 ;
        RECT 145.000 139.000 165.000 139.500 ;
        RECT 172.500 139.000 175.000 139.500 ;
        RECT 177.500 139.000 181.500 139.500 ;
        RECT 184.000 139.000 242.000 139.500 ;
        RECT 16.000 138.500 41.500 139.000 ;
        RECT 64.000 138.500 86.500 139.000 ;
        RECT 15.500 138.000 41.500 138.500 ;
        RECT 63.500 138.000 86.500 138.500 ;
        RECT 90.500 138.500 136.000 139.000 ;
        RECT 143.000 138.500 167.500 139.000 ;
        RECT 174.000 138.500 175.000 139.000 ;
        RECT 178.000 138.500 181.000 139.000 ;
        RECT 183.500 138.500 242.000 139.000 ;
        RECT 90.500 138.000 135.000 138.500 ;
        RECT 141.000 138.000 169.500 138.500 ;
        RECT 178.000 138.000 180.500 138.500 ;
        RECT 183.000 138.000 242.000 138.500 ;
        RECT 15.500 137.500 41.000 138.000 ;
        RECT 63.000 137.500 86.000 138.000 ;
        RECT 15.500 137.000 40.500 137.500 ;
        RECT 62.500 137.000 86.000 137.500 ;
        RECT 91.000 137.500 133.500 138.000 ;
        RECT 139.000 137.500 171.000 138.000 ;
        RECT 178.500 137.500 180.000 138.000 ;
        RECT 182.500 137.500 242.000 138.000 ;
        RECT 91.000 137.000 132.500 137.500 ;
        RECT 138.000 137.000 172.500 137.500 ;
        RECT 178.500 137.000 179.500 137.500 ;
        RECT 182.000 137.000 242.000 137.500 ;
        RECT 15.000 136.500 40.000 137.000 ;
        RECT 62.000 136.500 86.000 137.000 ;
        RECT 91.500 136.500 131.500 137.000 ;
        RECT 136.500 136.500 173.500 137.000 ;
        RECT 181.500 136.500 242.000 137.000 ;
        RECT 15.000 136.000 39.500 136.500 ;
        RECT 61.500 136.000 85.500 136.500 ;
        RECT 14.500 135.500 39.500 136.000 ;
        RECT 61.000 135.500 85.500 136.000 ;
        RECT 92.000 136.000 130.500 136.500 ;
        RECT 135.000 136.000 175.000 136.500 ;
        RECT 92.000 135.500 129.500 136.000 ;
        RECT 134.000 135.500 176.000 136.000 ;
        RECT 181.000 135.500 242.000 136.500 ;
        RECT 14.500 135.000 39.000 135.500 ;
        RECT 60.500 135.000 85.000 135.500 ;
        RECT 14.000 134.500 38.500 135.000 ;
        RECT 60.000 134.500 85.000 135.000 ;
        RECT 92.500 135.000 128.500 135.500 ;
        RECT 133.000 135.000 177.000 135.500 ;
        RECT 181.500 135.000 241.500 135.500 ;
        RECT 92.500 134.500 127.500 135.000 ;
        RECT 132.000 134.500 178.000 135.000 ;
        RECT 182.500 134.500 241.500 135.000 ;
        RECT 14.000 134.000 38.000 134.500 ;
        RECT 59.500 134.000 85.000 134.500 ;
        RECT 93.000 134.000 127.000 134.500 ;
        RECT 131.000 134.000 179.000 134.500 ;
        RECT 183.500 134.000 241.500 134.500 ;
        RECT 13.500 133.500 38.000 134.000 ;
        RECT 13.500 133.000 37.500 133.500 ;
        RECT 59.000 133.000 84.500 134.000 ;
        RECT 93.000 133.500 126.000 134.000 ;
        RECT 130.000 133.500 180.000 134.000 ;
        RECT 184.000 133.500 241.500 134.000 ;
        RECT 13.500 132.500 37.000 133.000 ;
        RECT 58.500 132.500 84.500 133.000 ;
        RECT 93.500 133.000 125.500 133.500 ;
        RECT 129.000 133.000 181.000 133.500 ;
        RECT 185.000 133.000 241.500 133.500 ;
        RECT 93.500 132.500 124.500 133.000 ;
        RECT 128.500 132.500 181.500 133.000 ;
        RECT 185.500 132.500 241.500 133.000 ;
        RECT 13.000 131.500 36.500 132.500 ;
        RECT 58.000 132.000 84.000 132.500 ;
        RECT 94.000 132.000 124.000 132.500 ;
        RECT 127.500 132.000 182.500 132.500 ;
        RECT 186.500 132.000 241.500 132.500 ;
        RECT 57.500 131.500 84.000 132.000 ;
        RECT 94.500 131.500 123.000 132.000 ;
        RECT 127.000 131.500 183.500 132.000 ;
        RECT 187.000 131.500 241.500 132.000 ;
        RECT 12.500 131.000 36.000 131.500 ;
        RECT 57.000 131.000 83.500 131.500 ;
        RECT 95.000 131.000 122.500 131.500 ;
        RECT 126.000 131.000 184.000 131.500 ;
        RECT 187.500 131.000 241.000 131.500 ;
        RECT 12.500 130.500 35.500 131.000 ;
        RECT 56.500 130.500 83.500 131.000 ;
        RECT 96.000 130.500 122.000 131.000 ;
        RECT 125.500 130.500 185.000 131.000 ;
        RECT 188.500 130.500 241.000 131.000 ;
        RECT 12.500 130.000 35.000 130.500 ;
        RECT 56.000 130.000 83.000 130.500 ;
        RECT 97.000 130.000 121.500 130.500 ;
        RECT 124.500 130.000 185.500 130.500 ;
        RECT 189.000 130.000 241.000 130.500 ;
        RECT 12.000 129.500 35.000 130.000 ;
        RECT 55.500 129.500 82.000 130.000 ;
        RECT 98.500 129.500 120.500 130.000 ;
        RECT 124.000 129.500 186.000 130.000 ;
        RECT 189.500 129.500 241.000 130.000 ;
        RECT 12.000 129.000 34.500 129.500 ;
        RECT 55.000 129.000 81.000 129.500 ;
        RECT 100.000 129.000 120.000 129.500 ;
        RECT 123.500 129.000 187.000 129.500 ;
        RECT 190.000 129.000 241.000 129.500 ;
        RECT 12.000 128.500 34.000 129.000 ;
        RECT 11.500 128.000 34.000 128.500 ;
        RECT 54.500 128.500 80.500 129.000 ;
        RECT 101.000 128.500 119.500 129.000 ;
        RECT 122.500 128.500 187.500 129.000 ;
        RECT 190.500 128.500 241.000 129.000 ;
        RECT 54.500 128.000 79.500 128.500 ;
        RECT 102.500 128.000 119.000 128.500 ;
        RECT 122.000 128.000 188.000 128.500 ;
        RECT 191.500 128.000 241.000 128.500 ;
        RECT 11.500 127.500 33.500 128.000 ;
        RECT 54.000 127.500 78.500 128.000 ;
        RECT 103.500 127.500 118.500 128.000 ;
        RECT 121.500 127.500 188.500 128.000 ;
        RECT 192.000 127.500 240.500 128.000 ;
        RECT 11.500 127.000 33.000 127.500 ;
        RECT 53.500 127.000 77.500 127.500 ;
        RECT 104.500 127.000 118.000 127.500 ;
        RECT 121.000 127.000 189.000 127.500 ;
        RECT 192.500 127.000 240.500 127.500 ;
        RECT 11.000 126.500 33.000 127.000 ;
        RECT 53.000 126.500 76.500 127.000 ;
        RECT 105.000 126.500 117.500 127.000 ;
        RECT 120.500 126.500 189.500 127.000 ;
        RECT 193.000 126.500 240.500 127.000 ;
        RECT 11.000 126.000 32.500 126.500 ;
        RECT 52.500 126.000 76.000 126.500 ;
        RECT 105.000 126.000 117.000 126.500 ;
        RECT 120.000 126.000 190.000 126.500 ;
        RECT 193.500 126.000 240.500 126.500 ;
        RECT 11.000 125.500 32.000 126.000 ;
        RECT 10.500 125.000 32.000 125.500 ;
        RECT 52.000 125.500 75.000 126.000 ;
        RECT 105.000 125.500 116.500 126.000 ;
        RECT 119.500 125.500 190.500 126.000 ;
        RECT 194.000 125.500 240.500 126.000 ;
        RECT 52.000 125.000 74.500 125.500 ;
        RECT 104.000 125.000 116.000 125.500 ;
        RECT 119.000 125.000 191.500 125.500 ;
        RECT 194.500 125.000 240.000 125.500 ;
        RECT 10.500 124.500 31.500 125.000 ;
        RECT 51.500 124.500 74.000 125.000 ;
        RECT 103.500 124.500 115.500 125.000 ;
        RECT 118.500 124.500 192.000 125.000 ;
        RECT 10.500 123.500 31.000 124.500 ;
        RECT 51.000 124.000 73.500 124.500 ;
        RECT 102.500 124.000 115.000 124.500 ;
        RECT 118.000 124.000 192.000 124.500 ;
        RECT 195.000 124.000 240.000 125.000 ;
        RECT 50.500 123.500 73.500 124.000 ;
        RECT 102.000 123.500 114.500 124.000 ;
        RECT 117.500 123.500 192.500 124.000 ;
        RECT 195.500 123.500 240.000 124.000 ;
        RECT 10.000 122.500 30.500 123.500 ;
        RECT 50.000 123.000 74.500 123.500 ;
        RECT 101.000 123.000 114.000 123.500 ;
        RECT 117.000 123.000 193.000 123.500 ;
        RECT 196.000 123.000 240.000 123.500 ;
        RECT 50.000 122.500 75.500 123.000 ;
        RECT 100.000 122.500 113.500 123.000 ;
        RECT 116.500 122.500 193.500 123.000 ;
        RECT 196.500 122.500 239.500 123.000 ;
        RECT 10.000 122.000 30.000 122.500 ;
        RECT 49.500 122.000 76.500 122.500 ;
        RECT 99.000 122.000 113.500 122.500 ;
        RECT 116.000 122.000 194.000 122.500 ;
        RECT 197.000 122.000 239.500 122.500 ;
        RECT 10.000 121.500 29.500 122.000 ;
        RECT 49.000 121.500 78.000 122.000 ;
        RECT 98.000 121.500 113.000 122.000 ;
        RECT 115.500 121.500 194.500 122.000 ;
        RECT 9.500 121.000 29.500 121.500 ;
        RECT 48.500 121.000 79.000 121.500 ;
        RECT 97.500 121.000 112.500 121.500 ;
        RECT 115.000 121.000 195.000 121.500 ;
        RECT 197.500 121.000 239.500 122.000 ;
        RECT 9.500 120.500 29.000 121.000 ;
        RECT 48.000 120.500 80.500 121.000 ;
        RECT 96.500 120.500 112.000 121.000 ;
        RECT 115.000 120.500 195.500 121.000 ;
        RECT 198.000 120.500 239.500 121.000 ;
        RECT 9.500 119.500 28.500 120.500 ;
        RECT 48.000 120.000 82.000 120.500 ;
        RECT 47.500 119.500 83.000 120.000 ;
        RECT 95.500 119.500 111.500 120.500 ;
        RECT 114.500 120.000 195.500 120.500 ;
        RECT 198.500 120.000 239.000 120.500 ;
        RECT 114.000 119.500 196.000 120.000 ;
        RECT 9.000 118.500 28.000 119.500 ;
        RECT 47.000 119.000 84.000 119.500 ;
        RECT 95.000 119.000 111.000 119.500 ;
        RECT 113.500 119.000 196.500 119.500 ;
        RECT 199.000 119.000 239.000 120.000 ;
        RECT 46.500 118.500 84.500 119.000 ;
        RECT 95.000 118.500 110.500 119.000 ;
        RECT 113.500 118.500 197.000 119.000 ;
        RECT 199.500 118.500 239.000 119.000 ;
        RECT 9.000 118.000 27.500 118.500 ;
        RECT 46.500 118.000 85.000 118.500 ;
        RECT 9.000 117.000 27.000 118.000 ;
        RECT 46.000 117.500 85.000 118.000 ;
        RECT 94.500 118.000 110.500 118.500 ;
        RECT 113.000 118.000 197.000 118.500 ;
        RECT 94.500 117.500 110.000 118.000 ;
        RECT 112.500 117.500 197.500 118.000 ;
        RECT 200.000 117.500 238.500 118.500 ;
        RECT 8.500 116.000 26.500 117.000 ;
        RECT 45.500 116.500 85.500 117.500 ;
        RECT 94.000 116.500 109.500 117.500 ;
        RECT 112.500 117.000 198.000 117.500 ;
        RECT 200.500 117.000 238.500 117.500 ;
        RECT 112.000 116.500 198.000 117.000 ;
        RECT 201.000 116.500 238.500 117.000 ;
        RECT 45.000 116.000 86.000 116.500 ;
        RECT 94.000 116.000 109.000 116.500 ;
        RECT 8.500 115.000 26.000 116.000 ;
        RECT 44.500 115.500 86.000 116.000 ;
        RECT 93.500 115.500 109.000 116.000 ;
        RECT 111.500 116.000 198.500 116.500 ;
        RECT 201.000 116.000 238.000 116.500 ;
        RECT 111.500 115.500 199.000 116.000 ;
        RECT 8.500 114.500 25.500 115.000 ;
        RECT 44.000 114.500 86.500 115.500 ;
        RECT 93.500 115.000 108.500 115.500 ;
        RECT 111.000 115.000 199.000 115.500 ;
        RECT 201.500 115.000 238.000 116.000 ;
        RECT 93.500 114.500 108.000 115.000 ;
        RECT 8.000 113.500 25.000 114.500 ;
        RECT 43.500 114.000 87.000 114.500 ;
        RECT 93.000 114.000 108.000 114.500 ;
        RECT 110.500 114.000 199.500 115.000 ;
        RECT 202.000 114.000 237.500 115.000 ;
        RECT 8.000 112.500 24.500 113.500 ;
        RECT 43.000 113.000 87.500 114.000 ;
        RECT 93.000 113.500 107.500 114.000 ;
        RECT 92.500 113.000 107.500 113.500 ;
        RECT 110.000 113.000 200.000 114.000 ;
        RECT 202.500 113.500 237.500 114.000 ;
        RECT 203.000 113.000 237.500 113.500 ;
        RECT 42.500 112.500 88.000 113.000 ;
        RECT 8.000 111.500 24.000 112.500 ;
        RECT 42.000 112.000 88.000 112.500 ;
        RECT 92.500 112.000 107.000 113.000 ;
        RECT 109.500 112.000 200.500 113.000 ;
        RECT 203.000 112.500 237.000 113.000 ;
        RECT 42.000 111.500 88.500 112.000 ;
        RECT 8.000 110.500 23.500 111.500 ;
        RECT 41.500 111.000 89.000 111.500 ;
        RECT 92.000 111.000 106.500 112.000 ;
        RECT 109.000 111.000 201.000 112.000 ;
        RECT 203.500 111.500 237.000 112.500 ;
        RECT 203.500 111.000 236.500 111.500 ;
        RECT 41.000 110.500 62.000 111.000 ;
        RECT 63.000 110.500 89.000 111.000 ;
        RECT 7.500 110.000 23.000 110.500 ;
        RECT 41.000 110.000 61.500 110.500 ;
        RECT 63.000 110.000 89.500 110.500 ;
        RECT 91.500 110.000 106.000 111.000 ;
        RECT 108.500 110.000 201.500 111.000 ;
        RECT 204.000 110.000 236.500 111.000 ;
        RECT 7.500 109.000 22.500 110.000 ;
        RECT 40.500 109.500 61.500 110.000 ;
        RECT 63.500 109.500 90.000 110.000 ;
        RECT 91.000 109.500 106.000 110.000 ;
        RECT 40.500 109.000 61.000 109.500 ;
        RECT 63.500 109.000 105.500 109.500 ;
        RECT 108.000 109.000 202.000 110.000 ;
        RECT 204.500 109.000 236.000 110.000 ;
        RECT 7.500 108.000 22.000 109.000 ;
        RECT 40.000 108.500 61.000 109.000 ;
        RECT 64.000 108.500 105.500 109.000 ;
        RECT 7.500 107.000 21.500 108.000 ;
        RECT 39.500 107.500 60.500 108.500 ;
        RECT 64.000 108.000 105.000 108.500 ;
        RECT 39.000 107.000 60.000 107.500 ;
        RECT 64.500 107.000 105.000 108.000 ;
        RECT 107.500 108.000 202.500 109.000 ;
        RECT 205.000 108.500 236.000 109.000 ;
        RECT 107.500 107.500 203.000 108.000 ;
        RECT 205.000 107.500 235.500 108.500 ;
        RECT 7.500 106.000 21.000 107.000 ;
        RECT 38.500 106.500 60.000 107.000 ;
        RECT 38.500 106.000 59.500 106.500 ;
        RECT 65.000 106.000 104.500 107.000 ;
        RECT 107.000 106.500 203.000 107.500 ;
        RECT 205.500 106.500 235.000 107.500 ;
        RECT 7.500 105.000 20.500 106.000 ;
        RECT 38.000 105.500 59.500 106.000 ;
        RECT 38.000 105.000 59.000 105.500 ;
        RECT 65.500 105.000 104.000 106.000 ;
        RECT 106.500 105.000 203.500 106.500 ;
        RECT 206.000 106.000 235.000 106.500 ;
        RECT 206.000 105.000 234.500 106.000 ;
        RECT 7.000 104.000 20.000 105.000 ;
        RECT 37.500 104.500 59.000 105.000 ;
        RECT 66.000 104.500 104.000 105.000 ;
        RECT 37.000 104.000 58.500 104.500 ;
        RECT 66.000 104.000 103.500 104.500 ;
        RECT 7.000 103.000 19.500 104.000 ;
        RECT 37.000 103.500 58.000 104.000 ;
        RECT 66.500 103.500 103.500 104.000 ;
        RECT 36.500 103.000 57.500 103.500 ;
        RECT 67.000 103.000 103.500 103.500 ;
        RECT 106.000 103.500 204.000 105.000 ;
        RECT 206.500 103.500 234.000 105.000 ;
        RECT 106.000 103.000 204.500 103.500 ;
        RECT 206.500 103.000 233.500 103.500 ;
        RECT 7.000 102.000 19.000 103.000 ;
        RECT 36.500 102.500 56.000 103.000 ;
        RECT 68.000 102.500 103.500 103.000 ;
        RECT 36.000 102.000 55.000 102.500 ;
        RECT 69.500 102.000 103.000 102.500 ;
        RECT 7.000 101.000 18.500 102.000 ;
        RECT 36.000 101.500 54.000 102.000 ;
        RECT 70.500 101.500 103.000 102.000 ;
        RECT 105.500 101.500 204.500 103.000 ;
        RECT 207.000 102.500 233.500 103.000 ;
        RECT 207.000 101.500 233.000 102.500 ;
        RECT 35.500 101.000 53.000 101.500 ;
        RECT 71.500 101.000 103.000 101.500 ;
        RECT 7.000 100.000 18.000 101.000 ;
        RECT 35.000 100.500 52.000 101.000 ;
        RECT 72.500 100.500 103.000 101.000 ;
        RECT 35.000 100.000 51.500 100.500 ;
        RECT 73.000 100.000 102.500 100.500 ;
        RECT 7.000 98.500 17.500 100.000 ;
        RECT 34.500 99.000 51.500 100.000 ;
        RECT 73.500 99.000 102.500 100.000 ;
        RECT 105.000 99.500 205.000 101.500 ;
        RECT 207.000 101.000 232.500 101.500 ;
        RECT 207.500 100.500 232.500 101.000 ;
        RECT 207.500 99.500 232.000 100.500 ;
        RECT 105.000 99.000 205.500 99.500 ;
        RECT 207.500 99.000 231.500 99.500 ;
        RECT 34.000 98.500 52.000 99.000 ;
        RECT 72.500 98.500 102.500 99.000 ;
        RECT 7.000 97.500 17.000 98.500 ;
        RECT 34.000 98.000 53.000 98.500 ;
        RECT 71.500 98.000 102.500 98.500 ;
        RECT 33.500 97.500 54.000 98.000 ;
        RECT 70.500 97.500 102.000 98.000 ;
        RECT 7.000 96.500 16.500 97.500 ;
        RECT 33.500 97.000 55.000 97.500 ;
        RECT 69.500 97.000 102.000 97.500 ;
        RECT 33.000 96.500 56.000 97.000 ;
        RECT 68.500 96.500 102.000 97.000 ;
        RECT 104.500 97.000 205.500 99.000 ;
        RECT 208.000 98.500 231.500 99.000 ;
        RECT 208.000 97.500 231.000 98.500 ;
        RECT 104.500 96.500 206.000 97.000 ;
        RECT 7.000 96.000 16.000 96.500 ;
        RECT 33.000 96.000 57.500 96.500 ;
        RECT 67.500 96.000 102.000 96.500 ;
        RECT 7.500 95.500 16.000 96.000 ;
        RECT 32.500 95.500 58.000 96.000 ;
        RECT 66.500 95.500 102.000 96.000 ;
        RECT 7.500 94.500 15.500 95.500 ;
        RECT 32.000 95.000 58.500 95.500 ;
        RECT 32.000 94.500 59.000 95.000 ;
        RECT 66.000 94.500 102.000 95.500 ;
        RECT 7.500 93.000 15.000 94.500 ;
        RECT 31.500 93.500 59.000 94.500 ;
        RECT 65.500 93.500 101.500 94.500 ;
        RECT 7.500 92.000 14.500 93.000 ;
        RECT 31.000 92.500 59.500 93.500 ;
        RECT 65.000 92.500 101.500 93.500 ;
        RECT 7.500 91.000 14.000 92.000 ;
        RECT 30.500 91.500 60.000 92.500 ;
        RECT 64.500 91.500 101.500 92.500 ;
        RECT 7.500 90.000 13.500 91.000 ;
        RECT 30.000 90.500 60.500 91.500 ;
        RECT 64.000 90.500 101.500 91.500 ;
        RECT 8.000 89.500 13.500 90.000 ;
        RECT 29.500 89.500 61.000 90.500 ;
        RECT 63.500 89.500 101.500 90.500 ;
        RECT 104.000 92.000 206.000 96.500 ;
        RECT 208.000 96.500 230.500 97.500 ;
        RECT 208.000 96.000 230.000 96.500 ;
        RECT 208.500 95.000 229.500 96.000 ;
        RECT 208.500 94.000 229.000 95.000 ;
        RECT 208.500 93.500 228.500 94.000 ;
        RECT 208.500 92.500 228.000 93.500 ;
        RECT 104.000 90.000 206.500 92.000 ;
        RECT 8.000 88.500 13.000 89.500 ;
        RECT 29.500 89.000 61.500 89.500 ;
        RECT 63.000 89.000 101.500 89.500 ;
        RECT 29.000 88.500 61.500 89.000 ;
        RECT 62.500 88.500 101.500 89.000 ;
        RECT 8.000 87.500 12.500 88.500 ;
        RECT 29.000 88.000 101.500 88.500 ;
        RECT 8.000 86.500 12.000 87.500 ;
        RECT 28.500 87.000 101.500 88.000 ;
        RECT 103.500 87.500 206.500 90.000 ;
        RECT 208.500 91.500 227.500 92.500 ;
        RECT 208.500 91.000 227.000 91.500 ;
        RECT 208.500 90.500 226.500 91.000 ;
        RECT 208.500 89.500 226.000 90.500 ;
        RECT 209.000 89.000 225.500 89.500 ;
        RECT 209.000 88.000 225.000 89.000 ;
        RECT 209.000 87.500 224.500 88.000 ;
        RECT 234.000 87.500 235.500 88.000 ;
        RECT 8.500 86.000 12.000 86.500 ;
        RECT 28.000 86.000 101.500 87.000 ;
        RECT 8.500 85.000 11.500 86.000 ;
        RECT 27.500 85.000 101.500 86.000 ;
        RECT 8.500 83.500 11.000 85.000 ;
        RECT 27.000 84.500 101.500 85.000 ;
        RECT 27.000 84.000 87.500 84.500 ;
        RECT 88.500 84.000 101.500 84.500 ;
        RECT 9.000 82.500 10.500 83.500 ;
        RECT 26.500 82.500 87.000 84.000 ;
        RECT 89.000 83.000 101.500 84.000 ;
        RECT 89.500 82.500 101.500 83.000 ;
        RECT 104.000 86.500 206.500 87.500 ;
        RECT 208.500 87.000 224.000 87.500 ;
        RECT 232.500 87.000 235.500 87.500 ;
        RECT 208.500 86.500 216.500 87.000 ;
        RECT 231.000 86.500 235.000 87.000 ;
        RECT 104.000 86.000 206.000 86.500 ;
        RECT 229.000 86.000 235.000 86.500 ;
        RECT 104.000 85.500 189.000 86.000 ;
        RECT 227.500 85.500 235.000 86.000 ;
        RECT 104.000 85.000 183.500 85.500 ;
        RECT 225.500 85.000 234.500 85.500 ;
        RECT 104.000 84.500 180.500 85.000 ;
        RECT 223.000 84.500 234.500 85.000 ;
        RECT 104.000 84.000 178.000 84.500 ;
        RECT 217.000 84.000 234.500 84.500 ;
        RECT 104.000 83.500 176.000 84.000 ;
        RECT 209.000 83.500 234.000 84.000 ;
        RECT 104.000 83.000 174.500 83.500 ;
        RECT 191.000 83.000 234.000 83.500 ;
        RECT 104.000 82.500 172.500 83.000 ;
        RECT 185.000 82.500 233.500 83.000 ;
        RECT 9.000 81.000 10.000 82.500 ;
        RECT 26.000 81.500 86.500 82.500 ;
        RECT 89.500 82.000 102.000 82.500 ;
        RECT 25.500 80.500 86.000 81.500 ;
        RECT 90.000 81.000 102.000 82.000 ;
        RECT 104.000 82.000 171.000 82.500 ;
        RECT 182.000 82.000 233.500 82.500 ;
        RECT 104.000 81.500 169.500 82.000 ;
        RECT 179.500 81.500 233.500 82.000 ;
        RECT 90.500 80.500 102.000 81.000 ;
        RECT 25.000 80.000 85.500 80.500 ;
        RECT 91.500 80.000 102.000 80.500 ;
        RECT 25.000 79.500 84.500 80.000 ;
        RECT 92.500 79.500 102.000 80.000 ;
        RECT 25.000 79.000 83.500 79.500 ;
        RECT 93.500 79.000 102.000 79.500 ;
        RECT 104.500 81.000 168.500 81.500 ;
        RECT 177.500 81.000 233.000 81.500 ;
        RECT 104.500 80.500 167.000 81.000 ;
        RECT 175.500 80.500 233.000 81.000 ;
        RECT 104.500 80.000 166.000 80.500 ;
        RECT 174.000 80.000 232.500 80.500 ;
        RECT 104.500 79.500 165.000 80.000 ;
        RECT 172.000 79.500 232.500 80.000 ;
        RECT 104.500 79.000 163.500 79.500 ;
        RECT 171.000 79.000 232.000 79.500 ;
        RECT 24.500 78.500 82.500 79.000 ;
        RECT 24.500 78.000 81.500 78.500 ;
        RECT 24.000 77.500 81.500 78.000 ;
        RECT 94.500 77.500 102.500 79.000 ;
        RECT 104.500 78.500 162.500 79.000 ;
        RECT 169.500 78.500 232.000 79.000 ;
        RECT 24.000 77.000 82.500 77.500 ;
        RECT 93.500 77.000 102.500 77.500 ;
        RECT 24.000 76.500 83.500 77.000 ;
        RECT 92.500 76.500 102.500 77.000 ;
        RECT 105.000 78.000 161.500 78.500 ;
        RECT 168.000 78.000 231.500 78.500 ;
        RECT 105.000 77.500 160.500 78.000 ;
        RECT 166.500 77.500 231.500 78.000 ;
        RECT 105.000 77.000 159.500 77.500 ;
        RECT 165.500 77.000 231.000 77.500 ;
        RECT 105.000 76.500 158.500 77.000 ;
        RECT 164.000 76.500 231.000 77.000 ;
        RECT 23.500 76.000 84.500 76.500 ;
        RECT 91.500 76.000 103.000 76.500 ;
        RECT 23.500 75.500 85.500 76.000 ;
        RECT 23.000 75.000 86.000 75.500 ;
        RECT 90.500 75.000 103.000 76.000 ;
        RECT 23.000 74.000 86.500 75.000 ;
        RECT 90.000 74.500 103.000 75.000 ;
        RECT 105.500 76.000 157.500 76.500 ;
        RECT 163.000 76.000 230.500 76.500 ;
        RECT 105.500 75.500 157.000 76.000 ;
        RECT 162.000 75.500 230.500 76.000 ;
        RECT 105.500 75.000 156.000 75.500 ;
        RECT 161.000 75.000 230.000 75.500 ;
        RECT 105.500 74.500 155.000 75.000 ;
        RECT 160.000 74.500 230.000 75.000 ;
        RECT 90.000 74.000 103.500 74.500 ;
        RECT 22.500 73.000 59.000 74.000 ;
        RECT 60.500 73.000 87.000 74.000 ;
        RECT 89.500 73.000 103.500 74.000 ;
        RECT 106.000 74.000 154.000 74.500 ;
        RECT 159.000 74.000 229.500 74.500 ;
        RECT 106.000 73.500 153.000 74.000 ;
        RECT 158.000 73.500 229.500 74.000 ;
        RECT 106.000 73.000 152.500 73.500 ;
        RECT 157.000 73.000 229.000 73.500 ;
        RECT 22.000 72.000 58.500 73.000 ;
        RECT 61.000 72.000 87.500 73.000 ;
        RECT 89.500 72.500 104.000 73.000 ;
        RECT 22.000 71.500 58.000 72.000 ;
        RECT 21.500 71.000 58.000 71.500 ;
        RECT 61.500 71.500 88.000 72.000 ;
        RECT 89.000 71.500 104.000 72.500 ;
        RECT 106.500 72.500 151.500 73.000 ;
        RECT 156.000 72.500 229.000 73.000 ;
        RECT 106.500 72.000 150.500 72.500 ;
        RECT 155.000 72.000 228.500 72.500 ;
        RECT 106.500 71.500 149.500 72.000 ;
        RECT 154.000 71.500 228.000 72.000 ;
        RECT 61.500 71.000 104.500 71.500 ;
        RECT 21.500 70.000 57.500 71.000 ;
        RECT 62.000 70.000 104.500 71.000 ;
        RECT 107.000 71.000 149.000 71.500 ;
        RECT 153.000 71.000 228.000 71.500 ;
        RECT 107.000 70.500 148.000 71.000 ;
        RECT 152.500 70.500 227.500 71.000 ;
        RECT 107.500 70.000 147.000 70.500 ;
        RECT 151.500 70.000 227.500 70.500 ;
        RECT 21.000 69.500 57.000 70.000 ;
        RECT 62.500 69.500 105.000 70.000 ;
        RECT 21.000 69.000 56.000 69.500 ;
        RECT 63.500 69.000 105.000 69.500 ;
        RECT 107.500 69.500 146.500 70.000 ;
        RECT 151.000 69.500 227.000 70.000 ;
        RECT 107.500 69.000 145.500 69.500 ;
        RECT 150.000 69.000 226.500 69.500 ;
        RECT 21.000 68.500 55.000 69.000 ;
        RECT 64.500 68.500 105.000 69.000 ;
        RECT 108.000 68.500 144.500 69.000 ;
        RECT 149.000 68.500 226.500 69.000 ;
        RECT 20.500 68.000 54.000 68.500 ;
        RECT 65.500 68.000 105.500 68.500 ;
        RECT 108.000 68.000 144.000 68.500 ;
        RECT 148.500 68.000 226.000 68.500 ;
        RECT 20.500 67.500 53.000 68.000 ;
        RECT 20.000 66.500 53.000 67.500 ;
        RECT 66.500 67.500 105.500 68.000 ;
        RECT 108.500 67.500 143.000 68.000 ;
        RECT 147.500 67.500 225.500 68.000 ;
        RECT 66.500 66.500 106.000 67.500 ;
        RECT 108.500 67.000 142.500 67.500 ;
        RECT 147.000 67.000 225.500 67.500 ;
        RECT 109.000 66.500 141.500 67.000 ;
        RECT 146.000 66.500 225.000 67.000 ;
        RECT 20.000 66.000 54.000 66.500 ;
        RECT 66.000 66.000 106.500 66.500 ;
        RECT 109.000 66.000 140.500 66.500 ;
        RECT 145.500 66.000 224.500 66.500 ;
        RECT 19.500 65.500 54.500 66.000 ;
        RECT 65.000 65.500 106.500 66.000 ;
        RECT 19.500 65.000 56.000 65.500 ;
        RECT 63.500 65.000 106.500 65.500 ;
        RECT 109.500 65.500 140.000 66.000 ;
        RECT 144.500 65.500 224.000 66.000 ;
        RECT 109.500 65.000 139.000 65.500 ;
        RECT 143.500 65.000 224.000 65.500 ;
        RECT 19.500 64.500 57.000 65.000 ;
        RECT 62.500 64.500 107.000 65.000 ;
        RECT 19.000 63.500 57.500 64.500 ;
        RECT 62.000 64.000 107.000 64.500 ;
        RECT 110.000 64.500 138.500 65.000 ;
        RECT 143.000 64.500 223.500 65.000 ;
        RECT 110.000 64.000 137.500 64.500 ;
        RECT 142.000 64.000 223.000 64.500 ;
        RECT 62.000 63.500 107.500 64.000 ;
        RECT 110.500 63.500 137.000 64.000 ;
        RECT 141.500 63.500 222.500 64.000 ;
        RECT 19.000 63.000 58.000 63.500 ;
        RECT 18.500 62.500 58.000 63.000 ;
        RECT 61.500 62.500 108.000 63.500 ;
        RECT 110.500 63.000 136.000 63.500 ;
        RECT 140.500 63.000 222.500 63.500 ;
        RECT 111.000 62.500 135.500 63.000 ;
        RECT 139.500 62.500 222.000 63.000 ;
        RECT 18.500 61.500 58.500 62.500 ;
        RECT 61.000 61.500 108.500 62.500 ;
        RECT 111.000 62.000 134.500 62.500 ;
        RECT 139.000 62.000 221.500 62.500 ;
        RECT 111.500 61.500 134.000 62.000 ;
        RECT 138.000 61.500 221.000 62.000 ;
        RECT 18.000 60.500 59.000 61.500 ;
        RECT 60.500 60.500 109.000 61.500 ;
        RECT 112.000 61.000 133.000 61.500 ;
        RECT 137.500 61.000 220.500 61.500 ;
        RECT 112.000 60.500 132.500 61.000 ;
        RECT 136.500 60.500 220.000 61.000 ;
        RECT 18.000 60.000 109.500 60.500 ;
        RECT 112.500 60.000 131.500 60.500 ;
        RECT 136.000 60.000 220.000 60.500 ;
        RECT 17.500 59.000 110.000 60.000 ;
        RECT 113.000 59.500 131.000 60.000 ;
        RECT 135.000 59.500 219.500 60.000 ;
        RECT 113.000 59.000 130.000 59.500 ;
        RECT 134.500 59.000 219.000 59.500 ;
        RECT 17.500 58.500 110.500 59.000 ;
        RECT 113.500 58.500 129.500 59.000 ;
        RECT 133.500 58.500 218.500 59.000 ;
        RECT 18.000 57.500 111.000 58.500 ;
        RECT 114.000 58.000 129.000 58.500 ;
        RECT 132.500 58.000 218.000 58.500 ;
        RECT 114.500 57.500 128.000 58.000 ;
        RECT 132.000 57.500 217.500 58.000 ;
        RECT 18.500 56.500 110.500 57.500 ;
        RECT 114.500 57.000 127.500 57.500 ;
        RECT 131.000 57.000 217.000 57.500 ;
        RECT 115.000 56.500 126.500 57.000 ;
        RECT 130.500 56.500 216.500 57.000 ;
        RECT 19.000 56.000 110.000 56.500 ;
        RECT 115.500 56.000 126.000 56.500 ;
        RECT 130.000 56.000 216.000 56.500 ;
        RECT 19.000 55.500 109.500 56.000 ;
        RECT 116.000 55.500 125.000 56.000 ;
        RECT 129.000 55.500 215.500 56.000 ;
        RECT 19.500 55.000 109.000 55.500 ;
        RECT 112.000 55.000 113.000 55.500 ;
        RECT 116.500 55.000 124.500 55.500 ;
        RECT 128.500 55.000 215.000 55.500 ;
        RECT 20.000 54.500 108.500 55.000 ;
        RECT 111.500 54.500 113.500 55.000 ;
        RECT 20.000 54.000 108.000 54.500 ;
        RECT 111.000 54.000 113.500 54.500 ;
        RECT 117.000 54.500 124.000 55.000 ;
        RECT 127.500 54.500 214.500 55.000 ;
        RECT 117.000 54.000 123.000 54.500 ;
        RECT 127.000 54.000 214.000 54.500 ;
        RECT 20.500 53.500 107.500 54.000 ;
        RECT 110.500 53.500 114.000 54.000 ;
        RECT 117.500 53.500 122.500 54.000 ;
        RECT 126.000 53.500 213.500 54.000 ;
        RECT 20.500 53.000 107.000 53.500 ;
        RECT 110.000 53.000 114.500 53.500 ;
        RECT 118.000 53.000 121.500 53.500 ;
        RECT 125.500 53.000 213.000 53.500 ;
        RECT 21.000 52.500 106.500 53.000 ;
        RECT 109.500 52.500 115.000 53.000 ;
        RECT 118.500 52.500 121.000 53.000 ;
        RECT 124.500 52.500 212.500 53.000 ;
        RECT 21.500 52.000 106.500 52.500 ;
        RECT 109.000 52.000 115.500 52.500 ;
        RECT 119.000 52.000 120.000 52.500 ;
        RECT 124.000 52.000 212.000 52.500 ;
        RECT 21.500 51.500 106.000 52.000 ;
        RECT 108.500 51.500 116.000 52.000 ;
        RECT 123.000 51.500 211.500 52.000 ;
        RECT 22.000 51.000 105.500 51.500 ;
        RECT 108.000 51.000 116.500 51.500 ;
        RECT 122.500 51.000 210.500 51.500 ;
        RECT 22.500 50.500 105.000 51.000 ;
        RECT 22.500 50.000 104.500 50.500 ;
        RECT 107.500 50.000 117.000 51.000 ;
        RECT 121.500 50.500 210.000 51.000 ;
        RECT 121.000 50.000 209.500 50.500 ;
        RECT 23.000 49.500 104.000 50.000 ;
        RECT 107.000 49.500 116.500 50.000 ;
        RECT 120.000 49.500 209.000 50.000 ;
        RECT 23.500 49.000 103.500 49.500 ;
        RECT 106.500 49.000 116.000 49.500 ;
        RECT 119.500 49.000 208.500 49.500 ;
        RECT 23.500 48.500 103.000 49.000 ;
        RECT 106.000 48.500 115.000 49.000 ;
        RECT 118.500 48.500 207.500 49.000 ;
        RECT 24.000 48.000 102.500 48.500 ;
        RECT 105.500 48.000 114.500 48.500 ;
        RECT 118.000 48.000 207.000 48.500 ;
        RECT 24.500 47.500 102.000 48.000 ;
        RECT 105.000 47.500 113.500 48.000 ;
        RECT 117.000 47.500 206.500 48.000 ;
        RECT 25.000 47.000 102.000 47.500 ;
        RECT 104.500 47.000 113.000 47.500 ;
        RECT 116.500 47.000 206.000 47.500 ;
        RECT 25.000 46.500 101.500 47.000 ;
        RECT 104.000 46.500 112.000 47.000 ;
        RECT 115.500 46.500 205.000 47.000 ;
        RECT 25.500 46.000 101.000 46.500 ;
        RECT 103.500 46.000 111.500 46.500 ;
        RECT 115.000 46.000 204.500 46.500 ;
        RECT 26.000 45.500 100.500 46.000 ;
        RECT 103.000 45.500 111.000 46.000 ;
        RECT 114.000 45.500 204.000 46.000 ;
        RECT 26.500 45.000 100.000 45.500 ;
        RECT 102.500 45.000 110.000 45.500 ;
        RECT 113.500 45.000 203.000 45.500 ;
        RECT 27.000 44.500 99.500 45.000 ;
        RECT 102.000 44.500 109.000 45.000 ;
        RECT 112.500 44.500 202.500 45.000 ;
        RECT 27.000 44.000 99.000 44.500 ;
        RECT 101.500 44.000 108.500 44.500 ;
        RECT 112.000 44.000 202.000 44.500 ;
        RECT 27.500 43.500 98.500 44.000 ;
        RECT 101.000 43.500 107.500 44.000 ;
        RECT 111.000 43.500 201.000 44.000 ;
        RECT 28.000 43.000 98.000 43.500 ;
        RECT 101.000 43.000 107.000 43.500 ;
        RECT 110.500 43.000 200.500 43.500 ;
        RECT 28.500 42.500 97.500 43.000 ;
        RECT 100.500 42.500 106.000 43.000 ;
        RECT 109.500 42.500 199.500 43.000 ;
        RECT 29.000 42.000 97.000 42.500 ;
        RECT 100.000 42.000 105.500 42.500 ;
        RECT 109.000 42.000 199.000 42.500 ;
        RECT 29.500 41.500 96.500 42.000 ;
        RECT 99.500 41.500 104.500 42.000 ;
        RECT 108.000 41.500 198.000 42.000 ;
        RECT 29.500 41.000 96.000 41.500 ;
        RECT 99.000 41.000 104.000 41.500 ;
        RECT 107.500 41.000 197.500 41.500 ;
        RECT 30.000 40.500 96.000 41.000 ;
        RECT 98.500 40.500 103.000 41.000 ;
        RECT 106.500 40.500 196.500 41.000 ;
        RECT 30.500 40.000 95.500 40.500 ;
        RECT 98.000 40.000 102.500 40.500 ;
        RECT 105.500 40.000 196.000 40.500 ;
        RECT 31.000 39.500 95.000 40.000 ;
        RECT 97.500 39.500 101.500 40.000 ;
        RECT 105.000 39.500 195.000 40.000 ;
        RECT 31.500 39.000 94.500 39.500 ;
        RECT 97.000 39.000 101.000 39.500 ;
        RECT 104.000 39.000 194.500 39.500 ;
        RECT 32.000 38.500 94.000 39.000 ;
        RECT 96.500 38.500 100.000 39.000 ;
        RECT 103.500 38.500 193.500 39.000 ;
        RECT 32.500 38.000 93.500 38.500 ;
        RECT 96.000 38.000 99.000 38.500 ;
        RECT 103.000 38.000 192.500 38.500 ;
        RECT 33.000 37.500 93.000 38.000 ;
        RECT 95.500 37.500 98.500 38.000 ;
        RECT 102.000 37.500 192.000 38.000 ;
        RECT 33.500 37.000 92.500 37.500 ;
        RECT 95.000 37.000 97.500 37.500 ;
        RECT 101.500 37.000 191.000 37.500 ;
        RECT 34.000 36.500 92.000 37.000 ;
        RECT 94.500 36.500 97.000 37.000 ;
        RECT 100.500 36.500 190.000 37.000 ;
        RECT 34.500 36.000 91.500 36.500 ;
        RECT 94.000 36.000 96.000 36.500 ;
        RECT 100.000 36.000 189.000 36.500 ;
        RECT 35.000 35.500 91.000 36.000 ;
        RECT 93.500 35.500 95.000 36.000 ;
        RECT 99.000 35.500 188.500 36.000 ;
        RECT 35.500 35.000 90.500 35.500 ;
        RECT 93.000 35.000 94.500 35.500 ;
        RECT 98.500 35.000 187.500 35.500 ;
        RECT 36.000 34.500 90.000 35.000 ;
        RECT 92.500 34.500 94.000 35.000 ;
        RECT 97.500 34.500 186.500 35.000 ;
        RECT 36.500 34.000 89.500 34.500 ;
        RECT 92.000 34.000 93.500 34.500 ;
        RECT 97.000 34.000 185.500 34.500 ;
        RECT 37.500 33.500 89.000 34.000 ;
        RECT 91.500 33.500 92.500 34.000 ;
        RECT 96.000 33.500 184.500 34.000 ;
        RECT 38.000 33.000 88.500 33.500 ;
        RECT 95.500 33.000 183.500 33.500 ;
        RECT 38.500 32.500 88.000 33.000 ;
        RECT 94.500 32.500 182.500 33.000 ;
        RECT 39.000 32.000 87.500 32.500 ;
        RECT 93.500 32.000 181.500 32.500 ;
        RECT 39.500 31.500 87.000 32.000 ;
        RECT 93.000 31.500 180.500 32.000 ;
        RECT 40.500 31.000 86.500 31.500 ;
        RECT 92.000 31.000 179.500 31.500 ;
        RECT 41.000 30.500 86.000 31.000 ;
        RECT 91.500 30.500 178.500 31.000 ;
        RECT 41.500 30.000 85.500 30.500 ;
        RECT 90.500 30.000 177.500 30.500 ;
        RECT 42.000 29.500 85.000 30.000 ;
        RECT 89.500 29.500 176.500 30.000 ;
        RECT 43.000 29.000 84.000 29.500 ;
        RECT 89.000 29.000 175.500 29.500 ;
        RECT 43.500 28.500 83.500 29.000 ;
        RECT 88.000 28.500 174.000 29.000 ;
        RECT 44.500 28.000 82.500 28.500 ;
        RECT 87.000 28.000 173.000 28.500 ;
        RECT 45.000 27.500 81.500 28.000 ;
        RECT 86.500 27.500 172.000 28.000 ;
        RECT 45.500 27.000 80.500 27.500 ;
        RECT 85.500 27.000 170.500 27.500 ;
        RECT 46.500 26.500 79.500 27.000 ;
        RECT 84.500 26.500 169.500 27.000 ;
        RECT 47.000 26.000 78.500 26.500 ;
        RECT 83.500 26.000 168.500 26.500 ;
        RECT 48.000 25.500 78.000 26.000 ;
        RECT 82.500 25.500 167.000 26.000 ;
        RECT 48.500 25.000 77.000 25.500 ;
        RECT 82.000 25.000 166.000 25.500 ;
        RECT 49.500 24.500 76.000 25.000 ;
        RECT 81.000 24.500 164.500 25.000 ;
        RECT 50.500 24.000 75.000 24.500 ;
        RECT 80.000 24.000 163.000 24.500 ;
        RECT 51.500 23.500 74.000 24.000 ;
        RECT 79.000 23.500 162.000 24.000 ;
        RECT 52.000 23.000 73.000 23.500 ;
        RECT 78.000 23.000 160.500 23.500 ;
        RECT 53.000 22.500 72.500 23.000 ;
        RECT 77.000 22.500 159.000 23.000 ;
        RECT 54.000 22.000 71.500 22.500 ;
        RECT 76.500 22.000 157.500 22.500 ;
        RECT 55.000 21.500 70.500 22.000 ;
        RECT 75.500 21.500 156.500 22.000 ;
        RECT 56.000 21.000 69.500 21.500 ;
        RECT 74.500 21.000 155.000 21.500 ;
        RECT 57.000 20.500 68.500 21.000 ;
        RECT 73.500 20.500 153.500 21.000 ;
        RECT 58.000 20.000 67.500 20.500 ;
        RECT 72.500 20.000 152.000 20.500 ;
        RECT 59.000 19.500 66.500 20.000 ;
        RECT 71.500 19.500 150.000 20.000 ;
        RECT 60.000 19.000 65.500 19.500 ;
        RECT 70.500 19.000 148.500 19.500 ;
        RECT 61.500 18.500 64.500 19.000 ;
        RECT 69.500 18.500 147.000 19.000 ;
        RECT 62.500 18.000 63.500 18.500 ;
        RECT 68.500 18.000 145.000 18.500 ;
        RECT 67.500 17.500 143.500 18.000 ;
        RECT 66.500 17.000 141.500 17.500 ;
        RECT 65.500 16.500 140.000 17.000 ;
        RECT 64.000 16.000 138.000 16.500 ;
        RECT 63.000 15.500 136.000 16.000 ;
        RECT 62.000 15.000 134.000 15.500 ;
        RECT 61.000 14.500 131.500 15.000 ;
        RECT 60.000 14.000 129.000 14.500 ;
        RECT 59.000 13.500 126.500 14.000 ;
        RECT 57.500 13.000 123.500 13.500 ;
        RECT 56.500 12.500 120.000 13.000 ;
        RECT 55.500 12.000 115.000 12.500 ;
        RECT 54.500 11.500 105.000 12.000 ;
        RECT 53.000 11.000 81.500 11.500 ;
        RECT 87.000 11.000 91.000 11.500 ;
        RECT 52.000 10.500 69.500 11.000 ;
        RECT 51.000 10.000 64.500 10.500 ;
        RECT 49.500 9.500 60.500 10.000 ;
        RECT 48.500 9.000 57.000 9.500 ;
        RECT 47.000 8.500 54.000 9.000 ;
        RECT 46.000 8.000 51.500 8.500 ;
        RECT 44.500 7.500 48.500 8.000 ;
        RECT 43.000 7.000 46.000 7.500 ;
        RECT 41.500 6.500 43.500 7.000 ;
        RECT 39.500 6.000 42.000 6.500 ;
        RECT 39.000 5.500 40.000 6.000 ;
  END
END aef2
END LIBRARY

