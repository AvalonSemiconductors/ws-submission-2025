magic
tech gf180mcuD
magscale 1 10
timestamp 1762867098
<< pwell >>
rect -996 -30488 996 30488
<< mvnmos >>
rect -732 10232 -612 30232
rect -508 10232 -388 30232
rect -284 10232 -164 30232
rect -60 10232 60 30232
rect 164 10232 284 30232
rect 388 10232 508 30232
rect 612 10232 732 30232
rect -732 -10000 -612 10000
rect -508 -10000 -388 10000
rect -284 -10000 -164 10000
rect -60 -10000 60 10000
rect 164 -10000 284 10000
rect 388 -10000 508 10000
rect 612 -10000 732 10000
rect -732 -30232 -612 -10232
rect -508 -30232 -388 -10232
rect -284 -30232 -164 -10232
rect -60 -30232 60 -10232
rect 164 -30232 284 -10232
rect 388 -30232 508 -10232
rect 612 -30232 732 -10232
<< mvndiff >>
rect -820 30219 -732 30232
rect -820 10245 -807 30219
rect -761 10245 -732 30219
rect -820 10232 -732 10245
rect -612 30219 -508 30232
rect -612 10245 -583 30219
rect -537 10245 -508 30219
rect -612 10232 -508 10245
rect -388 30219 -284 30232
rect -388 10245 -359 30219
rect -313 10245 -284 30219
rect -388 10232 -284 10245
rect -164 30219 -60 30232
rect -164 10245 -135 30219
rect -89 10245 -60 30219
rect -164 10232 -60 10245
rect 60 30219 164 30232
rect 60 10245 89 30219
rect 135 10245 164 30219
rect 60 10232 164 10245
rect 284 30219 388 30232
rect 284 10245 313 30219
rect 359 10245 388 30219
rect 284 10232 388 10245
rect 508 30219 612 30232
rect 508 10245 537 30219
rect 583 10245 612 30219
rect 508 10232 612 10245
rect 732 30219 820 30232
rect 732 10245 761 30219
rect 807 10245 820 30219
rect 732 10232 820 10245
rect -820 9987 -732 10000
rect -820 -9987 -807 9987
rect -761 -9987 -732 9987
rect -820 -10000 -732 -9987
rect -612 9987 -508 10000
rect -612 -9987 -583 9987
rect -537 -9987 -508 9987
rect -612 -10000 -508 -9987
rect -388 9987 -284 10000
rect -388 -9987 -359 9987
rect -313 -9987 -284 9987
rect -388 -10000 -284 -9987
rect -164 9987 -60 10000
rect -164 -9987 -135 9987
rect -89 -9987 -60 9987
rect -164 -10000 -60 -9987
rect 60 9987 164 10000
rect 60 -9987 89 9987
rect 135 -9987 164 9987
rect 60 -10000 164 -9987
rect 284 9987 388 10000
rect 284 -9987 313 9987
rect 359 -9987 388 9987
rect 284 -10000 388 -9987
rect 508 9987 612 10000
rect 508 -9987 537 9987
rect 583 -9987 612 9987
rect 508 -10000 612 -9987
rect 732 9987 820 10000
rect 732 -9987 761 9987
rect 807 -9987 820 9987
rect 732 -10000 820 -9987
rect -820 -10245 -732 -10232
rect -820 -30219 -807 -10245
rect -761 -30219 -732 -10245
rect -820 -30232 -732 -30219
rect -612 -10245 -508 -10232
rect -612 -30219 -583 -10245
rect -537 -30219 -508 -10245
rect -612 -30232 -508 -30219
rect -388 -10245 -284 -10232
rect -388 -30219 -359 -10245
rect -313 -30219 -284 -10245
rect -388 -30232 -284 -30219
rect -164 -10245 -60 -10232
rect -164 -30219 -135 -10245
rect -89 -30219 -60 -10245
rect -164 -30232 -60 -30219
rect 60 -10245 164 -10232
rect 60 -30219 89 -10245
rect 135 -30219 164 -10245
rect 60 -30232 164 -30219
rect 284 -10245 388 -10232
rect 284 -30219 313 -10245
rect 359 -30219 388 -10245
rect 284 -30232 388 -30219
rect 508 -10245 612 -10232
rect 508 -30219 537 -10245
rect 583 -30219 612 -10245
rect 508 -30232 612 -30219
rect 732 -10245 820 -10232
rect 732 -30219 761 -10245
rect 807 -30219 820 -10245
rect 732 -30232 820 -30219
<< mvndiffc >>
rect -807 10245 -761 30219
rect -583 10245 -537 30219
rect -359 10245 -313 30219
rect -135 10245 -89 30219
rect 89 10245 135 30219
rect 313 10245 359 30219
rect 537 10245 583 30219
rect 761 10245 807 30219
rect -807 -9987 -761 9987
rect -583 -9987 -537 9987
rect -359 -9987 -313 9987
rect -135 -9987 -89 9987
rect 89 -9987 135 9987
rect 313 -9987 359 9987
rect 537 -9987 583 9987
rect 761 -9987 807 9987
rect -807 -30219 -761 -10245
rect -583 -30219 -537 -10245
rect -359 -30219 -313 -10245
rect -135 -30219 -89 -10245
rect 89 -30219 135 -10245
rect 313 -30219 359 -10245
rect 537 -30219 583 -10245
rect 761 -30219 807 -10245
<< mvpsubdiff >>
rect -964 30384 964 30456
rect -964 30340 -892 30384
rect -964 -30340 -951 30340
rect -905 -30340 -892 30340
rect 892 30340 964 30384
rect -964 -30384 -892 -30340
rect 892 -30340 905 30340
rect 951 -30340 964 30340
rect 892 -30384 964 -30340
rect -964 -30456 964 -30384
<< mvpsubdiffcont >>
rect -951 -30340 -905 30340
rect 905 -30340 951 30340
<< polysilicon >>
rect -732 30311 -612 30324
rect -732 30265 -719 30311
rect -625 30265 -612 30311
rect -732 30232 -612 30265
rect -508 30311 -388 30324
rect -508 30265 -495 30311
rect -401 30265 -388 30311
rect -508 30232 -388 30265
rect -284 30311 -164 30324
rect -284 30265 -271 30311
rect -177 30265 -164 30311
rect -284 30232 -164 30265
rect -60 30311 60 30324
rect -60 30265 -47 30311
rect 47 30265 60 30311
rect -60 30232 60 30265
rect 164 30311 284 30324
rect 164 30265 177 30311
rect 271 30265 284 30311
rect 164 30232 284 30265
rect 388 30311 508 30324
rect 388 30265 401 30311
rect 495 30265 508 30311
rect 388 30232 508 30265
rect 612 30311 732 30324
rect 612 30265 625 30311
rect 719 30265 732 30311
rect 612 30232 732 30265
rect -732 10199 -612 10232
rect -732 10153 -715 10199
rect -629 10153 -612 10199
rect -732 10079 -612 10153
rect -732 10033 -715 10079
rect -629 10033 -612 10079
rect -732 10000 -612 10033
rect -508 10199 -388 10232
rect -508 10153 -491 10199
rect -405 10153 -388 10199
rect -508 10079 -388 10153
rect -508 10033 -491 10079
rect -405 10033 -388 10079
rect -508 10000 -388 10033
rect -284 10199 -164 10232
rect -284 10153 -267 10199
rect -181 10153 -164 10199
rect -284 10079 -164 10153
rect -284 10033 -267 10079
rect -181 10033 -164 10079
rect -284 10000 -164 10033
rect -60 10199 60 10232
rect -60 10153 -43 10199
rect 43 10153 60 10199
rect -60 10079 60 10153
rect -60 10033 -43 10079
rect 43 10033 60 10079
rect -60 10000 60 10033
rect 164 10199 284 10232
rect 164 10153 181 10199
rect 267 10153 284 10199
rect 164 10079 284 10153
rect 164 10033 181 10079
rect 267 10033 284 10079
rect 164 10000 284 10033
rect 388 10199 508 10232
rect 388 10153 405 10199
rect 491 10153 508 10199
rect 388 10079 508 10153
rect 388 10033 405 10079
rect 491 10033 508 10079
rect 388 10000 508 10033
rect 612 10199 732 10232
rect 612 10153 629 10199
rect 715 10153 732 10199
rect 612 10079 732 10153
rect 612 10033 629 10079
rect 715 10033 732 10079
rect 612 10000 732 10033
rect -732 -10033 -612 -10000
rect -732 -10079 -715 -10033
rect -629 -10079 -612 -10033
rect -732 -10153 -612 -10079
rect -732 -10199 -715 -10153
rect -629 -10199 -612 -10153
rect -732 -10232 -612 -10199
rect -508 -10033 -388 -10000
rect -508 -10079 -491 -10033
rect -405 -10079 -388 -10033
rect -508 -10153 -388 -10079
rect -508 -10199 -491 -10153
rect -405 -10199 -388 -10153
rect -508 -10232 -388 -10199
rect -284 -10033 -164 -10000
rect -284 -10079 -267 -10033
rect -181 -10079 -164 -10033
rect -284 -10153 -164 -10079
rect -284 -10199 -267 -10153
rect -181 -10199 -164 -10153
rect -284 -10232 -164 -10199
rect -60 -10033 60 -10000
rect -60 -10079 -43 -10033
rect 43 -10079 60 -10033
rect -60 -10153 60 -10079
rect -60 -10199 -43 -10153
rect 43 -10199 60 -10153
rect -60 -10232 60 -10199
rect 164 -10033 284 -10000
rect 164 -10079 181 -10033
rect 267 -10079 284 -10033
rect 164 -10153 284 -10079
rect 164 -10199 181 -10153
rect 267 -10199 284 -10153
rect 164 -10232 284 -10199
rect 388 -10033 508 -10000
rect 388 -10079 405 -10033
rect 491 -10079 508 -10033
rect 388 -10153 508 -10079
rect 388 -10199 405 -10153
rect 491 -10199 508 -10153
rect 388 -10232 508 -10199
rect 612 -10033 732 -10000
rect 612 -10079 629 -10033
rect 715 -10079 732 -10033
rect 612 -10153 732 -10079
rect 612 -10199 629 -10153
rect 715 -10199 732 -10153
rect 612 -10232 732 -10199
rect -732 -30265 -612 -30232
rect -732 -30311 -719 -30265
rect -625 -30311 -612 -30265
rect -732 -30324 -612 -30311
rect -508 -30265 -388 -30232
rect -508 -30311 -495 -30265
rect -401 -30311 -388 -30265
rect -508 -30324 -388 -30311
rect -284 -30265 -164 -30232
rect -284 -30311 -271 -30265
rect -177 -30311 -164 -30265
rect -284 -30324 -164 -30311
rect -60 -30265 60 -30232
rect -60 -30311 -47 -30265
rect 47 -30311 60 -30265
rect -60 -30324 60 -30311
rect 164 -30265 284 -30232
rect 164 -30311 177 -30265
rect 271 -30311 284 -30265
rect 164 -30324 284 -30311
rect 388 -30265 508 -30232
rect 388 -30311 401 -30265
rect 495 -30311 508 -30265
rect 388 -30324 508 -30311
rect 612 -30265 732 -30232
rect 612 -30311 625 -30265
rect 719 -30311 732 -30265
rect 612 -30324 732 -30311
<< polycontact >>
rect -719 30265 -625 30311
rect -495 30265 -401 30311
rect -271 30265 -177 30311
rect -47 30265 47 30311
rect 177 30265 271 30311
rect 401 30265 495 30311
rect 625 30265 719 30311
rect -715 10153 -629 10199
rect -715 10033 -629 10079
rect -491 10153 -405 10199
rect -491 10033 -405 10079
rect -267 10153 -181 10199
rect -267 10033 -181 10079
rect -43 10153 43 10199
rect -43 10033 43 10079
rect 181 10153 267 10199
rect 181 10033 267 10079
rect 405 10153 491 10199
rect 405 10033 491 10079
rect 629 10153 715 10199
rect 629 10033 715 10079
rect -715 -10079 -629 -10033
rect -715 -10199 -629 -10153
rect -491 -10079 -405 -10033
rect -491 -10199 -405 -10153
rect -267 -10079 -181 -10033
rect -267 -10199 -181 -10153
rect -43 -10079 43 -10033
rect -43 -10199 43 -10153
rect 181 -10079 267 -10033
rect 181 -10199 267 -10153
rect 405 -10079 491 -10033
rect 405 -10199 491 -10153
rect 629 -10079 715 -10033
rect 629 -10199 715 -10153
rect -719 -30311 -625 -30265
rect -495 -30311 -401 -30265
rect -271 -30311 -177 -30265
rect -47 -30311 47 -30265
rect 177 -30311 271 -30265
rect 401 -30311 495 -30265
rect 625 -30311 719 -30265
<< metal1 >>
rect -951 30397 951 30443
rect -951 30340 -905 30397
rect -730 30311 730 30351
rect -730 30265 -719 30311
rect -625 30302 -495 30311
rect -625 30265 -614 30302
rect -506 30265 -495 30302
rect -401 30302 -271 30311
rect -401 30265 -390 30302
rect -282 30265 -271 30302
rect -177 30302 -47 30311
rect -177 30265 -166 30302
rect -58 30265 -47 30302
rect 47 30302 177 30311
rect 47 30265 58 30302
rect 166 30265 177 30302
rect 271 30302 401 30311
rect 271 30265 282 30302
rect 390 30265 401 30302
rect 495 30302 625 30311
rect 495 30265 506 30302
rect 614 30265 625 30302
rect 719 30265 730 30311
rect 905 30340 951 30397
rect -807 30219 -761 30230
rect -807 9987 -761 10245
rect -583 30219 -537 30230
rect -715 10199 -629 10210
rect -715 10079 -629 10153
rect -715 10022 -629 10033
rect -807 -10245 -761 -9987
rect -583 9987 -537 10245
rect -359 30219 -313 30230
rect -491 10199 -405 10210
rect -491 10079 -405 10153
rect -491 10022 -405 10033
rect -715 -10033 -629 -10022
rect -715 -10153 -629 -10079
rect -715 -10210 -629 -10199
rect -807 -30230 -761 -30219
rect -583 -10245 -537 -9987
rect -359 9987 -313 10245
rect -135 30219 -89 30230
rect -267 10199 -181 10210
rect -267 10079 -181 10153
rect -267 10022 -181 10033
rect -491 -10033 -405 -10022
rect -491 -10153 -405 -10079
rect -491 -10210 -405 -10199
rect -583 -30230 -537 -30219
rect -359 -10245 -313 -9987
rect -135 9987 -89 10245
rect 89 30219 135 30230
rect -43 10199 43 10210
rect -43 10079 43 10153
rect -43 10022 43 10033
rect -267 -10033 -181 -10022
rect -267 -10153 -181 -10079
rect -267 -10210 -181 -10199
rect -359 -30230 -313 -30219
rect -135 -10245 -89 -9987
rect 89 9987 135 10245
rect 313 30219 359 30230
rect 181 10199 267 10210
rect 181 10079 267 10153
rect 181 10022 267 10033
rect -43 -10033 43 -10022
rect -43 -10153 43 -10079
rect -43 -10210 43 -10199
rect -135 -30230 -89 -30219
rect 89 -10245 135 -9987
rect 313 9987 359 10245
rect 537 30219 583 30230
rect 405 10199 491 10210
rect 405 10079 491 10153
rect 405 10022 491 10033
rect 181 -10033 267 -10022
rect 181 -10153 267 -10079
rect 181 -10210 267 -10199
rect 89 -30230 135 -30219
rect 313 -10245 359 -9987
rect 537 9987 583 10245
rect 761 30219 807 30230
rect 629 10199 715 10210
rect 629 10079 715 10153
rect 629 10022 715 10033
rect 405 -10033 491 -10022
rect 405 -10153 491 -10079
rect 405 -10210 491 -10199
rect 313 -30230 359 -30219
rect 537 -10245 583 -9987
rect 761 9987 807 10245
rect 629 -10033 715 -10022
rect 629 -10153 715 -10079
rect 629 -10210 715 -10199
rect 537 -30230 583 -30219
rect 761 -10245 807 -9987
rect 761 -30230 807 -30219
rect -951 -30397 -905 -30340
rect -730 -30311 -719 -30265
rect -625 -30302 -614 -30265
rect -506 -30302 -495 -30265
rect -625 -30311 -495 -30302
rect -401 -30302 -390 -30265
rect -282 -30302 -271 -30265
rect -401 -30311 -271 -30302
rect -177 -30302 -166 -30265
rect -58 -30302 -47 -30265
rect -177 -30311 -47 -30302
rect 47 -30302 58 -30265
rect 166 -30302 177 -30265
rect 47 -30311 177 -30302
rect 271 -30302 282 -30265
rect 390 -30302 401 -30265
rect 271 -30311 401 -30302
rect 495 -30302 506 -30265
rect 614 -30302 625 -30265
rect 495 -30311 625 -30302
rect 719 -30311 730 -30265
rect -730 -30351 730 -30311
rect 905 -30397 951 -30340
rect -951 -30443 951 -30397
<< properties >>
string FIXED_BBOX -928 -30420 928 30420
string gencell nfet_06v0
string library gf180mcu
string parameters w 100.0 l 0.6 m 3 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.6 wmin 0.3 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
