module aef2;
endmodule
