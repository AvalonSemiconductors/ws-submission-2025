`default_nettype none

module tholin_img(
	input [7:0] column,
	input [6:0] row,
	output [4:0] pixel
);

reg [4:0] rom;
assign pixel = rom;
always @(*) begin
	case({column, row})
		default: rom = 5'hxx;
		0: rom = 31;
		1: rom = 31;
		2: rom = 31;
		3: rom = 31;
		4: rom = 31;
		5: rom = 31;
		6: rom = 31;
		7: rom = 31;
		8: rom = 31;
		9: rom = 31;
		10: rom = 31;
		11: rom = 31;
		12: rom = 31;
		13: rom = 31;
		14: rom = 31;
		15: rom = 31;
		16: rom = 31;
		17: rom = 31;
		18: rom = 31;
		19: rom = 31;
		20: rom = 31;
		21: rom = 31;
		22: rom = 31;
		23: rom = 31;
		24: rom = 31;
		25: rom = 31;
		26: rom = 31;
		27: rom = 31;
		28: rom = 31;
		29: rom = 31;
		30: rom = 31;
		31: rom = 31;
		32: rom = 31;
		33: rom = 31;
		34: rom = 31;
		35: rom = 31;
		36: rom = 31;
		37: rom = 31;
		38: rom = 31;
		39: rom = 31;
		40: rom = 31;
		41: rom = 31;
		42: rom = 31;
		43: rom = 31;
		44: rom = 31;
		45: rom = 31;
		46: rom = 31;
		47: rom = 31;
		48: rom = 31;
		49: rom = 31;
		50: rom = 31;
		51: rom = 31;
		52: rom = 31;
		53: rom = 31;
		54: rom = 31;
		55: rom = 31;
		56: rom = 31;
		57: rom = 31;
		58: rom = 31;
		59: rom = 31;
		60: rom = 31;
		61: rom = 31;
		62: rom = 31;
		63: rom = 31;
		64: rom = 31;
		65: rom = 31;
		66: rom = 31;
		67: rom = 31;
		68: rom = 31;
		69: rom = 31;
		70: rom = 31;
		71: rom = 31;
		72: rom = 31;
		73: rom = 31;
		74: rom = 31;
		75: rom = 31;
		76: rom = 31;
		77: rom = 31;
		78: rom = 31;
		79: rom = 31;
		80: rom = 31;
		81: rom = 31;
		82: rom = 31;
		83: rom = 31;
		84: rom = 31;
		85: rom = 31;
		86: rom = 31;
		87: rom = 31;
		88: rom = 31;
		89: rom = 31;
		90: rom = 31;
		91: rom = 31;
		92: rom = 31;
		93: rom = 31;
		94: rom = 31;
		95: rom = 31;
		96: rom = 31;
		97: rom = 31;
		98: rom = 31;
		99: rom = 31;
		100: rom = 31;
		101: rom = 31;
		102: rom = 31;
		103: rom = 31;
		104: rom = 31;
		105: rom = 31;
		106: rom = 31;
		107: rom = 31;
		108: rom = 31;
		109: rom = 31;
		110: rom = 31;
		111: rom = 31;
		112: rom = 31;
		113: rom = 31;
		114: rom = 31;
		115: rom = 31;
		116: rom = 31;
		117: rom = 31;
		118: rom = 31;
		119: rom = 31;
		120: rom = 31;
		121: rom = 31;
		122: rom = 31;
		128: rom = 31;
		129: rom = 31;
		130: rom = 31;
		131: rom = 31;
		132: rom = 31;
		133: rom = 31;
		134: rom = 31;
		135: rom = 31;
		136: rom = 31;
		137: rom = 31;
		138: rom = 31;
		139: rom = 31;
		140: rom = 31;
		141: rom = 31;
		142: rom = 31;
		143: rom = 31;
		144: rom = 31;
		145: rom = 31;
		146: rom = 31;
		147: rom = 31;
		148: rom = 31;
		149: rom = 31;
		150: rom = 31;
		151: rom = 31;
		152: rom = 31;
		153: rom = 31;
		154: rom = 31;
		155: rom = 31;
		156: rom = 31;
		157: rom = 31;
		158: rom = 31;
		159: rom = 31;
		160: rom = 31;
		161: rom = 31;
		162: rom = 31;
		163: rom = 31;
		164: rom = 31;
		165: rom = 31;
		166: rom = 31;
		167: rom = 31;
		168: rom = 31;
		169: rom = 31;
		170: rom = 31;
		171: rom = 31;
		172: rom = 31;
		173: rom = 31;
		174: rom = 31;
		175: rom = 31;
		176: rom = 31;
		177: rom = 31;
		178: rom = 31;
		179: rom = 31;
		180: rom = 31;
		181: rom = 31;
		182: rom = 31;
		183: rom = 31;
		184: rom = 31;
		185: rom = 31;
		186: rom = 31;
		187: rom = 31;
		188: rom = 31;
		189: rom = 31;
		190: rom = 31;
		191: rom = 31;
		192: rom = 31;
		193: rom = 31;
		194: rom = 31;
		195: rom = 31;
		196: rom = 31;
		197: rom = 31;
		198: rom = 31;
		199: rom = 31;
		200: rom = 31;
		201: rom = 31;
		202: rom = 31;
		203: rom = 31;
		204: rom = 31;
		205: rom = 31;
		206: rom = 31;
		207: rom = 31;
		208: rom = 31;
		209: rom = 31;
		210: rom = 31;
		211: rom = 31;
		212: rom = 31;
		213: rom = 31;
		214: rom = 31;
		215: rom = 31;
		216: rom = 31;
		217: rom = 31;
		218: rom = 31;
		219: rom = 31;
		220: rom = 31;
		221: rom = 31;
		222: rom = 31;
		223: rom = 31;
		224: rom = 31;
		225: rom = 31;
		226: rom = 31;
		227: rom = 31;
		228: rom = 31;
		229: rom = 31;
		230: rom = 31;
		231: rom = 31;
		232: rom = 31;
		233: rom = 31;
		234: rom = 31;
		235: rom = 31;
		236: rom = 31;
		237: rom = 31;
		238: rom = 31;
		239: rom = 31;
		240: rom = 31;
		241: rom = 31;
		242: rom = 31;
		243: rom = 31;
		244: rom = 31;
		245: rom = 31;
		246: rom = 31;
		247: rom = 31;
		248: rom = 31;
		249: rom = 31;
		250: rom = 31;
		256: rom = 31;
		257: rom = 31;
		258: rom = 31;
		259: rom = 31;
		260: rom = 31;
		261: rom = 31;
		262: rom = 31;
		263: rom = 31;
		264: rom = 31;
		265: rom = 31;
		266: rom = 31;
		267: rom = 31;
		268: rom = 31;
		269: rom = 31;
		270: rom = 31;
		271: rom = 31;
		272: rom = 31;
		273: rom = 31;
		274: rom = 31;
		275: rom = 31;
		276: rom = 31;
		277: rom = 31;
		278: rom = 31;
		279: rom = 31;
		280: rom = 31;
		281: rom = 31;
		282: rom = 31;
		283: rom = 31;
		284: rom = 31;
		285: rom = 31;
		286: rom = 31;
		287: rom = 31;
		288: rom = 31;
		289: rom = 31;
		290: rom = 31;
		291: rom = 31;
		292: rom = 31;
		293: rom = 31;
		294: rom = 31;
		295: rom = 31;
		296: rom = 31;
		297: rom = 31;
		298: rom = 31;
		299: rom = 31;
		300: rom = 31;
		301: rom = 31;
		302: rom = 31;
		303: rom = 31;
		304: rom = 31;
		305: rom = 31;
		306: rom = 31;
		307: rom = 31;
		308: rom = 31;
		309: rom = 31;
		310: rom = 31;
		311: rom = 31;
		312: rom = 31;
		313: rom = 31;
		314: rom = 31;
		315: rom = 31;
		316: rom = 31;
		317: rom = 31;
		318: rom = 31;
		319: rom = 31;
		320: rom = 31;
		321: rom = 31;
		322: rom = 31;
		323: rom = 31;
		324: rom = 31;
		325: rom = 31;
		326: rom = 31;
		327: rom = 31;
		328: rom = 31;
		329: rom = 31;
		330: rom = 31;
		331: rom = 31;
		332: rom = 31;
		333: rom = 31;
		334: rom = 31;
		335: rom = 31;
		336: rom = 31;
		337: rom = 31;
		338: rom = 31;
		339: rom = 31;
		340: rom = 31;
		341: rom = 31;
		342: rom = 31;
		343: rom = 31;
		344: rom = 31;
		345: rom = 31;
		346: rom = 31;
		347: rom = 31;
		348: rom = 31;
		349: rom = 31;
		350: rom = 31;
		351: rom = 31;
		352: rom = 31;
		353: rom = 31;
		354: rom = 31;
		355: rom = 31;
		356: rom = 31;
		357: rom = 31;
		358: rom = 31;
		359: rom = 31;
		360: rom = 31;
		361: rom = 31;
		362: rom = 31;
		363: rom = 31;
		364: rom = 31;
		365: rom = 31;
		366: rom = 31;
		367: rom = 31;
		368: rom = 31;
		369: rom = 31;
		370: rom = 31;
		371: rom = 31;
		372: rom = 31;
		373: rom = 31;
		374: rom = 31;
		375: rom = 31;
		376: rom = 31;
		377: rom = 31;
		378: rom = 31;
		384: rom = 31;
		385: rom = 31;
		386: rom = 31;
		387: rom = 31;
		388: rom = 31;
		389: rom = 31;
		390: rom = 31;
		391: rom = 31;
		392: rom = 31;
		393: rom = 31;
		394: rom = 31;
		395: rom = 31;
		396: rom = 31;
		397: rom = 31;
		398: rom = 31;
		399: rom = 31;
		400: rom = 31;
		401: rom = 31;
		402: rom = 31;
		403: rom = 31;
		404: rom = 31;
		405: rom = 31;
		406: rom = 31;
		407: rom = 31;
		408: rom = 31;
		409: rom = 31;
		410: rom = 31;
		411: rom = 31;
		412: rom = 31;
		413: rom = 31;
		414: rom = 31;
		415: rom = 31;
		416: rom = 31;
		417: rom = 31;
		418: rom = 31;
		419: rom = 31;
		420: rom = 31;
		421: rom = 31;
		422: rom = 31;
		423: rom = 31;
		424: rom = 31;
		425: rom = 31;
		426: rom = 31;
		427: rom = 31;
		428: rom = 31;
		429: rom = 31;
		430: rom = 31;
		431: rom = 31;
		432: rom = 31;
		433: rom = 31;
		434: rom = 31;
		435: rom = 31;
		436: rom = 31;
		437: rom = 31;
		438: rom = 31;
		439: rom = 31;
		440: rom = 31;
		441: rom = 31;
		442: rom = 31;
		443: rom = 31;
		444: rom = 31;
		445: rom = 31;
		446: rom = 31;
		447: rom = 31;
		448: rom = 31;
		449: rom = 31;
		450: rom = 31;
		451: rom = 31;
		452: rom = 31;
		453: rom = 31;
		454: rom = 31;
		455: rom = 31;
		456: rom = 31;
		457: rom = 31;
		458: rom = 31;
		459: rom = 31;
		460: rom = 31;
		461: rom = 31;
		462: rom = 31;
		463: rom = 31;
		464: rom = 31;
		465: rom = 31;
		466: rom = 31;
		467: rom = 31;
		468: rom = 31;
		469: rom = 31;
		470: rom = 31;
		471: rom = 31;
		472: rom = 31;
		473: rom = 31;
		474: rom = 31;
		475: rom = 31;
		476: rom = 31;
		477: rom = 31;
		478: rom = 31;
		479: rom = 31;
		480: rom = 31;
		481: rom = 31;
		482: rom = 31;
		483: rom = 31;
		484: rom = 31;
		485: rom = 31;
		486: rom = 31;
		487: rom = 31;
		488: rom = 31;
		489: rom = 31;
		490: rom = 31;
		491: rom = 31;
		492: rom = 31;
		493: rom = 31;
		494: rom = 31;
		495: rom = 31;
		496: rom = 31;
		497: rom = 31;
		498: rom = 31;
		499: rom = 31;
		500: rom = 31;
		501: rom = 31;
		502: rom = 31;
		503: rom = 31;
		504: rom = 31;
		505: rom = 31;
		506: rom = 31;
		512: rom = 31;
		513: rom = 31;
		514: rom = 31;
		515: rom = 31;
		516: rom = 31;
		517: rom = 31;
		518: rom = 31;
		519: rom = 31;
		520: rom = 31;
		521: rom = 31;
		522: rom = 31;
		523: rom = 31;
		524: rom = 31;
		525: rom = 31;
		526: rom = 31;
		527: rom = 31;
		528: rom = 31;
		529: rom = 31;
		530: rom = 31;
		531: rom = 31;
		532: rom = 31;
		533: rom = 31;
		534: rom = 31;
		535: rom = 31;
		536: rom = 31;
		537: rom = 31;
		538: rom = 31;
		539: rom = 31;
		540: rom = 31;
		541: rom = 31;
		542: rom = 31;
		543: rom = 31;
		544: rom = 31;
		545: rom = 31;
		546: rom = 31;
		547: rom = 31;
		548: rom = 31;
		549: rom = 31;
		550: rom = 31;
		551: rom = 31;
		552: rom = 31;
		553: rom = 31;
		554: rom = 31;
		555: rom = 31;
		556: rom = 31;
		557: rom = 31;
		558: rom = 31;
		559: rom = 31;
		560: rom = 31;
		561: rom = 31;
		562: rom = 31;
		563: rom = 31;
		564: rom = 31;
		565: rom = 31;
		566: rom = 31;
		567: rom = 31;
		568: rom = 31;
		569: rom = 31;
		570: rom = 31;
		571: rom = 31;
		572: rom = 31;
		573: rom = 31;
		574: rom = 31;
		575: rom = 31;
		576: rom = 31;
		577: rom = 31;
		578: rom = 31;
		579: rom = 31;
		580: rom = 31;
		581: rom = 31;
		582: rom = 31;
		583: rom = 31;
		584: rom = 31;
		585: rom = 31;
		586: rom = 31;
		587: rom = 31;
		588: rom = 31;
		589: rom = 31;
		590: rom = 31;
		591: rom = 31;
		592: rom = 31;
		593: rom = 31;
		594: rom = 31;
		595: rom = 31;
		596: rom = 31;
		597: rom = 31;
		598: rom = 31;
		599: rom = 31;
		600: rom = 31;
		601: rom = 31;
		602: rom = 31;
		603: rom = 31;
		604: rom = 31;
		605: rom = 31;
		606: rom = 31;
		607: rom = 31;
		608: rom = 31;
		609: rom = 31;
		610: rom = 31;
		611: rom = 31;
		612: rom = 31;
		613: rom = 31;
		614: rom = 31;
		615: rom = 31;
		616: rom = 31;
		617: rom = 31;
		618: rom = 31;
		619: rom = 31;
		620: rom = 31;
		621: rom = 31;
		622: rom = 31;
		623: rom = 31;
		624: rom = 31;
		625: rom = 31;
		626: rom = 31;
		627: rom = 31;
		628: rom = 31;
		629: rom = 31;
		630: rom = 31;
		631: rom = 31;
		632: rom = 31;
		633: rom = 31;
		634: rom = 31;
		640: rom = 31;
		641: rom = 31;
		642: rom = 31;
		643: rom = 31;
		644: rom = 31;
		645: rom = 31;
		646: rom = 31;
		647: rom = 31;
		648: rom = 31;
		649: rom = 31;
		650: rom = 31;
		651: rom = 31;
		652: rom = 31;
		653: rom = 31;
		654: rom = 31;
		655: rom = 31;
		656: rom = 31;
		657: rom = 31;
		658: rom = 31;
		659: rom = 31;
		660: rom = 31;
		661: rom = 31;
		662: rom = 31;
		663: rom = 31;
		664: rom = 31;
		665: rom = 31;
		666: rom = 31;
		667: rom = 31;
		668: rom = 31;
		669: rom = 31;
		670: rom = 31;
		671: rom = 31;
		672: rom = 31;
		673: rom = 31;
		674: rom = 31;
		675: rom = 31;
		676: rom = 31;
		677: rom = 31;
		678: rom = 31;
		679: rom = 31;
		680: rom = 31;
		681: rom = 31;
		682: rom = 31;
		683: rom = 31;
		684: rom = 31;
		685: rom = 31;
		686: rom = 31;
		687: rom = 31;
		688: rom = 31;
		689: rom = 31;
		690: rom = 31;
		691: rom = 31;
		692: rom = 31;
		693: rom = 31;
		694: rom = 31;
		695: rom = 31;
		696: rom = 31;
		697: rom = 31;
		698: rom = 31;
		699: rom = 31;
		700: rom = 31;
		701: rom = 31;
		702: rom = 31;
		703: rom = 31;
		704: rom = 31;
		705: rom = 31;
		706: rom = 31;
		707: rom = 31;
		708: rom = 31;
		709: rom = 31;
		710: rom = 31;
		711: rom = 31;
		712: rom = 31;
		713: rom = 31;
		714: rom = 31;
		715: rom = 31;
		716: rom = 31;
		717: rom = 31;
		718: rom = 31;
		719: rom = 31;
		720: rom = 31;
		721: rom = 31;
		722: rom = 31;
		723: rom = 31;
		724: rom = 31;
		725: rom = 31;
		726: rom = 31;
		727: rom = 31;
		728: rom = 31;
		729: rom = 31;
		730: rom = 31;
		731: rom = 31;
		732: rom = 31;
		733: rom = 31;
		734: rom = 31;
		735: rom = 31;
		736: rom = 31;
		737: rom = 31;
		738: rom = 31;
		739: rom = 31;
		740: rom = 31;
		741: rom = 31;
		742: rom = 31;
		743: rom = 31;
		744: rom = 31;
		745: rom = 31;
		746: rom = 31;
		747: rom = 31;
		748: rom = 31;
		749: rom = 31;
		750: rom = 31;
		751: rom = 31;
		752: rom = 31;
		753: rom = 31;
		754: rom = 31;
		755: rom = 31;
		756: rom = 31;
		757: rom = 31;
		758: rom = 31;
		759: rom = 31;
		760: rom = 31;
		761: rom = 31;
		762: rom = 31;
		768: rom = 31;
		769: rom = 31;
		770: rom = 31;
		771: rom = 31;
		772: rom = 31;
		773: rom = 31;
		774: rom = 31;
		775: rom = 31;
		776: rom = 31;
		777: rom = 31;
		778: rom = 31;
		779: rom = 31;
		780: rom = 31;
		781: rom = 31;
		782: rom = 31;
		783: rom = 31;
		784: rom = 31;
		785: rom = 31;
		786: rom = 31;
		787: rom = 31;
		788: rom = 31;
		789: rom = 31;
		790: rom = 31;
		791: rom = 31;
		792: rom = 31;
		793: rom = 31;
		794: rom = 31;
		795: rom = 31;
		796: rom = 31;
		797: rom = 31;
		798: rom = 31;
		799: rom = 31;
		800: rom = 31;
		801: rom = 31;
		802: rom = 31;
		803: rom = 31;
		804: rom = 31;
		805: rom = 31;
		806: rom = 31;
		807: rom = 31;
		808: rom = 31;
		809: rom = 31;
		810: rom = 31;
		811: rom = 31;
		812: rom = 31;
		813: rom = 31;
		814: rom = 31;
		815: rom = 31;
		816: rom = 31;
		817: rom = 31;
		818: rom = 31;
		819: rom = 31;
		820: rom = 31;
		821: rom = 31;
		822: rom = 31;
		823: rom = 31;
		824: rom = 31;
		825: rom = 31;
		826: rom = 31;
		827: rom = 31;
		828: rom = 31;
		829: rom = 31;
		830: rom = 31;
		831: rom = 31;
		832: rom = 31;
		833: rom = 31;
		834: rom = 31;
		835: rom = 31;
		836: rom = 31;
		837: rom = 31;
		838: rom = 31;
		839: rom = 31;
		840: rom = 31;
		841: rom = 31;
		842: rom = 31;
		843: rom = 31;
		844: rom = 31;
		845: rom = 31;
		846: rom = 31;
		847: rom = 31;
		848: rom = 31;
		849: rom = 31;
		850: rom = 31;
		851: rom = 31;
		852: rom = 31;
		853: rom = 31;
		854: rom = 31;
		855: rom = 31;
		856: rom = 31;
		857: rom = 31;
		858: rom = 31;
		859: rom = 31;
		860: rom = 31;
		861: rom = 31;
		862: rom = 31;
		863: rom = 31;
		864: rom = 31;
		865: rom = 31;
		866: rom = 31;
		867: rom = 31;
		868: rom = 31;
		869: rom = 31;
		870: rom = 31;
		871: rom = 31;
		872: rom = 31;
		873: rom = 31;
		874: rom = 31;
		875: rom = 31;
		876: rom = 31;
		877: rom = 31;
		878: rom = 31;
		879: rom = 31;
		880: rom = 31;
		881: rom = 31;
		882: rom = 31;
		883: rom = 31;
		884: rom = 31;
		885: rom = 31;
		886: rom = 31;
		887: rom = 31;
		888: rom = 31;
		889: rom = 31;
		890: rom = 31;
		896: rom = 31;
		897: rom = 31;
		898: rom = 31;
		899: rom = 31;
		900: rom = 31;
		901: rom = 31;
		902: rom = 31;
		903: rom = 31;
		904: rom = 31;
		905: rom = 31;
		906: rom = 31;
		907: rom = 31;
		908: rom = 31;
		909: rom = 31;
		910: rom = 31;
		911: rom = 31;
		912: rom = 31;
		913: rom = 31;
		914: rom = 31;
		915: rom = 31;
		916: rom = 31;
		917: rom = 31;
		918: rom = 31;
		919: rom = 31;
		920: rom = 31;
		921: rom = 31;
		922: rom = 31;
		923: rom = 31;
		924: rom = 31;
		925: rom = 31;
		926: rom = 31;
		927: rom = 31;
		928: rom = 31;
		929: rom = 31;
		930: rom = 31;
		931: rom = 31;
		932: rom = 31;
		933: rom = 31;
		934: rom = 31;
		935: rom = 31;
		936: rom = 31;
		937: rom = 31;
		938: rom = 31;
		939: rom = 31;
		940: rom = 31;
		941: rom = 31;
		942: rom = 31;
		943: rom = 31;
		944: rom = 31;
		945: rom = 31;
		946: rom = 31;
		947: rom = 31;
		948: rom = 31;
		949: rom = 31;
		950: rom = 31;
		951: rom = 31;
		952: rom = 31;
		953: rom = 31;
		954: rom = 31;
		955: rom = 31;
		956: rom = 31;
		957: rom = 31;
		958: rom = 31;
		959: rom = 31;
		960: rom = 31;
		961: rom = 31;
		962: rom = 31;
		963: rom = 31;
		964: rom = 31;
		965: rom = 31;
		966: rom = 31;
		967: rom = 31;
		968: rom = 31;
		969: rom = 31;
		970: rom = 31;
		971: rom = 31;
		972: rom = 31;
		973: rom = 31;
		974: rom = 31;
		975: rom = 31;
		976: rom = 31;
		977: rom = 31;
		978: rom = 31;
		979: rom = 31;
		980: rom = 31;
		981: rom = 31;
		982: rom = 31;
		983: rom = 31;
		984: rom = 31;
		985: rom = 31;
		986: rom = 31;
		987: rom = 31;
		988: rom = 31;
		989: rom = 31;
		990: rom = 31;
		991: rom = 31;
		992: rom = 31;
		993: rom = 31;
		994: rom = 31;
		995: rom = 31;
		996: rom = 31;
		997: rom = 31;
		998: rom = 31;
		999: rom = 31;
		1000: rom = 31;
		1001: rom = 31;
		1002: rom = 31;
		1003: rom = 31;
		1004: rom = 31;
		1005: rom = 31;
		1006: rom = 31;
		1007: rom = 31;
		1008: rom = 31;
		1009: rom = 31;
		1010: rom = 31;
		1011: rom = 31;
		1012: rom = 31;
		1013: rom = 31;
		1014: rom = 31;
		1015: rom = 31;
		1016: rom = 31;
		1017: rom = 31;
		1018: rom = 31;
		1024: rom = 31;
		1025: rom = 31;
		1026: rom = 31;
		1027: rom = 31;
		1028: rom = 31;
		1029: rom = 31;
		1030: rom = 31;
		1031: rom = 31;
		1032: rom = 31;
		1033: rom = 31;
		1034: rom = 31;
		1035: rom = 31;
		1036: rom = 31;
		1037: rom = 31;
		1038: rom = 31;
		1039: rom = 31;
		1040: rom = 31;
		1041: rom = 31;
		1042: rom = 31;
		1043: rom = 31;
		1044: rom = 31;
		1045: rom = 31;
		1046: rom = 31;
		1047: rom = 31;
		1048: rom = 31;
		1049: rom = 31;
		1050: rom = 31;
		1051: rom = 31;
		1052: rom = 31;
		1053: rom = 31;
		1054: rom = 31;
		1055: rom = 31;
		1056: rom = 31;
		1057: rom = 31;
		1058: rom = 31;
		1059: rom = 31;
		1060: rom = 31;
		1061: rom = 31;
		1062: rom = 31;
		1063: rom = 31;
		1064: rom = 31;
		1065: rom = 31;
		1066: rom = 31;
		1067: rom = 31;
		1068: rom = 31;
		1069: rom = 31;
		1070: rom = 31;
		1071: rom = 31;
		1072: rom = 31;
		1073: rom = 31;
		1074: rom = 31;
		1075: rom = 31;
		1076: rom = 31;
		1077: rom = 31;
		1078: rom = 31;
		1079: rom = 31;
		1080: rom = 31;
		1081: rom = 31;
		1082: rom = 31;
		1083: rom = 31;
		1084: rom = 31;
		1085: rom = 31;
		1086: rom = 31;
		1087: rom = 31;
		1088: rom = 31;
		1089: rom = 31;
		1090: rom = 31;
		1091: rom = 31;
		1092: rom = 31;
		1093: rom = 31;
		1094: rom = 31;
		1095: rom = 31;
		1096: rom = 31;
		1097: rom = 31;
		1098: rom = 31;
		1099: rom = 31;
		1100: rom = 31;
		1101: rom = 31;
		1102: rom = 31;
		1103: rom = 31;
		1104: rom = 31;
		1105: rom = 31;
		1106: rom = 31;
		1107: rom = 31;
		1108: rom = 31;
		1109: rom = 31;
		1110: rom = 31;
		1111: rom = 31;
		1112: rom = 31;
		1113: rom = 31;
		1114: rom = 31;
		1115: rom = 31;
		1116: rom = 31;
		1117: rom = 31;
		1118: rom = 31;
		1119: rom = 31;
		1120: rom = 31;
		1121: rom = 31;
		1122: rom = 31;
		1123: rom = 31;
		1124: rom = 31;
		1125: rom = 31;
		1126: rom = 31;
		1127: rom = 31;
		1128: rom = 31;
		1129: rom = 31;
		1130: rom = 31;
		1131: rom = 31;
		1132: rom = 31;
		1133: rom = 31;
		1134: rom = 31;
		1135: rom = 31;
		1136: rom = 31;
		1137: rom = 31;
		1138: rom = 31;
		1139: rom = 31;
		1140: rom = 31;
		1141: rom = 31;
		1142: rom = 31;
		1143: rom = 31;
		1144: rom = 31;
		1145: rom = 31;
		1146: rom = 31;
		1152: rom = 27;
		1153: rom = 27;
		1154: rom = 27;
		1155: rom = 27;
		1156: rom = 27;
		1157: rom = 27;
		1158: rom = 27;
		1159: rom = 27;
		1160: rom = 27;
		1161: rom = 27;
		1162: rom = 27;
		1163: rom = 27;
		1164: rom = 27;
		1165: rom = 27;
		1166: rom = 27;
		1167: rom = 27;
		1168: rom = 27;
		1169: rom = 27;
		1170: rom = 27;
		1171: rom = 27;
		1172: rom = 27;
		1173: rom = 27;
		1174: rom = 27;
		1175: rom = 27;
		1176: rom = 27;
		1177: rom = 27;
		1178: rom = 27;
		1179: rom = 27;
		1180: rom = 27;
		1181: rom = 27;
		1182: rom = 27;
		1183: rom = 27;
		1184: rom = 27;
		1185: rom = 27;
		1186: rom = 27;
		1187: rom = 27;
		1188: rom = 27;
		1189: rom = 27;
		1190: rom = 27;
		1191: rom = 27;
		1192: rom = 27;
		1193: rom = 27;
		1194: rom = 27;
		1195: rom = 27;
		1196: rom = 27;
		1197: rom = 27;
		1198: rom = 27;
		1199: rom = 27;
		1200: rom = 27;
		1201: rom = 27;
		1202: rom = 27;
		1203: rom = 27;
		1204: rom = 27;
		1205: rom = 27;
		1206: rom = 27;
		1207: rom = 27;
		1208: rom = 27;
		1209: rom = 27;
		1210: rom = 27;
		1211: rom = 27;
		1212: rom = 27;
		1213: rom = 27;
		1214: rom = 27;
		1215: rom = 27;
		1216: rom = 27;
		1217: rom = 27;
		1218: rom = 27;
		1219: rom = 27;
		1220: rom = 27;
		1221: rom = 27;
		1222: rom = 27;
		1223: rom = 27;
		1224: rom = 27;
		1225: rom = 27;
		1226: rom = 27;
		1227: rom = 27;
		1228: rom = 27;
		1229: rom = 27;
		1230: rom = 27;
		1231: rom = 27;
		1232: rom = 27;
		1233: rom = 27;
		1234: rom = 27;
		1235: rom = 27;
		1236: rom = 27;
		1237: rom = 27;
		1238: rom = 27;
		1239: rom = 27;
		1240: rom = 27;
		1241: rom = 27;
		1242: rom = 27;
		1243: rom = 27;
		1244: rom = 27;
		1245: rom = 27;
		1246: rom = 27;
		1247: rom = 27;
		1248: rom = 27;
		1249: rom = 27;
		1250: rom = 27;
		1251: rom = 27;
		1252: rom = 27;
		1253: rom = 27;
		1254: rom = 27;
		1255: rom = 27;
		1256: rom = 27;
		1257: rom = 27;
		1258: rom = 27;
		1259: rom = 27;
		1260: rom = 27;
		1261: rom = 27;
		1262: rom = 27;
		1263: rom = 27;
		1264: rom = 27;
		1265: rom = 27;
		1266: rom = 27;
		1267: rom = 27;
		1268: rom = 27;
		1269: rom = 27;
		1270: rom = 27;
		1271: rom = 27;
		1272: rom = 27;
		1273: rom = 27;
		1274: rom = 27;
		1280: rom = 27;
		1281: rom = 27;
		1282: rom = 27;
		1283: rom = 27;
		1284: rom = 27;
		1285: rom = 27;
		1286: rom = 27;
		1287: rom = 23;
		1288: rom = 26;
		1289: rom = 27;
		1290: rom = 27;
		1291: rom = 27;
		1292: rom = 27;
		1293: rom = 27;
		1294: rom = 27;
		1295: rom = 27;
		1296: rom = 27;
		1297: rom = 27;
		1298: rom = 27;
		1299: rom = 27;
		1300: rom = 27;
		1301: rom = 27;
		1302: rom = 27;
		1303: rom = 27;
		1304: rom = 27;
		1305: rom = 27;
		1306: rom = 27;
		1307: rom = 27;
		1308: rom = 27;
		1309: rom = 27;
		1310: rom = 27;
		1311: rom = 27;
		1312: rom = 27;
		1313: rom = 27;
		1314: rom = 27;
		1315: rom = 27;
		1316: rom = 27;
		1317: rom = 27;
		1318: rom = 27;
		1319: rom = 27;
		1320: rom = 27;
		1321: rom = 27;
		1322: rom = 27;
		1323: rom = 27;
		1324: rom = 27;
		1325: rom = 27;
		1326: rom = 27;
		1327: rom = 27;
		1328: rom = 27;
		1329: rom = 27;
		1330: rom = 27;
		1331: rom = 27;
		1332: rom = 27;
		1333: rom = 27;
		1334: rom = 27;
		1335: rom = 27;
		1336: rom = 27;
		1337: rom = 27;
		1338: rom = 27;
		1339: rom = 27;
		1340: rom = 27;
		1341: rom = 27;
		1342: rom = 27;
		1343: rom = 27;
		1344: rom = 27;
		1345: rom = 27;
		1346: rom = 27;
		1347: rom = 27;
		1348: rom = 27;
		1349: rom = 27;
		1350: rom = 27;
		1351: rom = 27;
		1352: rom = 27;
		1353: rom = 27;
		1354: rom = 27;
		1355: rom = 27;
		1356: rom = 27;
		1357: rom = 27;
		1358: rom = 27;
		1359: rom = 27;
		1360: rom = 27;
		1361: rom = 27;
		1362: rom = 27;
		1363: rom = 27;
		1364: rom = 27;
		1365: rom = 27;
		1366: rom = 27;
		1367: rom = 27;
		1368: rom = 27;
		1369: rom = 27;
		1370: rom = 27;
		1371: rom = 27;
		1372: rom = 27;
		1373: rom = 27;
		1374: rom = 27;
		1375: rom = 27;
		1376: rom = 27;
		1377: rom = 27;
		1378: rom = 27;
		1379: rom = 27;
		1380: rom = 27;
		1381: rom = 27;
		1382: rom = 27;
		1383: rom = 27;
		1384: rom = 27;
		1385: rom = 27;
		1386: rom = 27;
		1387: rom = 27;
		1388: rom = 27;
		1389: rom = 27;
		1390: rom = 27;
		1391: rom = 27;
		1392: rom = 27;
		1393: rom = 27;
		1394: rom = 27;
		1395: rom = 27;
		1396: rom = 27;
		1397: rom = 27;
		1398: rom = 27;
		1399: rom = 27;
		1400: rom = 27;
		1401: rom = 27;
		1402: rom = 27;
		1408: rom = 27;
		1409: rom = 27;
		1410: rom = 27;
		1411: rom = 27;
		1412: rom = 27;
		1413: rom = 27;
		1414: rom = 27;
		1415: rom = 21;
		1416: rom = 7;
		1417: rom = 22;
		1418: rom = 27;
		1419: rom = 27;
		1420: rom = 27;
		1421: rom = 27;
		1422: rom = 27;
		1423: rom = 27;
		1424: rom = 27;
		1425: rom = 27;
		1426: rom = 27;
		1427: rom = 27;
		1428: rom = 27;
		1429: rom = 27;
		1430: rom = 27;
		1431: rom = 27;
		1432: rom = 27;
		1433: rom = 27;
		1434: rom = 27;
		1435: rom = 27;
		1436: rom = 27;
		1437: rom = 27;
		1438: rom = 27;
		1439: rom = 27;
		1440: rom = 27;
		1441: rom = 27;
		1442: rom = 27;
		1443: rom = 27;
		1444: rom = 27;
		1445: rom = 27;
		1446: rom = 27;
		1447: rom = 27;
		1448: rom = 27;
		1449: rom = 27;
		1450: rom = 27;
		1451: rom = 27;
		1452: rom = 27;
		1453: rom = 27;
		1454: rom = 27;
		1455: rom = 27;
		1456: rom = 27;
		1457: rom = 27;
		1458: rom = 27;
		1459: rom = 27;
		1460: rom = 27;
		1461: rom = 27;
		1462: rom = 27;
		1463: rom = 27;
		1464: rom = 27;
		1465: rom = 27;
		1466: rom = 27;
		1467: rom = 27;
		1468: rom = 27;
		1469: rom = 27;
		1470: rom = 27;
		1471: rom = 27;
		1472: rom = 27;
		1473: rom = 27;
		1474: rom = 27;
		1475: rom = 27;
		1476: rom = 27;
		1477: rom = 27;
		1478: rom = 27;
		1479: rom = 27;
		1480: rom = 27;
		1481: rom = 27;
		1482: rom = 27;
		1483: rom = 27;
		1484: rom = 27;
		1485: rom = 27;
		1486: rom = 27;
		1487: rom = 27;
		1488: rom = 27;
		1489: rom = 27;
		1490: rom = 20;
		1491: rom = 11;
		1492: rom = 11;
		1493: rom = 10;
		1494: rom = 10;
		1495: rom = 10;
		1496: rom = 12;
		1497: rom = 27;
		1498: rom = 27;
		1499: rom = 27;
		1500: rom = 27;
		1501: rom = 27;
		1502: rom = 27;
		1503: rom = 27;
		1504: rom = 27;
		1505: rom = 27;
		1506: rom = 27;
		1507: rom = 27;
		1508: rom = 27;
		1509: rom = 27;
		1510: rom = 27;
		1511: rom = 27;
		1512: rom = 27;
		1513: rom = 27;
		1514: rom = 27;
		1515: rom = 27;
		1516: rom = 27;
		1517: rom = 27;
		1518: rom = 27;
		1519: rom = 27;
		1520: rom = 27;
		1521: rom = 27;
		1522: rom = 27;
		1523: rom = 27;
		1524: rom = 27;
		1525: rom = 27;
		1526: rom = 27;
		1527: rom = 27;
		1528: rom = 27;
		1529: rom = 27;
		1530: rom = 27;
		1536: rom = 27;
		1537: rom = 27;
		1538: rom = 27;
		1539: rom = 27;
		1540: rom = 27;
		1541: rom = 27;
		1542: rom = 27;
		1543: rom = 27;
		1544: rom = 12;
		1545: rom = 13;
		1546: rom = 17;
		1547: rom = 27;
		1548: rom = 27;
		1549: rom = 27;
		1550: rom = 27;
		1551: rom = 27;
		1552: rom = 27;
		1553: rom = 27;
		1554: rom = 27;
		1555: rom = 27;
		1556: rom = 27;
		1557: rom = 27;
		1558: rom = 27;
		1559: rom = 27;
		1560: rom = 27;
		1561: rom = 27;
		1562: rom = 27;
		1563: rom = 27;
		1564: rom = 27;
		1565: rom = 27;
		1566: rom = 27;
		1567: rom = 27;
		1568: rom = 27;
		1569: rom = 27;
		1570: rom = 27;
		1571: rom = 27;
		1572: rom = 27;
		1573: rom = 27;
		1574: rom = 27;
		1575: rom = 27;
		1576: rom = 27;
		1577: rom = 27;
		1578: rom = 27;
		1579: rom = 27;
		1580: rom = 27;
		1581: rom = 27;
		1582: rom = 27;
		1583: rom = 27;
		1584: rom = 27;
		1585: rom = 27;
		1586: rom = 27;
		1587: rom = 27;
		1588: rom = 27;
		1589: rom = 27;
		1590: rom = 27;
		1591: rom = 27;
		1592: rom = 27;
		1593: rom = 27;
		1594: rom = 27;
		1595: rom = 27;
		1596: rom = 27;
		1597: rom = 27;
		1598: rom = 27;
		1599: rom = 27;
		1600: rom = 27;
		1601: rom = 27;
		1602: rom = 27;
		1603: rom = 27;
		1604: rom = 27;
		1605: rom = 27;
		1606: rom = 27;
		1607: rom = 27;
		1608: rom = 27;
		1609: rom = 27;
		1610: rom = 27;
		1611: rom = 27;
		1612: rom = 27;
		1613: rom = 27;
		1614: rom = 27;
		1615: rom = 27;
		1616: rom = 27;
		1617: rom = 27;
		1618: rom = 19;
		1619: rom = 0;
		1620: rom = 0;
		1621: rom = 0;
		1622: rom = 0;
		1623: rom = 0;
		1624: rom = 0;
		1625: rom = 20;
		1626: rom = 27;
		1627: rom = 27;
		1628: rom = 27;
		1629: rom = 27;
		1630: rom = 27;
		1631: rom = 27;
		1632: rom = 27;
		1633: rom = 27;
		1634: rom = 27;
		1635: rom = 27;
		1636: rom = 27;
		1637: rom = 27;
		1638: rom = 27;
		1639: rom = 27;
		1640: rom = 27;
		1641: rom = 27;
		1642: rom = 27;
		1643: rom = 27;
		1644: rom = 27;
		1645: rom = 27;
		1646: rom = 27;
		1647: rom = 27;
		1648: rom = 27;
		1649: rom = 27;
		1650: rom = 27;
		1651: rom = 27;
		1652: rom = 27;
		1653: rom = 27;
		1654: rom = 27;
		1655: rom = 27;
		1656: rom = 27;
		1657: rom = 27;
		1658: rom = 27;
		1664: rom = 27;
		1665: rom = 27;
		1666: rom = 27;
		1667: rom = 27;
		1668: rom = 27;
		1669: rom = 27;
		1670: rom = 27;
		1671: rom = 27;
		1672: rom = 20;
		1673: rom = 15;
		1674: rom = 16;
		1675: rom = 12;
		1676: rom = 23;
		1677: rom = 27;
		1678: rom = 27;
		1679: rom = 27;
		1680: rom = 27;
		1681: rom = 27;
		1682: rom = 27;
		1683: rom = 27;
		1684: rom = 27;
		1685: rom = 27;
		1686: rom = 27;
		1687: rom = 27;
		1688: rom = 27;
		1689: rom = 27;
		1690: rom = 27;
		1691: rom = 27;
		1692: rom = 27;
		1693: rom = 27;
		1694: rom = 27;
		1695: rom = 27;
		1696: rom = 27;
		1697: rom = 27;
		1698: rom = 27;
		1699: rom = 27;
		1700: rom = 27;
		1701: rom = 27;
		1702: rom = 27;
		1703: rom = 27;
		1704: rom = 27;
		1705: rom = 27;
		1706: rom = 27;
		1707: rom = 27;
		1708: rom = 27;
		1709: rom = 20;
		1710: rom = 27;
		1711: rom = 27;
		1712: rom = 27;
		1713: rom = 27;
		1714: rom = 27;
		1715: rom = 27;
		1716: rom = 27;
		1717: rom = 27;
		1718: rom = 27;
		1719: rom = 27;
		1720: rom = 27;
		1721: rom = 27;
		1722: rom = 27;
		1723: rom = 27;
		1724: rom = 27;
		1725: rom = 27;
		1726: rom = 27;
		1727: rom = 27;
		1728: rom = 27;
		1729: rom = 27;
		1730: rom = 27;
		1731: rom = 27;
		1732: rom = 27;
		1733: rom = 27;
		1734: rom = 27;
		1735: rom = 27;
		1736: rom = 27;
		1737: rom = 27;
		1738: rom = 27;
		1739: rom = 27;
		1740: rom = 27;
		1741: rom = 27;
		1742: rom = 27;
		1743: rom = 27;
		1744: rom = 27;
		1745: rom = 27;
		1746: rom = 19;
		1747: rom = 0;
		1748: rom = 0;
		1749: rom = 0;
		1750: rom = 0;
		1751: rom = 14;
		1752: rom = 18;
		1753: rom = 20;
		1754: rom = 27;
		1755: rom = 27;
		1756: rom = 27;
		1757: rom = 27;
		1758: rom = 27;
		1759: rom = 27;
		1760: rom = 27;
		1761: rom = 27;
		1762: rom = 27;
		1763: rom = 27;
		1764: rom = 27;
		1765: rom = 27;
		1766: rom = 27;
		1767: rom = 27;
		1768: rom = 27;
		1769: rom = 27;
		1770: rom = 27;
		1771: rom = 27;
		1772: rom = 27;
		1773: rom = 27;
		1774: rom = 27;
		1775: rom = 27;
		1776: rom = 27;
		1777: rom = 27;
		1778: rom = 27;
		1779: rom = 27;
		1780: rom = 27;
		1781: rom = 27;
		1782: rom = 27;
		1783: rom = 27;
		1784: rom = 27;
		1785: rom = 27;
		1786: rom = 27;
		1792: rom = 27;
		1793: rom = 27;
		1794: rom = 27;
		1795: rom = 27;
		1796: rom = 27;
		1797: rom = 27;
		1798: rom = 27;
		1799: rom = 27;
		1800: rom = 27;
		1801: rom = 12;
		1802: rom = 18;
		1803: rom = 18;
		1804: rom = 13;
		1805: rom = 16;
		1806: rom = 25;
		1807: rom = 27;
		1808: rom = 27;
		1809: rom = 27;
		1810: rom = 27;
		1811: rom = 27;
		1812: rom = 27;
		1813: rom = 27;
		1814: rom = 27;
		1815: rom = 27;
		1816: rom = 27;
		1817: rom = 27;
		1818: rom = 27;
		1819: rom = 27;
		1820: rom = 27;
		1821: rom = 27;
		1822: rom = 27;
		1823: rom = 27;
		1824: rom = 27;
		1825: rom = 27;
		1826: rom = 27;
		1827: rom = 27;
		1828: rom = 27;
		1829: rom = 27;
		1830: rom = 27;
		1831: rom = 27;
		1832: rom = 27;
		1833: rom = 27;
		1834: rom = 27;
		1835: rom = 27;
		1836: rom = 23;
		1837: rom = 15;
		1838: rom = 27;
		1839: rom = 27;
		1840: rom = 27;
		1841: rom = 27;
		1842: rom = 27;
		1843: rom = 27;
		1844: rom = 27;
		1845: rom = 27;
		1846: rom = 27;
		1847: rom = 27;
		1848: rom = 27;
		1849: rom = 27;
		1850: rom = 27;
		1851: rom = 27;
		1852: rom = 27;
		1853: rom = 27;
		1854: rom = 27;
		1855: rom = 27;
		1856: rom = 27;
		1857: rom = 27;
		1858: rom = 27;
		1859: rom = 27;
		1860: rom = 27;
		1861: rom = 27;
		1862: rom = 27;
		1863: rom = 27;
		1864: rom = 27;
		1865: rom = 27;
		1866: rom = 27;
		1867: rom = 27;
		1868: rom = 27;
		1869: rom = 27;
		1870: rom = 27;
		1871: rom = 27;
		1872: rom = 27;
		1873: rom = 27;
		1874: rom = 19;
		1875: rom = 0;
		1876: rom = 0;
		1877: rom = 0;
		1878: rom = 0;
		1879: rom = 8;
		1880: rom = 25;
		1881: rom = 27;
		1882: rom = 24;
		1883: rom = 10;
		1884: rom = 26;
		1885: rom = 27;
		1886: rom = 27;
		1887: rom = 27;
		1888: rom = 27;
		1889: rom = 27;
		1890: rom = 27;
		1891: rom = 27;
		1892: rom = 27;
		1893: rom = 27;
		1894: rom = 27;
		1895: rom = 27;
		1896: rom = 27;
		1897: rom = 27;
		1898: rom = 27;
		1899: rom = 27;
		1900: rom = 27;
		1901: rom = 27;
		1902: rom = 27;
		1903: rom = 27;
		1904: rom = 27;
		1905: rom = 27;
		1906: rom = 27;
		1907: rom = 27;
		1908: rom = 27;
		1909: rom = 27;
		1910: rom = 27;
		1911: rom = 27;
		1912: rom = 27;
		1913: rom = 27;
		1914: rom = 27;
		1920: rom = 27;
		1921: rom = 27;
		1922: rom = 27;
		1923: rom = 27;
		1924: rom = 27;
		1925: rom = 27;
		1926: rom = 27;
		1927: rom = 27;
		1928: rom = 27;
		1929: rom = 21;
		1930: rom = 15;
		1931: rom = 18;
		1932: rom = 18;
		1933: rom = 17;
		1934: rom = 11;
		1935: rom = 17;
		1936: rom = 26;
		1937: rom = 27;
		1938: rom = 27;
		1939: rom = 27;
		1940: rom = 27;
		1941: rom = 27;
		1942: rom = 27;
		1943: rom = 27;
		1944: rom = 27;
		1945: rom = 27;
		1946: rom = 27;
		1947: rom = 27;
		1948: rom = 27;
		1949: rom = 27;
		1950: rom = 27;
		1951: rom = 27;
		1952: rom = 27;
		1953: rom = 27;
		1954: rom = 27;
		1955: rom = 27;
		1956: rom = 27;
		1957: rom = 27;
		1958: rom = 27;
		1959: rom = 27;
		1960: rom = 27;
		1961: rom = 27;
		1962: rom = 27;
		1963: rom = 27;
		1964: rom = 13;
		1965: rom = 15;
		1966: rom = 27;
		1967: rom = 27;
		1968: rom = 27;
		1969: rom = 27;
		1970: rom = 27;
		1971: rom = 27;
		1972: rom = 27;
		1973: rom = 27;
		1974: rom = 27;
		1975: rom = 27;
		1976: rom = 27;
		1977: rom = 27;
		1978: rom = 27;
		1979: rom = 27;
		1980: rom = 27;
		1981: rom = 27;
		1982: rom = 27;
		1983: rom = 27;
		1984: rom = 27;
		1985: rom = 27;
		1986: rom = 27;
		1987: rom = 27;
		1988: rom = 27;
		1989: rom = 27;
		1990: rom = 27;
		1991: rom = 27;
		1992: rom = 27;
		1993: rom = 27;
		1994: rom = 27;
		1995: rom = 27;
		1996: rom = 27;
		1997: rom = 27;
		1998: rom = 27;
		1999: rom = 27;
		2000: rom = 27;
		2001: rom = 27;
		2002: rom = 19;
		2003: rom = 0;
		2004: rom = 0;
		2005: rom = 0;
		2006: rom = 0;
		2007: rom = 0;
		2008: rom = 11;
		2009: rom = 25;
		2010: rom = 9;
		2011: rom = 0;
		2012: rom = 13;
		2013: rom = 27;
		2014: rom = 27;
		2015: rom = 27;
		2016: rom = 27;
		2017: rom = 27;
		2018: rom = 27;
		2019: rom = 27;
		2020: rom = 27;
		2021: rom = 27;
		2022: rom = 27;
		2023: rom = 27;
		2024: rom = 27;
		2025: rom = 27;
		2026: rom = 27;
		2027: rom = 27;
		2028: rom = 27;
		2029: rom = 27;
		2030: rom = 27;
		2031: rom = 27;
		2032: rom = 27;
		2033: rom = 27;
		2034: rom = 27;
		2035: rom = 27;
		2036: rom = 27;
		2037: rom = 27;
		2038: rom = 27;
		2039: rom = 27;
		2040: rom = 27;
		2041: rom = 27;
		2042: rom = 27;
		2048: rom = 27;
		2049: rom = 27;
		2050: rom = 27;
		2051: rom = 27;
		2052: rom = 27;
		2053: rom = 27;
		2054: rom = 27;
		2055: rom = 27;
		2056: rom = 27;
		2057: rom = 27;
		2058: rom = 12;
		2059: rom = 18;
		2060: rom = 18;
		2061: rom = 18;
		2062: rom = 18;
		2063: rom = 17;
		2064: rom = 11;
		2065: rom = 17;
		2066: rom = 26;
		2067: rom = 27;
		2068: rom = 27;
		2069: rom = 27;
		2070: rom = 27;
		2071: rom = 27;
		2072: rom = 27;
		2073: rom = 27;
		2074: rom = 27;
		2075: rom = 27;
		2076: rom = 27;
		2077: rom = 27;
		2078: rom = 27;
		2079: rom = 27;
		2080: rom = 27;
		2081: rom = 27;
		2082: rom = 27;
		2083: rom = 27;
		2084: rom = 27;
		2085: rom = 27;
		2086: rom = 27;
		2087: rom = 27;
		2088: rom = 27;
		2089: rom = 27;
		2090: rom = 27;
		2091: rom = 20;
		2092: rom = 16;
		2093: rom = 15;
		2094: rom = 27;
		2095: rom = 27;
		2096: rom = 27;
		2097: rom = 27;
		2098: rom = 27;
		2099: rom = 27;
		2100: rom = 27;
		2101: rom = 27;
		2102: rom = 27;
		2103: rom = 27;
		2104: rom = 27;
		2105: rom = 27;
		2106: rom = 27;
		2107: rom = 27;
		2108: rom = 27;
		2109: rom = 27;
		2110: rom = 27;
		2111: rom = 27;
		2112: rom = 27;
		2113: rom = 27;
		2114: rom = 27;
		2115: rom = 27;
		2116: rom = 27;
		2117: rom = 27;
		2118: rom = 27;
		2119: rom = 27;
		2120: rom = 27;
		2121: rom = 27;
		2122: rom = 27;
		2123: rom = 27;
		2124: rom = 27;
		2125: rom = 27;
		2126: rom = 27;
		2127: rom = 27;
		2128: rom = 27;
		2129: rom = 27;
		2130: rom = 18;
		2131: rom = 0;
		2132: rom = 7;
		2133: rom = 0;
		2134: rom = 0;
		2135: rom = 0;
		2136: rom = 0;
		2137: rom = 3;
		2138: rom = 0;
		2139: rom = 0;
		2140: rom = 15;
		2141: rom = 27;
		2142: rom = 27;
		2143: rom = 27;
		2144: rom = 27;
		2145: rom = 27;
		2146: rom = 27;
		2147: rom = 27;
		2148: rom = 27;
		2149: rom = 27;
		2150: rom = 27;
		2151: rom = 27;
		2152: rom = 27;
		2153: rom = 27;
		2154: rom = 27;
		2155: rom = 27;
		2156: rom = 27;
		2157: rom = 27;
		2158: rom = 27;
		2159: rom = 27;
		2160: rom = 27;
		2161: rom = 27;
		2162: rom = 27;
		2163: rom = 27;
		2164: rom = 27;
		2165: rom = 27;
		2166: rom = 27;
		2167: rom = 27;
		2168: rom = 27;
		2169: rom = 27;
		2170: rom = 27;
		2176: rom = 27;
		2177: rom = 27;
		2178: rom = 27;
		2179: rom = 27;
		2180: rom = 27;
		2181: rom = 27;
		2182: rom = 27;
		2183: rom = 27;
		2184: rom = 27;
		2185: rom = 27;
		2186: rom = 22;
		2187: rom = 15;
		2188: rom = 18;
		2189: rom = 18;
		2190: rom = 18;
		2191: rom = 18;
		2192: rom = 18;
		2193: rom = 17;
		2194: rom = 11;
		2195: rom = 18;
		2196: rom = 26;
		2197: rom = 27;
		2198: rom = 27;
		2199: rom = 27;
		2200: rom = 27;
		2201: rom = 27;
		2202: rom = 27;
		2203: rom = 27;
		2204: rom = 27;
		2205: rom = 27;
		2206: rom = 27;
		2207: rom = 27;
		2208: rom = 27;
		2209: rom = 27;
		2210: rom = 27;
		2211: rom = 27;
		2212: rom = 27;
		2213: rom = 27;
		2214: rom = 27;
		2215: rom = 27;
		2216: rom = 27;
		2217: rom = 27;
		2218: rom = 25;
		2219: rom = 12;
		2220: rom = 18;
		2221: rom = 15;
		2222: rom = 27;
		2223: rom = 27;
		2224: rom = 27;
		2225: rom = 27;
		2226: rom = 27;
		2227: rom = 27;
		2228: rom = 27;
		2229: rom = 27;
		2230: rom = 27;
		2231: rom = 27;
		2232: rom = 27;
		2233: rom = 27;
		2234: rom = 27;
		2235: rom = 27;
		2236: rom = 27;
		2237: rom = 27;
		2238: rom = 27;
		2239: rom = 27;
		2240: rom = 27;
		2241: rom = 27;
		2242: rom = 27;
		2243: rom = 27;
		2244: rom = 27;
		2245: rom = 27;
		2246: rom = 27;
		2247: rom = 27;
		2248: rom = 27;
		2249: rom = 27;
		2250: rom = 27;
		2251: rom = 27;
		2252: rom = 27;
		2253: rom = 27;
		2254: rom = 27;
		2255: rom = 27;
		2256: rom = 27;
		2257: rom = 27;
		2258: rom = 18;
		2259: rom = 0;
		2260: rom = 19;
		2261: rom = 16;
		2262: rom = 0;
		2263: rom = 0;
		2264: rom = 0;
		2265: rom = 0;
		2266: rom = 0;
		2267: rom = 16;
		2268: rom = 27;
		2269: rom = 27;
		2270: rom = 27;
		2271: rom = 27;
		2272: rom = 26;
		2273: rom = 21;
		2274: rom = 18;
		2275: rom = 17;
		2276: rom = 17;
		2277: rom = 19;
		2278: rom = 24;
		2279: rom = 27;
		2280: rom = 27;
		2281: rom = 27;
		2282: rom = 27;
		2283: rom = 27;
		2284: rom = 27;
		2285: rom = 27;
		2286: rom = 27;
		2287: rom = 27;
		2288: rom = 27;
		2289: rom = 27;
		2290: rom = 27;
		2291: rom = 27;
		2292: rom = 27;
		2293: rom = 27;
		2294: rom = 27;
		2295: rom = 27;
		2296: rom = 27;
		2297: rom = 27;
		2298: rom = 27;
		2304: rom = 27;
		2305: rom = 27;
		2306: rom = 27;
		2307: rom = 27;
		2308: rom = 27;
		2309: rom = 27;
		2310: rom = 27;
		2311: rom = 27;
		2312: rom = 27;
		2313: rom = 27;
		2314: rom = 27;
		2315: rom = 13;
		2316: rom = 18;
		2317: rom = 18;
		2318: rom = 18;
		2319: rom = 18;
		2320: rom = 18;
		2321: rom = 18;
		2322: rom = 18;
		2323: rom = 16;
		2324: rom = 11;
		2325: rom = 20;
		2326: rom = 27;
		2327: rom = 27;
		2328: rom = 27;
		2329: rom = 27;
		2330: rom = 27;
		2331: rom = 27;
		2332: rom = 27;
		2333: rom = 27;
		2334: rom = 27;
		2335: rom = 27;
		2336: rom = 27;
		2337: rom = 27;
		2338: rom = 27;
		2339: rom = 27;
		2340: rom = 27;
		2341: rom = 27;
		2342: rom = 27;
		2343: rom = 27;
		2344: rom = 27;
		2345: rom = 27;
		2346: rom = 15;
		2347: rom = 17;
		2348: rom = 18;
		2349: rom = 15;
		2350: rom = 27;
		2351: rom = 27;
		2352: rom = 27;
		2353: rom = 27;
		2354: rom = 27;
		2355: rom = 27;
		2356: rom = 27;
		2357: rom = 27;
		2358: rom = 27;
		2359: rom = 27;
		2360: rom = 27;
		2361: rom = 27;
		2362: rom = 27;
		2363: rom = 27;
		2364: rom = 27;
		2365: rom = 27;
		2366: rom = 27;
		2367: rom = 27;
		2368: rom = 27;
		2369: rom = 27;
		2370: rom = 27;
		2371: rom = 27;
		2372: rom = 27;
		2373: rom = 27;
		2374: rom = 27;
		2375: rom = 27;
		2376: rom = 27;
		2377: rom = 27;
		2378: rom = 27;
		2379: rom = 27;
		2380: rom = 27;
		2381: rom = 27;
		2382: rom = 27;
		2383: rom = 27;
		2384: rom = 27;
		2385: rom = 27;
		2386: rom = 24;
		2387: rom = 4;
		2388: rom = 19;
		2389: rom = 27;
		2390: rom = 13;
		2391: rom = 0;
		2392: rom = 0;
		2393: rom = 0;
		2394: rom = 0;
		2395: rom = 21;
		2396: rom = 27;
		2397: rom = 27;
		2398: rom = 24;
		2399: rom = 15;
		2400: rom = 2;
		2401: rom = 0;
		2402: rom = 0;
		2403: rom = 0;
		2404: rom = 0;
		2405: rom = 0;
		2406: rom = 0;
		2407: rom = 8;
		2408: rom = 20;
		2409: rom = 27;
		2410: rom = 27;
		2411: rom = 27;
		2412: rom = 27;
		2413: rom = 27;
		2414: rom = 27;
		2415: rom = 27;
		2416: rom = 27;
		2417: rom = 27;
		2418: rom = 27;
		2419: rom = 27;
		2420: rom = 27;
		2421: rom = 27;
		2422: rom = 27;
		2423: rom = 27;
		2424: rom = 27;
		2425: rom = 27;
		2426: rom = 27;
		2432: rom = 27;
		2433: rom = 27;
		2434: rom = 27;
		2435: rom = 27;
		2436: rom = 27;
		2437: rom = 27;
		2438: rom = 27;
		2439: rom = 27;
		2440: rom = 27;
		2441: rom = 27;
		2442: rom = 27;
		2443: rom = 23;
		2444: rom = 14;
		2445: rom = 18;
		2446: rom = 18;
		2447: rom = 18;
		2448: rom = 18;
		2449: rom = 18;
		2450: rom = 18;
		2451: rom = 18;
		2452: rom = 18;
		2453: rom = 15;
		2454: rom = 12;
		2455: rom = 23;
		2456: rom = 27;
		2457: rom = 27;
		2458: rom = 27;
		2459: rom = 27;
		2460: rom = 27;
		2461: rom = 27;
		2462: rom = 27;
		2463: rom = 27;
		2464: rom = 27;
		2465: rom = 27;
		2466: rom = 27;
		2467: rom = 27;
		2468: rom = 27;
		2469: rom = 27;
		2470: rom = 27;
		2471: rom = 27;
		2472: rom = 27;
		2473: rom = 22;
		2474: rom = 14;
		2475: rom = 18;
		2476: rom = 18;
		2477: rom = 15;
		2478: rom = 27;
		2479: rom = 27;
		2480: rom = 27;
		2481: rom = 27;
		2482: rom = 27;
		2483: rom = 27;
		2484: rom = 27;
		2485: rom = 27;
		2486: rom = 27;
		2487: rom = 27;
		2488: rom = 27;
		2489: rom = 27;
		2490: rom = 27;
		2491: rom = 27;
		2492: rom = 27;
		2493: rom = 27;
		2494: rom = 27;
		2495: rom = 27;
		2496: rom = 27;
		2497: rom = 27;
		2498: rom = 27;
		2499: rom = 27;
		2500: rom = 27;
		2501: rom = 27;
		2502: rom = 27;
		2503: rom = 27;
		2504: rom = 27;
		2505: rom = 27;
		2506: rom = 27;
		2507: rom = 27;
		2508: rom = 27;
		2509: rom = 27;
		2510: rom = 27;
		2511: rom = 27;
		2512: rom = 27;
		2513: rom = 27;
		2514: rom = 27;
		2515: rom = 25;
		2516: rom = 23;
		2517: rom = 27;
		2518: rom = 19;
		2519: rom = 0;
		2520: rom = 0;
		2521: rom = 0;
		2522: rom = 0;
		2523: rom = 3;
		2524: rom = 22;
		2525: rom = 18;
		2526: rom = 1;
		2527: rom = 0;
		2528: rom = 0;
		2529: rom = 0;
		2530: rom = 0;
		2531: rom = 0;
		2532: rom = 0;
		2533: rom = 0;
		2534: rom = 0;
		2535: rom = 0;
		2536: rom = 0;
		2537: rom = 9;
		2538: rom = 23;
		2539: rom = 27;
		2540: rom = 27;
		2541: rom = 27;
		2542: rom = 27;
		2543: rom = 27;
		2544: rom = 27;
		2545: rom = 27;
		2546: rom = 27;
		2547: rom = 27;
		2548: rom = 27;
		2549: rom = 27;
		2550: rom = 27;
		2551: rom = 27;
		2552: rom = 27;
		2553: rom = 27;
		2554: rom = 27;
		2560: rom = 27;
		2561: rom = 27;
		2562: rom = 27;
		2563: rom = 27;
		2564: rom = 27;
		2565: rom = 27;
		2566: rom = 27;
		2567: rom = 27;
		2568: rom = 27;
		2569: rom = 27;
		2570: rom = 27;
		2571: rom = 27;
		2572: rom = 14;
		2573: rom = 18;
		2574: rom = 18;
		2575: rom = 18;
		2576: rom = 18;
		2577: rom = 18;
		2578: rom = 18;
		2579: rom = 18;
		2580: rom = 18;
		2581: rom = 18;
		2582: rom = 18;
		2583: rom = 13;
		2584: rom = 16;
		2585: rom = 26;
		2586: rom = 27;
		2587: rom = 27;
		2588: rom = 27;
		2589: rom = 27;
		2590: rom = 27;
		2591: rom = 27;
		2592: rom = 27;
		2593: rom = 27;
		2594: rom = 27;
		2595: rom = 27;
		2596: rom = 27;
		2597: rom = 27;
		2598: rom = 27;
		2599: rom = 27;
		2600: rom = 26;
		2601: rom = 12;
		2602: rom = 18;
		2603: rom = 18;
		2604: rom = 18;
		2605: rom = 16;
		2606: rom = 27;
		2607: rom = 27;
		2608: rom = 27;
		2609: rom = 27;
		2610: rom = 27;
		2611: rom = 27;
		2612: rom = 27;
		2613: rom = 27;
		2614: rom = 27;
		2615: rom = 27;
		2616: rom = 27;
		2617: rom = 27;
		2618: rom = 27;
		2619: rom = 27;
		2620: rom = 27;
		2621: rom = 27;
		2622: rom = 27;
		2623: rom = 27;
		2624: rom = 27;
		2625: rom = 27;
		2626: rom = 27;
		2627: rom = 27;
		2628: rom = 27;
		2629: rom = 27;
		2630: rom = 27;
		2631: rom = 27;
		2632: rom = 27;
		2633: rom = 27;
		2634: rom = 27;
		2635: rom = 27;
		2636: rom = 27;
		2637: rom = 27;
		2638: rom = 27;
		2639: rom = 27;
		2640: rom = 27;
		2641: rom = 27;
		2642: rom = 27;
		2643: rom = 27;
		2644: rom = 27;
		2645: rom = 19;
		2646: rom = 0;
		2647: rom = 0;
		2648: rom = 0;
		2649: rom = 0;
		2650: rom = 0;
		2651: rom = 0;
		2652: rom = 0;
		2653: rom = 0;
		2654: rom = 0;
		2655: rom = 0;
		2656: rom = 0;
		2657: rom = 0;
		2658: rom = 0;
		2659: rom = 0;
		2660: rom = 0;
		2661: rom = 0;
		2662: rom = 0;
		2663: rom = 0;
		2664: rom = 0;
		2665: rom = 0;
		2666: rom = 2;
		2667: rom = 21;
		2668: rom = 27;
		2669: rom = 27;
		2670: rom = 27;
		2671: rom = 27;
		2672: rom = 27;
		2673: rom = 27;
		2674: rom = 27;
		2675: rom = 27;
		2676: rom = 27;
		2677: rom = 27;
		2678: rom = 27;
		2679: rom = 27;
		2680: rom = 27;
		2681: rom = 27;
		2682: rom = 27;
		2688: rom = 27;
		2689: rom = 27;
		2690: rom = 27;
		2691: rom = 27;
		2692: rom = 27;
		2693: rom = 27;
		2694: rom = 27;
		2695: rom = 27;
		2696: rom = 27;
		2697: rom = 27;
		2698: rom = 27;
		2699: rom = 27;
		2700: rom = 24;
		2701: rom = 13;
		2702: rom = 18;
		2703: rom = 18;
		2704: rom = 18;
		2705: rom = 18;
		2706: rom = 19;
		2707: rom = 20;
		2708: rom = 20;
		2709: rom = 20;
		2710: rom = 19;
		2711: rom = 19;
		2712: rom = 17;
		2713: rom = 11;
		2714: rom = 23;
		2715: rom = 27;
		2716: rom = 27;
		2717: rom = 27;
		2718: rom = 27;
		2719: rom = 27;
		2720: rom = 27;
		2721: rom = 27;
		2722: rom = 27;
		2723: rom = 27;
		2724: rom = 27;
		2725: rom = 27;
		2726: rom = 27;
		2727: rom = 27;
		2728: rom = 17;
		2729: rom = 17;
		2730: rom = 18;
		2731: rom = 18;
		2732: rom = 18;
		2733: rom = 12;
		2734: rom = 27;
		2735: rom = 27;
		2736: rom = 27;
		2737: rom = 27;
		2738: rom = 27;
		2739: rom = 27;
		2740: rom = 27;
		2741: rom = 27;
		2742: rom = 27;
		2743: rom = 27;
		2744: rom = 27;
		2745: rom = 27;
		2746: rom = 27;
		2747: rom = 27;
		2748: rom = 27;
		2749: rom = 27;
		2750: rom = 27;
		2751: rom = 27;
		2752: rom = 27;
		2753: rom = 27;
		2754: rom = 27;
		2755: rom = 27;
		2756: rom = 27;
		2757: rom = 27;
		2758: rom = 27;
		2759: rom = 27;
		2760: rom = 27;
		2761: rom = 27;
		2762: rom = 24;
		2763: rom = 25;
		2764: rom = 27;
		2765: rom = 27;
		2766: rom = 27;
		2767: rom = 27;
		2768: rom = 27;
		2769: rom = 27;
		2770: rom = 27;
		2771: rom = 27;
		2772: rom = 26;
		2773: rom = 7;
		2774: rom = 0;
		2775: rom = 3;
		2776: rom = 22;
		2777: rom = 10;
		2778: rom = 0;
		2779: rom = 0;
		2780: rom = 0;
		2781: rom = 0;
		2782: rom = 0;
		2783: rom = 0;
		2784: rom = 2;
		2785: rom = 13;
		2786: rom = 19;
		2787: rom = 20;
		2788: rom = 20;
		2789: rom = 18;
		2790: rom = 9;
		2791: rom = 0;
		2792: rom = 0;
		2793: rom = 0;
		2794: rom = 0;
		2795: rom = 0;
		2796: rom = 21;
		2797: rom = 27;
		2798: rom = 27;
		2799: rom = 27;
		2800: rom = 27;
		2801: rom = 27;
		2802: rom = 27;
		2803: rom = 27;
		2804: rom = 27;
		2805: rom = 27;
		2806: rom = 27;
		2807: rom = 27;
		2808: rom = 27;
		2809: rom = 27;
		2810: rom = 27;
		2816: rom = 27;
		2817: rom = 27;
		2818: rom = 27;
		2819: rom = 27;
		2820: rom = 27;
		2821: rom = 27;
		2822: rom = 27;
		2823: rom = 27;
		2824: rom = 27;
		2825: rom = 27;
		2826: rom = 27;
		2827: rom = 27;
		2828: rom = 27;
		2829: rom = 16;
		2830: rom = 17;
		2831: rom = 18;
		2832: rom = 21;
		2833: rom = 24;
		2834: rom = 25;
		2835: rom = 25;
		2836: rom = 25;
		2837: rom = 25;
		2838: rom = 25;
		2839: rom = 25;
		2840: rom = 24;
		2841: rom = 22;
		2842: rom = 15;
		2843: rom = 19;
		2844: rom = 27;
		2845: rom = 27;
		2846: rom = 27;
		2847: rom = 27;
		2848: rom = 27;
		2849: rom = 27;
		2850: rom = 27;
		2851: rom = 27;
		2852: rom = 27;
		2853: rom = 27;
		2854: rom = 27;
		2855: rom = 24;
		2856: rom = 5;
		2857: rom = 11;
		2858: rom = 18;
		2859: rom = 18;
		2860: rom = 18;
		2861: rom = 11;
		2862: rom = 27;
		2863: rom = 27;
		2864: rom = 27;
		2865: rom = 27;
		2866: rom = 27;
		2867: rom = 27;
		2868: rom = 27;
		2869: rom = 27;
		2870: rom = 27;
		2871: rom = 27;
		2872: rom = 27;
		2873: rom = 27;
		2874: rom = 27;
		2875: rom = 27;
		2876: rom = 27;
		2877: rom = 27;
		2878: rom = 27;
		2879: rom = 27;
		2880: rom = 27;
		2881: rom = 27;
		2882: rom = 27;
		2883: rom = 27;
		2884: rom = 27;
		2885: rom = 27;
		2886: rom = 27;
		2887: rom = 27;
		2888: rom = 27;
		2889: rom = 26;
		2890: rom = 14;
		2891: rom = 15;
		2892: rom = 27;
		2893: rom = 27;
		2894: rom = 27;
		2895: rom = 27;
		2896: rom = 27;
		2897: rom = 27;
		2898: rom = 27;
		2899: rom = 27;
		2900: rom = 27;
		2901: rom = 24;
		2902: rom = 4;
		2903: rom = 20;
		2904: rom = 27;
		2905: rom = 25;
		2906: rom = 5;
		2907: rom = 0;
		2908: rom = 0;
		2909: rom = 0;
		2910: rom = 0;
		2911: rom = 15;
		2912: rom = 25;
		2913: rom = 27;
		2914: rom = 27;
		2915: rom = 27;
		2916: rom = 27;
		2917: rom = 27;
		2918: rom = 27;
		2919: rom = 22;
		2920: rom = 9;
		2921: rom = 0;
		2922: rom = 0;
		2923: rom = 0;
		2924: rom = 3;
		2925: rom = 25;
		2926: rom = 27;
		2927: rom = 27;
		2928: rom = 27;
		2929: rom = 27;
		2930: rom = 27;
		2931: rom = 27;
		2932: rom = 27;
		2933: rom = 27;
		2934: rom = 27;
		2935: rom = 27;
		2936: rom = 27;
		2937: rom = 27;
		2938: rom = 27;
		2944: rom = 27;
		2945: rom = 27;
		2946: rom = 27;
		2947: rom = 27;
		2948: rom = 27;
		2949: rom = 27;
		2950: rom = 27;
		2951: rom = 27;
		2952: rom = 27;
		2953: rom = 27;
		2954: rom = 27;
		2955: rom = 27;
		2956: rom = 27;
		2957: rom = 25;
		2958: rom = 12;
		2959: rom = 21;
		2960: rom = 25;
		2961: rom = 25;
		2962: rom = 25;
		2963: rom = 24;
		2964: rom = 23;
		2965: rom = 23;
		2966: rom = 24;
		2967: rom = 25;
		2968: rom = 25;
		2969: rom = 25;
		2970: rom = 25;
		2971: rom = 21;
		2972: rom = 15;
		2973: rom = 26;
		2974: rom = 27;
		2975: rom = 27;
		2976: rom = 27;
		2977: rom = 27;
		2978: rom = 27;
		2979: rom = 27;
		2980: rom = 27;
		2981: rom = 27;
		2982: rom = 27;
		2983: rom = 13;
		2984: rom = 17;
		2985: rom = 13;
		2986: rom = 17;
		2987: rom = 18;
		2988: rom = 18;
		2989: rom = 13;
		2990: rom = 26;
		2991: rom = 27;
		2992: rom = 27;
		2993: rom = 27;
		2994: rom = 27;
		2995: rom = 27;
		2996: rom = 27;
		2997: rom = 27;
		2998: rom = 27;
		2999: rom = 27;
		3000: rom = 27;
		3001: rom = 27;
		3002: rom = 27;
		3003: rom = 27;
		3004: rom = 27;
		3005: rom = 27;
		3006: rom = 27;
		3007: rom = 27;
		3008: rom = 27;
		3009: rom = 27;
		3010: rom = 27;
		3011: rom = 27;
		3012: rom = 27;
		3013: rom = 27;
		3014: rom = 27;
		3015: rom = 27;
		3016: rom = 27;
		3017: rom = 21;
		3018: rom = 21;
		3019: rom = 15;
		3020: rom = 26;
		3021: rom = 27;
		3022: rom = 27;
		3023: rom = 27;
		3024: rom = 27;
		3025: rom = 27;
		3026: rom = 27;
		3027: rom = 27;
		3028: rom = 27;
		3029: rom = 27;
		3030: rom = 24;
		3031: rom = 27;
		3032: rom = 27;
		3033: rom = 24;
		3034: rom = 1;
		3035: rom = 0;
		3036: rom = 0;
		3037: rom = 0;
		3038: rom = 20;
		3039: rom = 27;
		3040: rom = 27;
		3041: rom = 27;
		3042: rom = 27;
		3043: rom = 27;
		3044: rom = 27;
		3045: rom = 27;
		3046: rom = 27;
		3047: rom = 27;
		3048: rom = 26;
		3049: rom = 14;
		3050: rom = 0;
		3051: rom = 0;
		3052: rom = 0;
		3053: rom = 13;
		3054: rom = 27;
		3055: rom = 27;
		3056: rom = 27;
		3057: rom = 27;
		3058: rom = 27;
		3059: rom = 27;
		3060: rom = 27;
		3061: rom = 27;
		3062: rom = 27;
		3063: rom = 27;
		3064: rom = 27;
		3065: rom = 27;
		3066: rom = 27;
		3072: rom = 27;
		3073: rom = 27;
		3074: rom = 27;
		3075: rom = 27;
		3076: rom = 27;
		3077: rom = 27;
		3078: rom = 27;
		3079: rom = 27;
		3080: rom = 27;
		3081: rom = 27;
		3082: rom = 27;
		3083: rom = 27;
		3084: rom = 27;
		3085: rom = 27;
		3086: rom = 18;
		3087: rom = 22;
		3088: rom = 25;
		3089: rom = 21;
		3090: rom = 18;
		3091: rom = 18;
		3092: rom = 18;
		3093: rom = 18;
		3094: rom = 18;
		3095: rom = 18;
		3096: rom = 20;
		3097: rom = 22;
		3098: rom = 24;
		3099: rom = 25;
		3100: rom = 23;
		3101: rom = 14;
		3102: rom = 26;
		3103: rom = 27;
		3104: rom = 27;
		3105: rom = 27;
		3106: rom = 27;
		3107: rom = 27;
		3108: rom = 27;
		3109: rom = 27;
		3110: rom = 20;
		3111: rom = 15;
		3112: rom = 18;
		3113: rom = 11;
		3114: rom = 12;
		3115: rom = 11;
		3116: rom = 18;
		3117: rom = 15;
		3118: rom = 24;
		3119: rom = 27;
		3120: rom = 27;
		3121: rom = 27;
		3122: rom = 27;
		3123: rom = 27;
		3124: rom = 27;
		3125: rom = 27;
		3126: rom = 27;
		3127: rom = 27;
		3128: rom = 27;
		3129: rom = 27;
		3130: rom = 27;
		3131: rom = 27;
		3132: rom = 27;
		3133: rom = 27;
		3134: rom = 27;
		3135: rom = 27;
		3136: rom = 27;
		3137: rom = 27;
		3138: rom = 27;
		3139: rom = 27;
		3140: rom = 27;
		3141: rom = 27;
		3142: rom = 27;
		3143: rom = 27;
		3144: rom = 27;
		3145: rom = 16;
		3146: rom = 24;
		3147: rom = 19;
		3148: rom = 24;
		3149: rom = 27;
		3150: rom = 27;
		3151: rom = 27;
		3152: rom = 27;
		3153: rom = 27;
		3154: rom = 27;
		3155: rom = 27;
		3156: rom = 27;
		3157: rom = 27;
		3158: rom = 27;
		3159: rom = 27;
		3160: rom = 27;
		3161: rom = 15;
		3162: rom = 0;
		3163: rom = 0;
		3164: rom = 0;
		3165: rom = 19;
		3166: rom = 27;
		3167: rom = 27;
		3168: rom = 27;
		3169: rom = 27;
		3170: rom = 27;
		3171: rom = 27;
		3172: rom = 27;
		3173: rom = 27;
		3174: rom = 27;
		3175: rom = 27;
		3176: rom = 27;
		3177: rom = 27;
		3178: rom = 12;
		3179: rom = 0;
		3180: rom = 0;
		3181: rom = 0;
		3182: rom = 23;
		3183: rom = 27;
		3184: rom = 27;
		3185: rom = 27;
		3186: rom = 27;
		3187: rom = 23;
		3188: rom = 22;
		3189: rom = 22;
		3190: rom = 25;
		3191: rom = 27;
		3192: rom = 27;
		3193: rom = 27;
		3194: rom = 27;
		3200: rom = 27;
		3201: rom = 27;
		3202: rom = 27;
		3203: rom = 27;
		3204: rom = 27;
		3205: rom = 27;
		3206: rom = 27;
		3207: rom = 27;
		3208: rom = 27;
		3209: rom = 27;
		3210: rom = 27;
		3211: rom = 27;
		3212: rom = 27;
		3213: rom = 27;
		3214: rom = 26;
		3215: rom = 15;
		3216: rom = 25;
		3217: rom = 18;
		3218: rom = 18;
		3219: rom = 18;
		3220: rom = 18;
		3221: rom = 18;
		3222: rom = 18;
		3223: rom = 18;
		3224: rom = 18;
		3225: rom = 18;
		3226: rom = 18;
		3227: rom = 20;
		3228: rom = 23;
		3229: rom = 23;
		3230: rom = 14;
		3231: rom = 26;
		3232: rom = 27;
		3233: rom = 27;
		3234: rom = 27;
		3235: rom = 27;
		3236: rom = 27;
		3237: rom = 26;
		3238: rom = 11;
		3239: rom = 18;
		3240: rom = 17;
		3241: rom = 14;
		3242: rom = 14;
		3243: rom = 19;
		3244: rom = 14;
		3245: rom = 16;
		3246: rom = 20;
		3247: rom = 27;
		3248: rom = 27;
		3249: rom = 27;
		3250: rom = 27;
		3251: rom = 27;
		3252: rom = 27;
		3253: rom = 27;
		3254: rom = 27;
		3255: rom = 27;
		3256: rom = 27;
		3257: rom = 27;
		3258: rom = 27;
		3259: rom = 27;
		3260: rom = 27;
		3261: rom = 27;
		3262: rom = 27;
		3263: rom = 27;
		3264: rom = 27;
		3265: rom = 27;
		3266: rom = 27;
		3267: rom = 18;
		3268: rom = 18;
		3269: rom = 27;
		3270: rom = 27;
		3271: rom = 27;
		3272: rom = 27;
		3273: rom = 15;
		3274: rom = 24;
		3275: rom = 21;
		3276: rom = 21;
		3277: rom = 27;
		3278: rom = 27;
		3279: rom = 27;
		3280: rom = 27;
		3281: rom = 27;
		3282: rom = 27;
		3283: rom = 27;
		3284: rom = 27;
		3285: rom = 27;
		3286: rom = 27;
		3287: rom = 27;
		3288: rom = 25;
		3289: rom = 1;
		3290: rom = 0;
		3291: rom = 0;
		3292: rom = 13;
		3293: rom = 27;
		3294: rom = 27;
		3295: rom = 27;
		3296: rom = 27;
		3297: rom = 27;
		3298: rom = 27;
		3299: rom = 27;
		3300: rom = 27;
		3301: rom = 27;
		3302: rom = 27;
		3303: rom = 27;
		3304: rom = 27;
		3305: rom = 27;
		3306: rom = 25;
		3307: rom = 4;
		3308: rom = 0;
		3309: rom = 0;
		3310: rom = 14;
		3311: rom = 27;
		3312: rom = 27;
		3313: rom = 27;
		3314: rom = 27;
		3315: rom = 11;
		3316: rom = 0;
		3317: rom = 0;
		3318: rom = 19;
		3319: rom = 27;
		3320: rom = 27;
		3321: rom = 27;
		3322: rom = 27;
		3328: rom = 27;
		3329: rom = 27;
		3330: rom = 27;
		3331: rom = 27;
		3332: rom = 27;
		3333: rom = 27;
		3334: rom = 27;
		3335: rom = 27;
		3336: rom = 27;
		3337: rom = 27;
		3338: rom = 27;
		3339: rom = 27;
		3340: rom = 27;
		3341: rom = 27;
		3342: rom = 27;
		3343: rom = 21;
		3344: rom = 21;
		3345: rom = 19;
		3346: rom = 18;
		3347: rom = 18;
		3348: rom = 18;
		3349: rom = 18;
		3350: rom = 18;
		3351: rom = 18;
		3352: rom = 18;
		3353: rom = 18;
		3354: rom = 18;
		3355: rom = 18;
		3356: rom = 18;
		3357: rom = 19;
		3358: rom = 21;
		3359: rom = 14;
		3360: rom = 26;
		3361: rom = 27;
		3362: rom = 27;
		3363: rom = 27;
		3364: rom = 27;
		3365: rom = 17;
		3366: rom = 16;
		3367: rom = 18;
		3368: rom = 14;
		3369: rom = 20;
		3370: rom = 22;
		3371: rom = 21;
		3372: rom = 14;
		3373: rom = 18;
		3374: rom = 18;
		3375: rom = 27;
		3376: rom = 27;
		3377: rom = 27;
		3378: rom = 27;
		3379: rom = 27;
		3380: rom = 27;
		3381: rom = 27;
		3382: rom = 27;
		3383: rom = 27;
		3384: rom = 27;
		3385: rom = 27;
		3386: rom = 27;
		3387: rom = 27;
		3388: rom = 27;
		3389: rom = 27;
		3390: rom = 27;
		3391: rom = 27;
		3392: rom = 27;
		3393: rom = 27;
		3394: rom = 27;
		3395: rom = 15;
		3396: rom = 15;
		3397: rom = 27;
		3398: rom = 27;
		3399: rom = 27;
		3400: rom = 23;
		3401: rom = 19;
		3402: rom = 24;
		3403: rom = 23;
		3404: rom = 19;
		3405: rom = 27;
		3406: rom = 27;
		3407: rom = 27;
		3408: rom = 27;
		3409: rom = 27;
		3410: rom = 27;
		3411: rom = 27;
		3412: rom = 27;
		3413: rom = 27;
		3414: rom = 27;
		3415: rom = 27;
		3416: rom = 20;
		3417: rom = 0;
		3418: rom = 0;
		3419: rom = 0;
		3420: rom = 24;
		3421: rom = 27;
		3422: rom = 27;
		3423: rom = 27;
		3424: rom = 27;
		3425: rom = 27;
		3426: rom = 27;
		3427: rom = 27;
		3428: rom = 27;
		3429: rom = 27;
		3430: rom = 27;
		3431: rom = 27;
		3432: rom = 27;
		3433: rom = 27;
		3434: rom = 27;
		3435: rom = 18;
		3436: rom = 0;
		3437: rom = 0;
		3438: rom = 1;
		3439: rom = 26;
		3440: rom = 27;
		3441: rom = 27;
		3442: rom = 27;
		3443: rom = 11;
		3444: rom = 0;
		3445: rom = 0;
		3446: rom = 19;
		3447: rom = 27;
		3448: rom = 27;
		3449: rom = 27;
		3450: rom = 27;
		3456: rom = 27;
		3457: rom = 27;
		3458: rom = 27;
		3459: rom = 27;
		3460: rom = 27;
		3461: rom = 27;
		3462: rom = 27;
		3463: rom = 27;
		3464: rom = 27;
		3465: rom = 27;
		3466: rom = 27;
		3467: rom = 27;
		3468: rom = 27;
		3469: rom = 27;
		3470: rom = 27;
		3471: rom = 27;
		3472: rom = 15;
		3473: rom = 21;
		3474: rom = 18;
		3475: rom = 18;
		3476: rom = 18;
		3477: rom = 18;
		3478: rom = 18;
		3479: rom = 18;
		3480: rom = 18;
		3481: rom = 18;
		3482: rom = 18;
		3483: rom = 18;
		3484: rom = 18;
		3485: rom = 18;
		3486: rom = 18;
		3487: rom = 18;
		3488: rom = 13;
		3489: rom = 26;
		3490: rom = 27;
		3491: rom = 27;
		3492: rom = 25;
		3493: rom = 12;
		3494: rom = 18;
		3495: rom = 18;
		3496: rom = 12;
		3497: rom = 23;
		3498: rom = 24;
		3499: rom = 17;
		3500: rom = 17;
		3501: rom = 18;
		3502: rom = 15;
		3503: rom = 27;
		3504: rom = 27;
		3505: rom = 27;
		3506: rom = 27;
		3507: rom = 27;
		3508: rom = 27;
		3509: rom = 27;
		3510: rom = 27;
		3511: rom = 27;
		3512: rom = 27;
		3513: rom = 27;
		3514: rom = 27;
		3515: rom = 27;
		3516: rom = 27;
		3517: rom = 27;
		3518: rom = 27;
		3519: rom = 27;
		3520: rom = 27;
		3521: rom = 27;
		3522: rom = 24;
		3523: rom = 19;
		3524: rom = 19;
		3525: rom = 23;
		3526: rom = 27;
		3527: rom = 27;
		3528: rom = 19;
		3529: rom = 22;
		3530: rom = 24;
		3531: rom = 24;
		3532: rom = 15;
		3533: rom = 27;
		3534: rom = 27;
		3535: rom = 27;
		3536: rom = 27;
		3537: rom = 27;
		3538: rom = 27;
		3539: rom = 27;
		3540: rom = 27;
		3541: rom = 27;
		3542: rom = 27;
		3543: rom = 27;
		3544: rom = 13;
		3545: rom = 0;
		3546: rom = 0;
		3547: rom = 13;
		3548: rom = 27;
		3549: rom = 27;
		3550: rom = 27;
		3551: rom = 27;
		3552: rom = 27;
		3553: rom = 27;
		3554: rom = 27;
		3555: rom = 27;
		3556: rom = 27;
		3557: rom = 27;
		3558: rom = 27;
		3559: rom = 27;
		3560: rom = 27;
		3561: rom = 27;
		3562: rom = 27;
		3563: rom = 25;
		3564: rom = 0;
		3565: rom = 0;
		3566: rom = 0;
		3567: rom = 22;
		3568: rom = 27;
		3569: rom = 27;
		3570: rom = 27;
		3571: rom = 11;
		3572: rom = 0;
		3573: rom = 0;
		3574: rom = 19;
		3575: rom = 27;
		3576: rom = 27;
		3577: rom = 27;
		3578: rom = 27;
		3584: rom = 27;
		3585: rom = 27;
		3586: rom = 27;
		3587: rom = 27;
		3588: rom = 27;
		3589: rom = 27;
		3590: rom = 27;
		3591: rom = 27;
		3592: rom = 27;
		3593: rom = 27;
		3594: rom = 27;
		3595: rom = 27;
		3596: rom = 27;
		3597: rom = 27;
		3598: rom = 27;
		3599: rom = 27;
		3600: rom = 24;
		3601: rom = 16;
		3602: rom = 18;
		3603: rom = 18;
		3604: rom = 18;
		3605: rom = 18;
		3606: rom = 18;
		3607: rom = 18;
		3608: rom = 18;
		3609: rom = 18;
		3610: rom = 18;
		3611: rom = 18;
		3612: rom = 18;
		3613: rom = 18;
		3614: rom = 18;
		3615: rom = 18;
		3616: rom = 16;
		3617: rom = 14;
		3618: rom = 27;
		3619: rom = 27;
		3620: rom = 15;
		3621: rom = 17;
		3622: rom = 18;
		3623: rom = 17;
		3624: rom = 10;
		3625: rom = 10;
		3626: rom = 22;
		3627: rom = 13;
		3628: rom = 18;
		3629: rom = 18;
		3630: rom = 11;
		3631: rom = 27;
		3632: rom = 27;
		3633: rom = 27;
		3634: rom = 27;
		3635: rom = 27;
		3636: rom = 27;
		3637: rom = 27;
		3638: rom = 27;
		3639: rom = 27;
		3640: rom = 27;
		3641: rom = 27;
		3642: rom = 27;
		3643: rom = 27;
		3644: rom = 27;
		3645: rom = 27;
		3646: rom = 27;
		3647: rom = 27;
		3648: rom = 27;
		3649: rom = 27;
		3650: rom = 20;
		3651: rom = 21;
		3652: rom = 22;
		3653: rom = 20;
		3654: rom = 27;
		3655: rom = 27;
		3656: rom = 16;
		3657: rom = 24;
		3658: rom = 24;
		3659: rom = 24;
		3660: rom = 17;
		3661: rom = 27;
		3662: rom = 27;
		3663: rom = 27;
		3664: rom = 27;
		3665: rom = 27;
		3666: rom = 27;
		3667: rom = 27;
		3668: rom = 27;
		3669: rom = 27;
		3670: rom = 27;
		3671: rom = 27;
		3672: rom = 3;
		3673: rom = 0;
		3674: rom = 0;
		3675: rom = 20;
		3676: rom = 27;
		3677: rom = 27;
		3678: rom = 27;
		3679: rom = 27;
		3680: rom = 27;
		3681: rom = 27;
		3682: rom = 27;
		3683: rom = 27;
		3684: rom = 27;
		3685: rom = 27;
		3686: rom = 27;
		3687: rom = 27;
		3688: rom = 27;
		3689: rom = 27;
		3690: rom = 27;
		3691: rom = 27;
		3692: rom = 12;
		3693: rom = 0;
		3694: rom = 0;
		3695: rom = 18;
		3696: rom = 27;
		3697: rom = 27;
		3698: rom = 27;
		3699: rom = 11;
		3700: rom = 0;
		3701: rom = 0;
		3702: rom = 19;
		3703: rom = 27;
		3704: rom = 27;
		3705: rom = 27;
		3706: rom = 27;
		3712: rom = 27;
		3713: rom = 27;
		3714: rom = 27;
		3715: rom = 27;
		3716: rom = 27;
		3717: rom = 27;
		3718: rom = 27;
		3719: rom = 27;
		3720: rom = 27;
		3721: rom = 27;
		3722: rom = 27;
		3723: rom = 27;
		3724: rom = 27;
		3725: rom = 27;
		3726: rom = 27;
		3727: rom = 27;
		3728: rom = 27;
		3729: rom = 17;
		3730: rom = 17;
		3731: rom = 18;
		3732: rom = 18;
		3733: rom = 18;
		3734: rom = 18;
		3735: rom = 18;
		3736: rom = 18;
		3737: rom = 18;
		3738: rom = 18;
		3739: rom = 18;
		3740: rom = 18;
		3741: rom = 18;
		3742: rom = 18;
		3743: rom = 18;
		3744: rom = 18;
		3745: rom = 15;
		3746: rom = 18;
		3747: rom = 24;
		3748: rom = 13;
		3749: rom = 18;
		3750: rom = 18;
		3751: rom = 18;
		3752: rom = 18;
		3753: rom = 16;
		3754: rom = 17;
		3755: rom = 16;
		3756: rom = 17;
		3757: rom = 18;
		3758: rom = 12;
		3759: rom = 27;
		3760: rom = 27;
		3761: rom = 27;
		3762: rom = 27;
		3763: rom = 27;
		3764: rom = 27;
		3765: rom = 27;
		3766: rom = 27;
		3767: rom = 27;
		3768: rom = 27;
		3769: rom = 27;
		3770: rom = 27;
		3771: rom = 27;
		3772: rom = 27;
		3773: rom = 27;
		3774: rom = 27;
		3775: rom = 27;
		3776: rom = 27;
		3777: rom = 27;
		3778: rom = 16;
		3779: rom = 24;
		3780: rom = 24;
		3781: rom = 16;
		3782: rom = 27;
		3783: rom = 27;
		3784: rom = 15;
		3785: rom = 24;
		3786: rom = 24;
		3787: rom = 24;
		3788: rom = 14;
		3789: rom = 27;
		3790: rom = 27;
		3791: rom = 27;
		3792: rom = 27;
		3793: rom = 27;
		3794: rom = 27;
		3795: rom = 27;
		3796: rom = 27;
		3797: rom = 27;
		3798: rom = 27;
		3799: rom = 25;
		3800: rom = 0;
		3801: rom = 0;
		3802: rom = 0;
		3803: rom = 23;
		3804: rom = 27;
		3805: rom = 27;
		3806: rom = 27;
		3807: rom = 27;
		3808: rom = 27;
		3809: rom = 27;
		3810: rom = 27;
		3811: rom = 27;
		3812: rom = 27;
		3813: rom = 27;
		3814: rom = 27;
		3815: rom = 27;
		3816: rom = 27;
		3817: rom = 27;
		3818: rom = 27;
		3819: rom = 27;
		3820: rom = 17;
		3821: rom = 0;
		3822: rom = 0;
		3823: rom = 7;
		3824: rom = 14;
		3825: rom = 14;
		3826: rom = 14;
		3827: rom = 5;
		3828: rom = 0;
		3829: rom = 0;
		3830: rom = 11;
		3831: rom = 16;
		3832: rom = 16;
		3833: rom = 16;
		3834: rom = 21;
		3840: rom = 27;
		3841: rom = 27;
		3842: rom = 27;
		3843: rom = 27;
		3844: rom = 27;
		3845: rom = 27;
		3846: rom = 27;
		3847: rom = 27;
		3848: rom = 27;
		3849: rom = 27;
		3850: rom = 27;
		3851: rom = 27;
		3852: rom = 27;
		3853: rom = 27;
		3854: rom = 27;
		3855: rom = 27;
		3856: rom = 27;
		3857: rom = 25;
		3858: rom = 11;
		3859: rom = 18;
		3860: rom = 18;
		3861: rom = 18;
		3862: rom = 18;
		3863: rom = 18;
		3864: rom = 15;
		3865: rom = 11;
		3866: rom = 11;
		3867: rom = 11;
		3868: rom = 11;
		3869: rom = 17;
		3870: rom = 18;
		3871: rom = 18;
		3872: rom = 18;
		3873: rom = 18;
		3874: rom = 13;
		3875: rom = 11;
		3876: rom = 17;
		3877: rom = 18;
		3878: rom = 18;
		3879: rom = 18;
		3880: rom = 18;
		3881: rom = 16;
		3882: rom = 18;
		3883: rom = 14;
		3884: rom = 18;
		3885: rom = 18;
		3886: rom = 13;
		3887: rom = 27;
		3888: rom = 27;
		3889: rom = 27;
		3890: rom = 27;
		3891: rom = 27;
		3892: rom = 27;
		3893: rom = 27;
		3894: rom = 27;
		3895: rom = 27;
		3896: rom = 27;
		3897: rom = 27;
		3898: rom = 27;
		3899: rom = 27;
		3900: rom = 27;
		3901: rom = 27;
		3902: rom = 27;
		3903: rom = 27;
		3904: rom = 27;
		3905: rom = 27;
		3906: rom = 17;
		3907: rom = 24;
		3908: rom = 24;
		3909: rom = 15;
		3910: rom = 27;
		3911: rom = 25;
		3912: rom = 17;
		3913: rom = 24;
		3914: rom = 24;
		3915: rom = 24;
		3916: rom = 13;
		3917: rom = 27;
		3918: rom = 27;
		3919: rom = 27;
		3920: rom = 27;
		3921: rom = 27;
		3922: rom = 27;
		3923: rom = 27;
		3924: rom = 27;
		3925: rom = 27;
		3926: rom = 27;
		3927: rom = 24;
		3928: rom = 0;
		3929: rom = 0;
		3930: rom = 0;
		3931: rom = 25;
		3932: rom = 27;
		3933: rom = 27;
		3934: rom = 27;
		3935: rom = 27;
		3936: rom = 27;
		3937: rom = 27;
		3938: rom = 27;
		3939: rom = 27;
		3940: rom = 27;
		3941: rom = 27;
		3942: rom = 27;
		3943: rom = 27;
		3944: rom = 27;
		3945: rom = 27;
		3946: rom = 27;
		3947: rom = 27;
		3948: rom = 20;
		3949: rom = 0;
		3950: rom = 0;
		3951: rom = 0;
		3952: rom = 0;
		3953: rom = 0;
		3954: rom = 0;
		3955: rom = 0;
		3956: rom = 0;
		3957: rom = 0;
		3958: rom = 0;
		3959: rom = 0;
		3960: rom = 0;
		3961: rom = 0;
		3962: rom = 17;
		3968: rom = 27;
		3969: rom = 27;
		3970: rom = 27;
		3971: rom = 27;
		3972: rom = 27;
		3973: rom = 27;
		3974: rom = 27;
		3975: rom = 27;
		3976: rom = 27;
		3977: rom = 27;
		3978: rom = 27;
		3979: rom = 27;
		3980: rom = 27;
		3981: rom = 27;
		3982: rom = 27;
		3983: rom = 27;
		3984: rom = 27;
		3985: rom = 27;
		3986: rom = 19;
		3987: rom = 15;
		3988: rom = 18;
		3989: rom = 18;
		3990: rom = 17;
		3991: rom = 12;
		3992: rom = 15;
		3993: rom = 22;
		3994: rom = 24;
		3995: rom = 24;
		3996: rom = 21;
		3997: rom = 11;
		3998: rom = 11;
		3999: rom = 10;
		4000: rom = 10;
		4001: rom = 10;
		4002: rom = 15;
		4003: rom = 10;
		4004: rom = 17;
		4005: rom = 18;
		4006: rom = 18;
		4007: rom = 18;
		4008: rom = 18;
		4009: rom = 11;
		4010: rom = 20;
		4011: rom = 9;
		4012: rom = 18;
		4013: rom = 18;
		4014: rom = 12;
		4015: rom = 27;
		4016: rom = 27;
		4017: rom = 27;
		4018: rom = 27;
		4019: rom = 27;
		4020: rom = 27;
		4021: rom = 27;
		4022: rom = 27;
		4023: rom = 27;
		4024: rom = 27;
		4025: rom = 27;
		4026: rom = 27;
		4027: rom = 27;
		4028: rom = 27;
		4029: rom = 27;
		4030: rom = 27;
		4031: rom = 27;
		4032: rom = 27;
		4033: rom = 27;
		4034: rom = 13;
		4035: rom = 24;
		4036: rom = 24;
		4037: rom = 15;
		4038: rom = 27;
		4039: rom = 23;
		4040: rom = 20;
		4041: rom = 24;
		4042: rom = 24;
		4043: rom = 24;
		4044: rom = 15;
		4045: rom = 27;
		4046: rom = 27;
		4047: rom = 27;
		4048: rom = 27;
		4049: rom = 19;
		4050: rom = 22;
		4051: rom = 27;
		4052: rom = 27;
		4053: rom = 27;
		4054: rom = 27;
		4055: rom = 24;
		4056: rom = 0;
		4057: rom = 0;
		4058: rom = 0;
		4059: rom = 26;
		4060: rom = 27;
		4061: rom = 27;
		4062: rom = 27;
		4063: rom = 27;
		4064: rom = 27;
		4065: rom = 27;
		4066: rom = 27;
		4067: rom = 27;
		4068: rom = 27;
		4069: rom = 27;
		4070: rom = 27;
		4071: rom = 27;
		4072: rom = 27;
		4073: rom = 27;
		4074: rom = 27;
		4075: rom = 27;
		4076: rom = 20;
		4077: rom = 0;
		4078: rom = 0;
		4079: rom = 0;
		4080: rom = 0;
		4081: rom = 0;
		4082: rom = 0;
		4083: rom = 0;
		4084: rom = 0;
		4085: rom = 0;
		4086: rom = 0;
		4087: rom = 0;
		4088: rom = 0;
		4089: rom = 0;
		4090: rom = 17;
		4096: rom = 27;
		4097: rom = 27;
		4098: rom = 27;
		4099: rom = 27;
		4100: rom = 27;
		4101: rom = 27;
		4102: rom = 27;
		4103: rom = 27;
		4104: rom = 27;
		4105: rom = 27;
		4106: rom = 27;
		4107: rom = 27;
		4108: rom = 27;
		4109: rom = 27;
		4110: rom = 27;
		4111: rom = 27;
		4112: rom = 27;
		4113: rom = 27;
		4114: rom = 27;
		4115: rom = 12;
		4116: rom = 18;
		4117: rom = 18;
		4118: rom = 12;
		4119: rom = 19;
		4120: rom = 24;
		4121: rom = 24;
		4122: rom = 24;
		4123: rom = 24;
		4124: rom = 24;
		4125: rom = 22;
		4126: rom = 14;
		4127: rom = 24;
		4128: rom = 24;
		4129: rom = 23;
		4130: rom = 16;
		4131: rom = 10;
		4132: rom = 11;
		4133: rom = 18;
		4134: rom = 18;
		4135: rom = 18;
		4136: rom = 14;
		4137: rom = 17;
		4138: rom = 24;
		4139: rom = 18;
		4140: rom = 16;
		4141: rom = 18;
		4142: rom = 11;
		4143: rom = 27;
		4144: rom = 27;
		4145: rom = 27;
		4146: rom = 27;
		4147: rom = 27;
		4148: rom = 27;
		4149: rom = 27;
		4150: rom = 27;
		4151: rom = 27;
		4152: rom = 27;
		4153: rom = 27;
		4154: rom = 27;
		4155: rom = 27;
		4156: rom = 25;
		4157: rom = 10;
		4158: rom = 23;
		4159: rom = 27;
		4160: rom = 27;
		4161: rom = 27;
		4162: rom = 16;
		4163: rom = 24;
		4164: rom = 24;
		4165: rom = 18;
		4166: rom = 25;
		4167: rom = 19;
		4168: rom = 22;
		4169: rom = 24;
		4170: rom = 24;
		4171: rom = 24;
		4172: rom = 17;
		4173: rom = 27;
		4174: rom = 27;
		4175: rom = 27;
		4176: rom = 23;
		4177: rom = 17;
		4178: rom = 17;
		4179: rom = 27;
		4180: rom = 27;
		4181: rom = 27;
		4182: rom = 27;
		4183: rom = 24;
		4184: rom = 0;
		4185: rom = 0;
		4186: rom = 0;
		4187: rom = 25;
		4188: rom = 27;
		4189: rom = 27;
		4190: rom = 27;
		4191: rom = 27;
		4192: rom = 27;
		4193: rom = 27;
		4194: rom = 27;
		4195: rom = 27;
		4196: rom = 27;
		4197: rom = 27;
		4198: rom = 27;
		4199: rom = 27;
		4200: rom = 27;
		4201: rom = 27;
		4202: rom = 27;
		4203: rom = 27;
		4204: rom = 20;
		4205: rom = 0;
		4206: rom = 0;
		4207: rom = 0;
		4208: rom = 0;
		4209: rom = 0;
		4210: rom = 0;
		4211: rom = 0;
		4212: rom = 0;
		4213: rom = 0;
		4214: rom = 0;
		4215: rom = 0;
		4216: rom = 0;
		4217: rom = 0;
		4218: rom = 17;
		4224: rom = 27;
		4225: rom = 27;
		4226: rom = 27;
		4227: rom = 27;
		4228: rom = 27;
		4229: rom = 27;
		4230: rom = 27;
		4231: rom = 27;
		4232: rom = 27;
		4233: rom = 27;
		4234: rom = 27;
		4235: rom = 27;
		4236: rom = 27;
		4237: rom = 27;
		4238: rom = 27;
		4239: rom = 27;
		4240: rom = 27;
		4241: rom = 27;
		4242: rom = 27;
		4243: rom = 22;
		4244: rom = 14;
		4245: rom = 15;
		4246: rom = 16;
		4247: rom = 24;
		4248: rom = 24;
		4249: rom = 24;
		4250: rom = 24;
		4251: rom = 24;
		4252: rom = 24;
		4253: rom = 24;
		4254: rom = 17;
		4255: rom = 21;
		4256: rom = 24;
		4257: rom = 24;
		4258: rom = 24;
		4259: rom = 16;
		4260: rom = 7;
		4261: rom = 13;
		4262: rom = 13;
		4263: rom = 15;
		4264: rom = 9;
		4265: rom = 22;
		4266: rom = 23;
		4267: rom = 12;
		4268: rom = 18;
		4269: rom = 18;
		4270: rom = 15;
		4271: rom = 27;
		4272: rom = 27;
		4273: rom = 27;
		4274: rom = 27;
		4275: rom = 27;
		4276: rom = 27;
		4277: rom = 27;
		4278: rom = 27;
		4279: rom = 27;
		4280: rom = 27;
		4281: rom = 27;
		4282: rom = 27;
		4283: rom = 27;
		4284: rom = 21;
		4285: rom = 21;
		4286: rom = 14;
		4287: rom = 26;
		4288: rom = 27;
		4289: rom = 25;
		4290: rom = 17;
		4291: rom = 24;
		4292: rom = 24;
		4293: rom = 20;
		4294: rom = 23;
		4295: rom = 17;
		4296: rom = 24;
		4297: rom = 24;
		4298: rom = 24;
		4299: rom = 24;
		4300: rom = 17;
		4301: rom = 26;
		4302: rom = 27;
		4303: rom = 27;
		4304: rom = 14;
		4305: rom = 23;
		4306: rom = 17;
		4307: rom = 27;
		4308: rom = 27;
		4309: rom = 27;
		4310: rom = 27;
		4311: rom = 26;
		4312: rom = 0;
		4313: rom = 0;
		4314: rom = 0;
		4315: rom = 23;
		4316: rom = 27;
		4317: rom = 27;
		4318: rom = 27;
		4319: rom = 27;
		4320: rom = 27;
		4321: rom = 27;
		4322: rom = 27;
		4323: rom = 27;
		4324: rom = 27;
		4325: rom = 27;
		4326: rom = 27;
		4327: rom = 27;
		4328: rom = 27;
		4329: rom = 27;
		4330: rom = 27;
		4331: rom = 27;
		4332: rom = 16;
		4333: rom = 0;
		4334: rom = 0;
		4335: rom = 12;
		4336: rom = 23;
		4337: rom = 23;
		4338: rom = 23;
		4339: rom = 6;
		4340: rom = 0;
		4341: rom = 0;
		4342: rom = 15;
		4343: rom = 22;
		4344: rom = 22;
		4345: rom = 22;
		4346: rom = 24;
		4352: rom = 26;
		4353: rom = 13;
		4354: rom = 18;
		4355: rom = 22;
		4356: rom = 25;
		4357: rom = 27;
		4358: rom = 27;
		4359: rom = 27;
		4360: rom = 27;
		4361: rom = 27;
		4362: rom = 27;
		4363: rom = 27;
		4364: rom = 27;
		4365: rom = 27;
		4366: rom = 27;
		4367: rom = 27;
		4368: rom = 27;
		4369: rom = 27;
		4370: rom = 27;
		4371: rom = 27;
		4372: rom = 13;
		4373: rom = 11;
		4374: rom = 23;
		4375: rom = 24;
		4376: rom = 24;
		4377: rom = 24;
		4378: rom = 24;
		4379: rom = 22;
		4380: rom = 19;
		4381: rom = 17;
		4382: rom = 17;
		4383: rom = 17;
		4384: rom = 24;
		4385: rom = 24;
		4386: rom = 24;
		4387: rom = 14;
		4388: rom = 21;
		4389: rom = 19;
		4390: rom = 16;
		4391: rom = 14;
		4392: rom = 6;
		4393: rom = 15;
		4394: rom = 12;
		4395: rom = 16;
		4396: rom = 18;
		4397: rom = 17;
		4398: rom = 17;
		4399: rom = 27;
		4400: rom = 27;
		4401: rom = 27;
		4402: rom = 27;
		4403: rom = 27;
		4404: rom = 27;
		4405: rom = 27;
		4406: rom = 27;
		4407: rom = 27;
		4408: rom = 27;
		4409: rom = 27;
		4410: rom = 27;
		4411: rom = 27;
		4412: rom = 18;
		4413: rom = 23;
		4414: rom = 22;
		4415: rom = 18;
		4416: rom = 27;
		4417: rom = 24;
		4418: rom = 18;
		4419: rom = 24;
		4420: rom = 24;
		4421: rom = 21;
		4422: rom = 21;
		4423: rom = 15;
		4424: rom = 24;
		4425: rom = 24;
		4426: rom = 24;
		4427: rom = 24;
		4428: rom = 17;
		4429: rom = 26;
		4430: rom = 27;
		4431: rom = 22;
		4432: rom = 19;
		4433: rom = 24;
		4434: rom = 17;
		4435: rom = 27;
		4436: rom = 27;
		4437: rom = 27;
		4438: rom = 27;
		4439: rom = 27;
		4440: rom = 9;
		4441: rom = 0;
		4442: rom = 0;
		4443: rom = 19;
		4444: rom = 27;
		4445: rom = 27;
		4446: rom = 27;
		4447: rom = 27;
		4448: rom = 27;
		4449: rom = 27;
		4450: rom = 27;
		4451: rom = 27;
		4452: rom = 27;
		4453: rom = 27;
		4454: rom = 27;
		4455: rom = 27;
		4456: rom = 27;
		4457: rom = 27;
		4458: rom = 27;
		4459: rom = 27;
		4460: rom = 9;
		4461: rom = 0;
		4462: rom = 0;
		4463: rom = 20;
		4464: rom = 27;
		4465: rom = 27;
		4466: rom = 27;
		4467: rom = 8;
		4468: rom = 0;
		4469: rom = 0;
		4470: rom = 19;
		4471: rom = 27;
		4472: rom = 27;
		4473: rom = 27;
		4474: rom = 27;
		4480: rom = 27;
		4481: rom = 21;
		4482: rom = 14;
		4483: rom = 15;
		4484: rom = 13;
		4485: rom = 10;
		4486: rom = 10;
		4487: rom = 12;
		4488: rom = 12;
		4489: rom = 12;
		4490: rom = 13;
		4491: rom = 15;
		4492: rom = 16;
		4493: rom = 18;
		4494: rom = 20;
		4495: rom = 24;
		4496: rom = 26;
		4497: rom = 27;
		4498: rom = 27;
		4499: rom = 20;
		4500: rom = 15;
		4501: rom = 14;
		4502: rom = 24;
		4503: rom = 24;
		4504: rom = 24;
		4505: rom = 23;
		4506: rom = 15;
		4507: rom = 14;
		4508: rom = 19;
		4509: rom = 21;
		4510: rom = 20;
		4511: rom = 22;
		4512: rom = 24;
		4513: rom = 24;
		4514: rom = 16;
		4515: rom = 17;
		4516: rom = 25;
		4517: rom = 22;
		4518: rom = 18;
		4519: rom = 18;
		4520: rom = 11;
		4521: rom = 17;
		4522: rom = 16;
		4523: rom = 17;
		4524: rom = 18;
		4525: rom = 14;
		4526: rom = 23;
		4527: rom = 27;
		4528: rom = 27;
		4529: rom = 27;
		4530: rom = 27;
		4531: rom = 27;
		4532: rom = 27;
		4533: rom = 27;
		4534: rom = 26;
		4535: rom = 18;
		4536: rom = 12;
		4537: rom = 15;
		4538: rom = 20;
		4539: rom = 26;
		4540: rom = 17;
		4541: rom = 24;
		4542: rom = 24;
		4543: rom = 15;
		4544: rom = 26;
		4545: rom = 23;
		4546: rom = 21;
		4547: rom = 24;
		4548: rom = 24;
		4549: rom = 22;
		4550: rom = 19;
		4551: rom = 15;
		4552: rom = 24;
		4553: rom = 24;
		4554: rom = 24;
		4555: rom = 24;
		4556: rom = 17;
		4557: rom = 26;
		4558: rom = 27;
		4559: rom = 14;
		4560: rom = 23;
		4561: rom = 24;
		4562: rom = 17;
		4563: rom = 27;
		4564: rom = 27;
		4565: rom = 27;
		4566: rom = 27;
		4567: rom = 27;
		4568: rom = 17;
		4569: rom = 0;
		4570: rom = 0;
		4571: rom = 10;
		4572: rom = 27;
		4573: rom = 27;
		4574: rom = 27;
		4575: rom = 27;
		4576: rom = 27;
		4577: rom = 27;
		4578: rom = 27;
		4579: rom = 27;
		4580: rom = 27;
		4581: rom = 27;
		4582: rom = 27;
		4583: rom = 27;
		4584: rom = 27;
		4585: rom = 27;
		4586: rom = 27;
		4587: rom = 24;
		4588: rom = 0;
		4589: rom = 0;
		4590: rom = 0;
		4591: rom = 24;
		4592: rom = 27;
		4593: rom = 27;
		4594: rom = 27;
		4595: rom = 8;
		4596: rom = 0;
		4597: rom = 0;
		4598: rom = 19;
		4599: rom = 27;
		4600: rom = 27;
		4601: rom = 27;
		4602: rom = 27;
		4608: rom = 27;
		4609: rom = 27;
		4610: rom = 15;
		4611: rom = 17;
		4612: rom = 18;
		4613: rom = 18;
		4614: rom = 18;
		4615: rom = 18;
		4616: rom = 18;
		4617: rom = 18;
		4618: rom = 18;
		4619: rom = 18;
		4620: rom = 18;
		4621: rom = 17;
		4622: rom = 16;
		4623: rom = 14;
		4624: rom = 10;
		4625: rom = 15;
		4626: rom = 22;
		4627: rom = 15;
		4628: rom = 14;
		4629: rom = 17;
		4630: rom = 24;
		4631: rom = 24;
		4632: rom = 22;
		4633: rom = 12;
		4634: rom = 21;
		4635: rom = 24;
		4636: rom = 24;
		4637: rom = 24;
		4638: rom = 24;
		4639: rom = 24;
		4640: rom = 24;
		4641: rom = 17;
		4642: rom = 13;
		4643: rom = 20;
		4644: rom = 25;
		4645: rom = 22;
		4646: rom = 18;
		4647: rom = 18;
		4648: rom = 14;
		4649: rom = 16;
		4650: rom = 10;
		4651: rom = 12;
		4652: rom = 18;
		4653: rom = 11;
		4654: rom = 27;
		4655: rom = 27;
		4656: rom = 27;
		4657: rom = 27;
		4658: rom = 27;
		4659: rom = 27;
		4660: rom = 27;
		4661: rom = 24;
		4662: rom = 11;
		4663: rom = 16;
		4664: rom = 18;
		4665: rom = 17;
		4666: rom = 15;
		4667: rom = 10;
		4668: rom = 11;
		4669: rom = 24;
		4670: rom = 24;
		4671: rom = 21;
		4672: rom = 21;
		4673: rom = 21;
		4674: rom = 21;
		4675: rom = 24;
		4676: rom = 24;
		4677: rom = 22;
		4678: rom = 14;
		4679: rom = 18;
		4680: rom = 24;
		4681: rom = 24;
		4682: rom = 24;
		4683: rom = 24;
		4684: rom = 17;
		4685: rom = 27;
		4686: rom = 23;
		4687: rom = 18;
		4688: rom = 24;
		4689: rom = 24;
		4690: rom = 17;
		4691: rom = 27;
		4692: rom = 27;
		4693: rom = 27;
		4694: rom = 27;
		4695: rom = 27;
		4696: rom = 23;
		4697: rom = 0;
		4698: rom = 0;
		4699: rom = 0;
		4700: rom = 23;
		4701: rom = 27;
		4702: rom = 27;
		4703: rom = 27;
		4704: rom = 27;
		4705: rom = 27;
		4706: rom = 27;
		4707: rom = 27;
		4708: rom = 27;
		4709: rom = 27;
		4710: rom = 27;
		4711: rom = 27;
		4712: rom = 27;
		4713: rom = 27;
		4714: rom = 27;
		4715: rom = 16;
		4716: rom = 0;
		4717: rom = 0;
		4718: rom = 8;
		4719: rom = 27;
		4720: rom = 27;
		4721: rom = 27;
		4722: rom = 27;
		4723: rom = 8;
		4724: rom = 0;
		4725: rom = 0;
		4726: rom = 19;
		4727: rom = 27;
		4728: rom = 27;
		4729: rom = 27;
		4730: rom = 27;
		4736: rom = 27;
		4737: rom = 27;
		4738: rom = 26;
		4739: rom = 12;
		4740: rom = 18;
		4741: rom = 18;
		4742: rom = 18;
		4743: rom = 18;
		4744: rom = 18;
		4745: rom = 18;
		4746: rom = 18;
		4747: rom = 18;
		4748: rom = 18;
		4749: rom = 18;
		4750: rom = 18;
		4751: rom = 18;
		4752: rom = 18;
		4753: rom = 18;
		4754: rom = 15;
		4755: rom = 13;
		4756: rom = 21;
		4757: rom = 17;
		4758: rom = 24;
		4759: rom = 23;
		4760: rom = 13;
		4761: rom = 21;
		4762: rom = 22;
		4763: rom = 24;
		4764: rom = 24;
		4765: rom = 24;
		4766: rom = 24;
		4767: rom = 23;
		4768: rom = 15;
		4769: rom = 13;
		4770: rom = 18;
		4771: rom = 20;
		4772: rom = 25;
		4773: rom = 22;
		4774: rom = 18;
		4775: rom = 18;
		4776: rom = 14;
		4777: rom = 8;
		4778: rom = 16;
		4779: rom = 11;
		4780: rom = 17;
		4781: rom = 18;
		4782: rom = 27;
		4783: rom = 27;
		4784: rom = 27;
		4785: rom = 27;
		4786: rom = 27;
		4787: rom = 27;
		4788: rom = 24;
		4789: rom = 11;
		4790: rom = 17;
		4791: rom = 18;
		4792: rom = 18;
		4793: rom = 18;
		4794: rom = 18;
		4795: rom = 17;
		4796: rom = 9;
		4797: rom = 23;
		4798: rom = 24;
		4799: rom = 23;
		4800: rom = 16;
		4801: rom = 20;
		4802: rom = 21;
		4803: rom = 24;
		4804: rom = 24;
		4805: rom = 23;
		4806: rom = 7;
		4807: rom = 20;
		4808: rom = 24;
		4809: rom = 24;
		4810: rom = 24;
		4811: rom = 24;
		4812: rom = 15;
		4813: rom = 27;
		4814: rom = 15;
		4815: rom = 23;
		4816: rom = 24;
		4817: rom = 24;
		4818: rom = 16;
		4819: rom = 27;
		4820: rom = 27;
		4821: rom = 27;
		4822: rom = 27;
		4823: rom = 27;
		4824: rom = 27;
		4825: rom = 9;
		4826: rom = 0;
		4827: rom = 0;
		4828: rom = 10;
		4829: rom = 27;
		4830: rom = 27;
		4831: rom = 27;
		4832: rom = 27;
		4833: rom = 27;
		4834: rom = 27;
		4835: rom = 27;
		4836: rom = 27;
		4837: rom = 27;
		4838: rom = 27;
		4839: rom = 27;
		4840: rom = 27;
		4841: rom = 27;
		4842: rom = 23;
		4843: rom = 0;
		4844: rom = 0;
		4845: rom = 0;
		4846: rom = 19;
		4847: rom = 27;
		4848: rom = 27;
		4849: rom = 27;
		4850: rom = 27;
		4851: rom = 10;
		4852: rom = 6;
		4853: rom = 6;
		4854: rom = 19;
		4855: rom = 27;
		4856: rom = 27;
		4857: rom = 27;
		4858: rom = 27;
		4864: rom = 27;
		4865: rom = 27;
		4866: rom = 27;
		4867: rom = 24;
		4868: rom = 12;
		4869: rom = 18;
		4870: rom = 18;
		4871: rom = 18;
		4872: rom = 18;
		4873: rom = 18;
		4874: rom = 18;
		4875: rom = 18;
		4876: rom = 19;
		4877: rom = 19;
		4878: rom = 18;
		4879: rom = 18;
		4880: rom = 18;
		4881: rom = 18;
		4882: rom = 18;
		4883: rom = 12;
		4884: rom = 23;
		4885: rom = 14;
		4886: rom = 24;
		4887: rom = 18;
		4888: rom = 8;
		4889: rom = 13;
		4890: rom = 14;
		4891: rom = 14;
		4892: rom = 14;
		4893: rom = 20;
		4894: rom = 19;
		4895: rom = 11;
		4896: rom = 12;
		4897: rom = 12;
		4898: rom = 15;
		4899: rom = 19;
		4900: rom = 25;
		4901: rom = 22;
		4902: rom = 18;
		4903: rom = 18;
		4904: rom = 13;
		4905: rom = 16;
		4906: rom = 18;
		4907: rom = 11;
		4908: rom = 12;
		4909: rom = 25;
		4910: rom = 27;
		4911: rom = 27;
		4912: rom = 27;
		4913: rom = 27;
		4914: rom = 27;
		4915: rom = 26;
		4916: rom = 11;
		4917: rom = 17;
		4918: rom = 18;
		4919: rom = 18;
		4920: rom = 18;
		4921: rom = 18;
		4922: rom = 18;
		4923: rom = 18;
		4924: rom = 13;
		4925: rom = 22;
		4926: rom = 24;
		4927: rom = 24;
		4928: rom = 15;
		4929: rom = 18;
		4930: rom = 21;
		4931: rom = 24;
		4932: rom = 24;
		4933: rom = 23;
		4934: rom = 2;
		4935: rom = 22;
		4936: rom = 24;
		4937: rom = 24;
		4938: rom = 24;
		4939: rom = 24;
		4940: rom = 14;
		4941: rom = 25;
		4942: rom = 17;
		4943: rom = 24;
		4944: rom = 24;
		4945: rom = 23;
		4946: rom = 18;
		4947: rom = 27;
		4948: rom = 27;
		4949: rom = 27;
		4950: rom = 27;
		4951: rom = 27;
		4952: rom = 27;
		4953: rom = 21;
		4954: rom = 0;
		4955: rom = 0;
		4956: rom = 0;
		4957: rom = 16;
		4958: rom = 27;
		4959: rom = 27;
		4960: rom = 27;
		4961: rom = 27;
		4962: rom = 27;
		4963: rom = 27;
		4964: rom = 27;
		4965: rom = 27;
		4966: rom = 27;
		4967: rom = 27;
		4968: rom = 27;
		4969: rom = 25;
		4970: rom = 8;
		4971: rom = 0;
		4972: rom = 0;
		4973: rom = 5;
		4974: rom = 26;
		4975: rom = 27;
		4976: rom = 27;
		4977: rom = 27;
		4978: rom = 27;
		4979: rom = 27;
		4980: rom = 27;
		4981: rom = 27;
		4982: rom = 27;
		4983: rom = 27;
		4984: rom = 27;
		4985: rom = 27;
		4986: rom = 27;
		4992: rom = 27;
		4993: rom = 27;
		4994: rom = 27;
		4995: rom = 27;
		4996: rom = 21;
		4997: rom = 14;
		4998: rom = 18;
		4999: rom = 18;
		5000: rom = 19;
		5001: rom = 22;
		5002: rom = 24;
		5003: rom = 25;
		5004: rom = 25;
		5005: rom = 25;
		5006: rom = 25;
		5007: rom = 24;
		5008: rom = 23;
		5009: rom = 22;
		5010: rom = 19;
		5011: rom = 14;
		5012: rom = 20;
		5013: rom = 14;
		5014: rom = 21;
		5015: rom = 14;
		5016: rom = 23;
		5017: rom = 24;
		5018: rom = 24;
		5019: rom = 24;
		5020: rom = 23;
		5021: rom = 18;
		5022: rom = 9;
		5023: rom = 22;
		5024: rom = 24;
		5025: rom = 21;
		5026: rom = 18;
		5027: rom = 14;
		5028: rom = 13;
		5029: rom = 13;
		5030: rom = 18;
		5031: rom = 18;
		5032: rom = 17;
		5033: rom = 18;
		5034: rom = 18;
		5035: rom = 7;
		5036: rom = 8;
		5037: rom = 20;
		5038: rom = 27;
		5039: rom = 27;
		5040: rom = 27;
		5041: rom = 27;
		5042: rom = 27;
		5043: rom = 17;
		5044: rom = 16;
		5045: rom = 18;
		5046: rom = 18;
		5047: rom = 18;
		5048: rom = 18;
		5049: rom = 18;
		5050: rom = 18;
		5051: rom = 18;
		5052: rom = 14;
		5053: rom = 20;
		5054: rom = 24;
		5055: rom = 24;
		5056: rom = 19;
		5057: rom = 11;
		5058: rom = 22;
		5059: rom = 24;
		5060: rom = 24;
		5061: rom = 23;
		5062: rom = 3;
		5063: rom = 23;
		5064: rom = 24;
		5065: rom = 24;
		5066: rom = 24;
		5067: rom = 24;
		5068: rom = 16;
		5069: rom = 17;
		5070: rom = 22;
		5071: rom = 24;
		5072: rom = 24;
		5073: rom = 22;
		5074: rom = 19;
		5075: rom = 27;
		5076: rom = 27;
		5077: rom = 27;
		5078: rom = 27;
		5079: rom = 27;
		5080: rom = 27;
		5081: rom = 26;
		5082: rom = 3;
		5083: rom = 0;
		5084: rom = 0;
		5085: rom = 0;
		5086: rom = 16;
		5087: rom = 27;
		5088: rom = 27;
		5089: rom = 27;
		5090: rom = 27;
		5091: rom = 27;
		5092: rom = 27;
		5093: rom = 27;
		5094: rom = 27;
		5095: rom = 27;
		5096: rom = 25;
		5097: rom = 9;
		5098: rom = 0;
		5099: rom = 0;
		5100: rom = 0;
		5101: rom = 20;
		5102: rom = 27;
		5103: rom = 27;
		5104: rom = 27;
		5105: rom = 27;
		5106: rom = 27;
		5107: rom = 27;
		5108: rom = 27;
		5109: rom = 27;
		5110: rom = 27;
		5111: rom = 27;
		5112: rom = 27;
		5113: rom = 27;
		5114: rom = 27;
		5120: rom = 27;
		5121: rom = 27;
		5122: rom = 27;
		5123: rom = 27;
		5124: rom = 27;
		5125: rom = 18;
		5126: rom = 15;
		5127: rom = 19;
		5128: rom = 24;
		5129: rom = 25;
		5130: rom = 25;
		5131: rom = 25;
		5132: rom = 25;
		5133: rom = 25;
		5134: rom = 25;
		5135: rom = 25;
		5136: rom = 25;
		5137: rom = 25;
		5138: rom = 25;
		5139: rom = 19;
		5140: rom = 13;
		5141: rom = 17;
		5142: rom = 21;
		5143: rom = 23;
		5144: rom = 24;
		5145: rom = 24;
		5146: rom = 24;
		5147: rom = 24;
		5148: rom = 24;
		5149: rom = 24;
		5150: rom = 22;
		5151: rom = 14;
		5152: rom = 24;
		5153: rom = 24;
		5154: rom = 24;
		5155: rom = 24;
		5156: rom = 24;
		5157: rom = 20;
		5158: rom = 9;
		5159: rom = 15;
		5160: rom = 18;
		5161: rom = 18;
		5162: rom = 17;
		5163: rom = 13;
		5164: rom = 16;
		5165: rom = 21;
		5166: rom = 27;
		5167: rom = 27;
		5168: rom = 27;
		5169: rom = 27;
		5170: rom = 25;
		5171: rom = 12;
		5172: rom = 18;
		5173: rom = 18;
		5174: rom = 18;
		5175: rom = 18;
		5176: rom = 18;
		5177: rom = 18;
		5178: rom = 18;
		5179: rom = 18;
		5180: rom = 16;
		5181: rom = 16;
		5182: rom = 24;
		5183: rom = 24;
		5184: rom = 21;
		5185: rom = 1;
		5186: rom = 22;
		5187: rom = 24;
		5188: rom = 24;
		5189: rom = 23;
		5190: rom = 10;
		5191: rom = 24;
		5192: rom = 24;
		5193: rom = 24;
		5194: rom = 24;
		5195: rom = 24;
		5196: rom = 16;
		5197: rom = 15;
		5198: rom = 24;
		5199: rom = 24;
		5200: rom = 24;
		5201: rom = 21;
		5202: rom = 21;
		5203: rom = 27;
		5204: rom = 27;
		5205: rom = 27;
		5206: rom = 27;
		5207: rom = 27;
		5208: rom = 27;
		5209: rom = 15;
		5210: rom = 0;
		5211: rom = 0;
		5212: rom = 0;
		5213: rom = 0;
		5214: rom = 0;
		5215: rom = 10;
		5216: rom = 22;
		5217: rom = 27;
		5218: rom = 27;
		5219: rom = 27;
		5220: rom = 27;
		5221: rom = 27;
		5222: rom = 26;
		5223: rom = 19;
		5224: rom = 4;
		5225: rom = 0;
		5226: rom = 0;
		5227: rom = 0;
		5228: rom = 14;
		5229: rom = 27;
		5230: rom = 27;
		5231: rom = 27;
		5232: rom = 27;
		5233: rom = 27;
		5234: rom = 27;
		5235: rom = 27;
		5236: rom = 27;
		5237: rom = 27;
		5238: rom = 27;
		5239: rom = 27;
		5240: rom = 27;
		5241: rom = 27;
		5242: rom = 27;
		5248: rom = 27;
		5249: rom = 27;
		5250: rom = 27;
		5251: rom = 27;
		5252: rom = 27;
		5253: rom = 27;
		5254: rom = 16;
		5255: rom = 20;
		5256: rom = 25;
		5257: rom = 23;
		5258: rom = 20;
		5259: rom = 18;
		5260: rom = 18;
		5261: rom = 18;
		5262: rom = 18;
		5263: rom = 19;
		5264: rom = 21;
		5265: rom = 22;
		5266: rom = 24;
		5267: rom = 13;
		5268: rom = 11;
		5269: rom = 21;
		5270: rom = 24;
		5271: rom = 24;
		5272: rom = 24;
		5273: rom = 24;
		5274: rom = 24;
		5275: rom = 24;
		5276: rom = 24;
		5277: rom = 24;
		5278: rom = 23;
		5279: rom = 13;
		5280: rom = 24;
		5281: rom = 24;
		5282: rom = 24;
		5283: rom = 24;
		5284: rom = 24;
		5285: rom = 18;
		5286: rom = 5;
		5287: rom = 5;
		5288: rom = 14;
		5289: rom = 18;
		5290: rom = 17;
		5291: rom = 18;
		5292: rom = 14;
		5293: rom = 24;
		5294: rom = 27;
		5295: rom = 27;
		5296: rom = 27;
		5297: rom = 27;
		5298: rom = 17;
		5299: rom = 17;
		5300: rom = 18;
		5301: rom = 18;
		5302: rom = 18;
		5303: rom = 22;
		5304: rom = 24;
		5305: rom = 23;
		5306: rom = 19;
		5307: rom = 18;
		5308: rom = 18;
		5309: rom = 14;
		5310: rom = 24;
		5311: rom = 24;
		5312: rom = 23;
		5313: rom = 4;
		5314: rom = 23;
		5315: rom = 24;
		5316: rom = 24;
		5317: rom = 23;
		5318: rom = 14;
		5319: rom = 24;
		5320: rom = 24;
		5321: rom = 24;
		5322: rom = 24;
		5323: rom = 24;
		5324: rom = 8;
		5325: rom = 21;
		5326: rom = 24;
		5327: rom = 24;
		5328: rom = 24;
		5329: rom = 20;
		5330: rom = 23;
		5331: rom = 27;
		5332: rom = 27;
		5333: rom = 27;
		5334: rom = 27;
		5335: rom = 27;
		5336: rom = 18;
		5337: rom = 0;
		5338: rom = 0;
		5339: rom = 0;
		5340: rom = 0;
		5341: rom = 0;
		5342: rom = 0;
		5343: rom = 0;
		5344: rom = 0;
		5345: rom = 6;
		5346: rom = 15;
		5347: rom = 17;
		5348: rom = 16;
		5349: rom = 13;
		5350: rom = 0;
		5351: rom = 0;
		5352: rom = 0;
		5353: rom = 0;
		5354: rom = 0;
		5355: rom = 12;
		5356: rom = 26;
		5357: rom = 27;
		5358: rom = 27;
		5359: rom = 27;
		5360: rom = 27;
		5361: rom = 27;
		5362: rom = 27;
		5363: rom = 27;
		5364: rom = 27;
		5365: rom = 27;
		5366: rom = 27;
		5367: rom = 27;
		5368: rom = 27;
		5369: rom = 27;
		5370: rom = 27;
		5376: rom = 27;
		5377: rom = 27;
		5378: rom = 27;
		5379: rom = 27;
		5380: rom = 27;
		5381: rom = 27;
		5382: rom = 27;
		5383: rom = 16;
		5384: rom = 21;
		5385: rom = 18;
		5386: rom = 18;
		5387: rom = 18;
		5388: rom = 18;
		5389: rom = 18;
		5390: rom = 18;
		5391: rom = 18;
		5392: rom = 18;
		5393: rom = 18;
		5394: rom = 18;
		5395: rom = 12;
		5396: rom = 21;
		5397: rom = 15;
		5398: rom = 24;
		5399: rom = 24;
		5400: rom = 24;
		5401: rom = 24;
		5402: rom = 24;
		5403: rom = 24;
		5404: rom = 24;
		5405: rom = 20;
		5406: rom = 12;
		5407: rom = 19;
		5408: rom = 24;
		5409: rom = 24;
		5410: rom = 24;
		5411: rom = 24;
		5412: rom = 20;
		5413: rom = 4;
		5414: rom = 7;
		5415: rom = 7;
		5416: rom = 14;
		5417: rom = 18;
		5418: rom = 18;
		5419: rom = 18;
		5420: rom = 11;
		5421: rom = 27;
		5422: rom = 27;
		5423: rom = 27;
		5424: rom = 27;
		5425: rom = 25;
		5426: rom = 12;
		5427: rom = 18;
		5428: rom = 18;
		5429: rom = 18;
		5430: rom = 23;
		5431: rom = 25;
		5432: rom = 25;
		5433: rom = 25;
		5434: rom = 25;
		5435: rom = 19;
		5436: rom = 18;
		5437: rom = 18;
		5438: rom = 23;
		5439: rom = 24;
		5440: rom = 24;
		5441: rom = 12;
		5442: rom = 23;
		5443: rom = 24;
		5444: rom = 24;
		5445: rom = 22;
		5446: rom = 16;
		5447: rom = 24;
		5448: rom = 24;
		5449: rom = 24;
		5450: rom = 24;
		5451: rom = 23;
		5452: rom = 10;
		5453: rom = 24;
		5454: rom = 24;
		5455: rom = 24;
		5456: rom = 24;
		5457: rom = 18;
		5458: rom = 25;
		5459: rom = 27;
		5460: rom = 26;
		5461: rom = 27;
		5462: rom = 27;
		5463: rom = 20;
		5464: rom = 0;
		5465: rom = 0;
		5466: rom = 0;
		5467: rom = 0;
		5468: rom = 11;
		5469: rom = 7;
		5470: rom = 0;
		5471: rom = 0;
		5472: rom = 0;
		5473: rom = 0;
		5474: rom = 0;
		5475: rom = 0;
		5476: rom = 0;
		5477: rom = 0;
		5478: rom = 0;
		5479: rom = 0;
		5480: rom = 0;
		5481: rom = 0;
		5482: rom = 15;
		5483: rom = 26;
		5484: rom = 27;
		5485: rom = 27;
		5486: rom = 27;
		5487: rom = 27;
		5488: rom = 27;
		5489: rom = 27;
		5490: rom = 27;
		5491: rom = 27;
		5492: rom = 27;
		5493: rom = 27;
		5494: rom = 27;
		5495: rom = 27;
		5496: rom = 27;
		5497: rom = 27;
		5498: rom = 27;
		5504: rom = 27;
		5505: rom = 27;
		5506: rom = 27;
		5507: rom = 27;
		5508: rom = 27;
		5509: rom = 27;
		5510: rom = 27;
		5511: rom = 27;
		5512: rom = 16;
		5513: rom = 15;
		5514: rom = 18;
		5515: rom = 18;
		5516: rom = 18;
		5517: rom = 18;
		5518: rom = 18;
		5519: rom = 18;
		5520: rom = 18;
		5521: rom = 18;
		5522: rom = 18;
		5523: rom = 13;
		5524: rom = 21;
		5525: rom = 16;
		5526: rom = 22;
		5527: rom = 24;
		5528: rom = 24;
		5529: rom = 24;
		5530: rom = 24;
		5531: rom = 22;
		5532: rom = 13;
		5533: rom = 17;
		5534: rom = 23;
		5535: rom = 24;
		5536: rom = 24;
		5537: rom = 24;
		5538: rom = 24;
		5539: rom = 20;
		5540: rom = 13;
		5541: rom = 14;
		5542: rom = 6;
		5543: rom = 7;
		5544: rom = 16;
		5545: rom = 18;
		5546: rom = 18;
		5547: rom = 18;
		5548: rom = 8;
		5549: rom = 16;
		5550: rom = 25;
		5551: rom = 27;
		5552: rom = 26;
		5553: rom = 16;
		5554: rom = 16;
		5555: rom = 18;
		5556: rom = 18;
		5557: rom = 21;
		5558: rom = 25;
		5559: rom = 24;
		5560: rom = 20;
		5561: rom = 23;
		5562: rom = 25;
		5563: rom = 23;
		5564: rom = 18;
		5565: rom = 18;
		5566: rom = 19;
		5567: rom = 23;
		5568: rom = 24;
		5569: rom = 16;
		5570: rom = 23;
		5571: rom = 24;
		5572: rom = 24;
		5573: rom = 21;
		5574: rom = 19;
		5575: rom = 24;
		5576: rom = 24;
		5577: rom = 24;
		5578: rom = 24;
		5579: rom = 20;
		5580: rom = 18;
		5581: rom = 24;
		5582: rom = 24;
		5583: rom = 24;
		5584: rom = 24;
		5585: rom = 16;
		5586: rom = 25;
		5587: rom = 16;
		5588: rom = 18;
		5589: rom = 27;
		5590: rom = 22;
		5591: rom = 1;
		5592: rom = 0;
		5593: rom = 0;
		5594: rom = 0;
		5595: rom = 9;
		5596: rom = 26;
		5597: rom = 26;
		5598: rom = 16;
		5599: rom = 0;
		5600: rom = 0;
		5601: rom = 0;
		5602: rom = 0;
		5603: rom = 0;
		5604: rom = 0;
		5605: rom = 0;
		5606: rom = 0;
		5607: rom = 0;
		5608: rom = 7;
		5609: rom = 21;
		5610: rom = 27;
		5611: rom = 27;
		5612: rom = 27;
		5613: rom = 27;
		5614: rom = 27;
		5615: rom = 27;
		5616: rom = 27;
		5617: rom = 27;
		5618: rom = 27;
		5619: rom = 27;
		5620: rom = 27;
		5621: rom = 27;
		5622: rom = 27;
		5623: rom = 27;
		5624: rom = 27;
		5625: rom = 27;
		5626: rom = 27;
		5632: rom = 27;
		5633: rom = 27;
		5634: rom = 27;
		5635: rom = 27;
		5636: rom = 27;
		5637: rom = 27;
		5638: rom = 27;
		5639: rom = 27;
		5640: rom = 27;
		5641: rom = 16;
		5642: rom = 15;
		5643: rom = 18;
		5644: rom = 18;
		5645: rom = 18;
		5646: rom = 18;
		5647: rom = 18;
		5648: rom = 18;
		5649: rom = 18;
		5650: rom = 18;
		5651: rom = 16;
		5652: rom = 16;
		5653: rom = 22;
		5654: rom = 18;
		5655: rom = 24;
		5656: rom = 24;
		5657: rom = 24;
		5658: rom = 21;
		5659: rom = 13;
		5660: rom = 22;
		5661: rom = 24;
		5662: rom = 24;
		5663: rom = 24;
		5664: rom = 24;
		5665: rom = 24;
		5666: rom = 17;
		5667: rom = 15;
		5668: rom = 22;
		5669: rom = 20;
		5670: rom = 5;
		5671: rom = 9;
		5672: rom = 18;
		5673: rom = 18;
		5674: rom = 18;
		5675: rom = 18;
		5676: rom = 13;
		5677: rom = 16;
		5678: rom = 12;
		5679: rom = 10;
		5680: rom = 10;
		5681: rom = 9;
		5682: rom = 18;
		5683: rom = 16;
		5684: rom = 18;
		5685: rom = 24;
		5686: rom = 25;
		5687: rom = 20;
		5688: rom = 18;
		5689: rom = 18;
		5690: rom = 24;
		5691: rom = 25;
		5692: rom = 19;
		5693: rom = 18;
		5694: rom = 18;
		5695: rom = 20;
		5696: rom = 24;
		5697: rom = 17;
		5698: rom = 23;
		5699: rom = 24;
		5700: rom = 24;
		5701: rom = 18;
		5702: rom = 21;
		5703: rom = 24;
		5704: rom = 24;
		5705: rom = 24;
		5706: rom = 24;
		5707: rom = 15;
		5708: rom = 23;
		5709: rom = 24;
		5710: rom = 24;
		5711: rom = 24;
		5712: rom = 24;
		5713: rom = 15;
		5714: rom = 19;
		5715: rom = 0;
		5716: rom = 18;
		5717: rom = 24;
		5718: rom = 4;
		5719: rom = 0;
		5720: rom = 0;
		5721: rom = 0;
		5722: rom = 7;
		5723: rom = 25;
		5724: rom = 27;
		5725: rom = 27;
		5726: rom = 27;
		5727: rom = 25;
		5728: rom = 19;
		5729: rom = 12;
		5730: rom = 3;
		5731: rom = 0;
		5732: rom = 0;
		5733: rom = 6;
		5734: rom = 14;
		5735: rom = 21;
		5736: rom = 27;
		5737: rom = 27;
		5738: rom = 27;
		5739: rom = 27;
		5740: rom = 27;
		5741: rom = 27;
		5742: rom = 27;
		5743: rom = 27;
		5744: rom = 27;
		5745: rom = 27;
		5746: rom = 27;
		5747: rom = 27;
		5748: rom = 27;
		5749: rom = 27;
		5750: rom = 27;
		5751: rom = 27;
		5752: rom = 27;
		5753: rom = 27;
		5754: rom = 27;
		5760: rom = 27;
		5761: rom = 27;
		5762: rom = 27;
		5763: rom = 27;
		5764: rom = 27;
		5765: rom = 27;
		5766: rom = 27;
		5767: rom = 27;
		5768: rom = 27;
		5769: rom = 27;
		5770: rom = 17;
		5771: rom = 14;
		5772: rom = 18;
		5773: rom = 18;
		5774: rom = 18;
		5775: rom = 18;
		5776: rom = 18;
		5777: rom = 18;
		5778: rom = 18;
		5779: rom = 17;
		5780: rom = 10;
		5781: rom = 19;
		5782: rom = 18;
		5783: rom = 24;
		5784: rom = 24;
		5785: rom = 22;
		5786: rom = 13;
		5787: rom = 23;
		5788: rom = 24;
		5789: rom = 24;
		5790: rom = 24;
		5791: rom = 24;
		5792: rom = 22;
		5793: rom = 12;
		5794: rom = 17;
		5795: rom = 23;
		5796: rom = 23;
		5797: rom = 17;
		5798: rom = 5;
		5799: rom = 14;
		5800: rom = 18;
		5801: rom = 18;
		5802: rom = 18;
		5803: rom = 18;
		5804: rom = 18;
		5805: rom = 18;
		5806: rom = 18;
		5807: rom = 18;
		5808: rom = 18;
		5809: rom = 16;
		5810: rom = 18;
		5811: rom = 12;
		5812: rom = 24;
		5813: rom = 25;
		5814: rom = 22;
		5815: rom = 18;
		5816: rom = 18;
		5817: rom = 18;
		5818: rom = 21;
		5819: rom = 25;
		5820: rom = 22;
		5821: rom = 18;
		5822: rom = 18;
		5823: rom = 18;
		5824: rom = 22;
		5825: rom = 17;
		5826: rom = 23;
		5827: rom = 24;
		5828: rom = 24;
		5829: rom = 16;
		5830: rom = 23;
		5831: rom = 24;
		5832: rom = 24;
		5833: rom = 24;
		5834: rom = 23;
		5835: rom = 16;
		5836: rom = 24;
		5837: rom = 24;
		5838: rom = 24;
		5839: rom = 24;
		5840: rom = 24;
		5841: rom = 16;
		5842: rom = 19;
		5843: rom = 0;
		5844: rom = 14;
		5845: rom = 7;
		5846: rom = 0;
		5847: rom = 0;
		5848: rom = 0;
		5849: rom = 5;
		5850: rom = 24;
		5851: rom = 27;
		5852: rom = 27;
		5853: rom = 27;
		5854: rom = 27;
		5855: rom = 27;
		5856: rom = 27;
		5857: rom = 27;
		5858: rom = 27;
		5859: rom = 26;
		5860: rom = 26;
		5861: rom = 27;
		5862: rom = 27;
		5863: rom = 27;
		5864: rom = 27;
		5865: rom = 27;
		5866: rom = 27;
		5867: rom = 27;
		5868: rom = 27;
		5869: rom = 27;
		5870: rom = 27;
		5871: rom = 27;
		5872: rom = 27;
		5873: rom = 27;
		5874: rom = 27;
		5875: rom = 27;
		5876: rom = 27;
		5877: rom = 27;
		5878: rom = 27;
		5879: rom = 27;
		5880: rom = 27;
		5881: rom = 27;
		5882: rom = 27;
		5888: rom = 27;
		5889: rom = 27;
		5890: rom = 27;
		5891: rom = 27;
		5892: rom = 27;
		5893: rom = 27;
		5894: rom = 27;
		5895: rom = 27;
		5896: rom = 27;
		5897: rom = 27;
		5898: rom = 27;
		5899: rom = 19;
		5900: rom = 12;
		5901: rom = 18;
		5902: rom = 18;
		5903: rom = 18;
		5904: rom = 18;
		5905: rom = 18;
		5906: rom = 17;
		5907: rom = 11;
		5908: rom = 18;
		5909: rom = 19;
		5910: rom = 16;
		5911: rom = 15;
		5912: rom = 23;
		5913: rom = 15;
		5914: rom = 22;
		5915: rom = 19;
		5916: rom = 20;
		5917: rom = 21;
		5918: rom = 19;
		5919: rom = 14;
		5920: rom = 5;
		5921: rom = 4;
		5922: rom = 5;
		5923: rom = 11;
		5924: rom = 11;
		5925: rom = 4;
		5926: rom = 9;
		5927: rom = 18;
		5928: rom = 18;
		5929: rom = 18;
		5930: rom = 18;
		5931: rom = 18;
		5932: rom = 25;
		5933: rom = 24;
		5934: rom = 22;
		5935: rom = 20;
		5936: rom = 19;
		5937: rom = 20;
		5938: rom = 23;
		5939: rom = 15;
		5940: rom = 25;
		5941: rom = 24;
		5942: rom = 18;
		5943: rom = 14;
		5944: rom = 18;
		5945: rom = 18;
		5946: rom = 19;
		5947: rom = 25;
		5948: rom = 24;
		5949: rom = 18;
		5950: rom = 18;
		5951: rom = 18;
		5952: rom = 19;
		5953: rom = 17;
		5954: rom = 22;
		5955: rom = 24;
		5956: rom = 24;
		5957: rom = 14;
		5958: rom = 24;
		5959: rom = 24;
		5960: rom = 24;
		5961: rom = 24;
		5962: rom = 18;
		5963: rom = 21;
		5964: rom = 24;
		5965: rom = 24;
		5966: rom = 24;
		5967: rom = 24;
		5968: rom = 23;
		5969: rom = 17;
		5970: rom = 19;
		5971: rom = 0;
		5972: rom = 0;
		5973: rom = 0;
		5974: rom = 0;
		5975: rom = 0;
		5976: rom = 2;
		5977: rom = 23;
		5978: rom = 27;
		5979: rom = 27;
		5980: rom = 27;
		5981: rom = 27;
		5982: rom = 27;
		5983: rom = 27;
		5984: rom = 27;
		5985: rom = 27;
		5986: rom = 27;
		5987: rom = 27;
		5988: rom = 27;
		5989: rom = 27;
		5990: rom = 27;
		5991: rom = 27;
		5992: rom = 27;
		5993: rom = 27;
		5994: rom = 27;
		5995: rom = 27;
		5996: rom = 27;
		5997: rom = 27;
		5998: rom = 27;
		5999: rom = 27;
		6000: rom = 27;
		6001: rom = 27;
		6002: rom = 27;
		6003: rom = 27;
		6004: rom = 27;
		6005: rom = 27;
		6006: rom = 27;
		6007: rom = 27;
		6008: rom = 27;
		6009: rom = 27;
		6010: rom = 27;
		6016: rom = 27;
		6017: rom = 27;
		6018: rom = 27;
		6019: rom = 27;
		6020: rom = 27;
		6021: rom = 27;
		6022: rom = 27;
		6023: rom = 27;
		6024: rom = 27;
		6025: rom = 27;
		6026: rom = 27;
		6027: rom = 27;
		6028: rom = 22;
		6029: rom = 11;
		6030: rom = 17;
		6031: rom = 18;
		6032: rom = 18;
		6033: rom = 18;
		6034: rom = 17;
		6035: rom = 11;
		6036: rom = 16;
		6037: rom = 22;
		6038: rom = 24;
		6039: rom = 22;
		6040: rom = 13;
		6041: rom = 19;
		6042: rom = 24;
		6043: rom = 23;
		6044: rom = 19;
		6045: rom = 17;
		6046: rom = 19;
		6047: rom = 22;
		6048: rom = 10;
		6049: rom = 7;
		6050: rom = 7;
		6051: rom = 6;
		6052: rom = 7;
		6053: rom = 7;
		6054: rom = 16;
		6055: rom = 18;
		6056: rom = 18;
		6057: rom = 18;
		6058: rom = 18;
		6059: rom = 18;
		6060: rom = 22;
		6061: rom = 25;
		6062: rom = 25;
		6063: rom = 25;
		6064: rom = 25;
		6065: rom = 25;
		6066: rom = 25;
		6067: rom = 15;
		6068: rom = 23;
		6069: rom = 19;
		6070: rom = 18;
		6071: rom = 12;
		6072: rom = 18;
		6073: rom = 18;
		6074: rom = 18;
		6075: rom = 23;
		6076: rom = 25;
		6077: rom = 21;
		6078: rom = 18;
		6079: rom = 18;
		6080: rom = 18;
		6081: rom = 16;
		6082: rom = 22;
		6083: rom = 24;
		6084: rom = 24;
		6085: rom = 15;
		6086: rom = 24;
		6087: rom = 24;
		6088: rom = 24;
		6089: rom = 24;
		6090: rom = 13;
		6091: rom = 24;
		6092: rom = 24;
		6093: rom = 24;
		6094: rom = 24;
		6095: rom = 24;
		6096: rom = 21;
		6097: rom = 21;
		6098: rom = 19;
		6099: rom = 0;
		6100: rom = 0;
		6101: rom = 0;
		6102: rom = 0;
		6103: rom = 0;
		6104: rom = 21;
		6105: rom = 27;
		6106: rom = 27;
		6107: rom = 27;
		6108: rom = 27;
		6109: rom = 27;
		6110: rom = 27;
		6111: rom = 27;
		6112: rom = 27;
		6113: rom = 27;
		6114: rom = 27;
		6115: rom = 27;
		6116: rom = 27;
		6117: rom = 27;
		6118: rom = 27;
		6119: rom = 27;
		6120: rom = 27;
		6121: rom = 27;
		6122: rom = 27;
		6123: rom = 27;
		6124: rom = 27;
		6125: rom = 27;
		6126: rom = 27;
		6127: rom = 27;
		6128: rom = 27;
		6129: rom = 27;
		6130: rom = 27;
		6131: rom = 27;
		6132: rom = 27;
		6133: rom = 27;
		6134: rom = 27;
		6135: rom = 27;
		6136: rom = 27;
		6137: rom = 27;
		6138: rom = 27;
		6144: rom = 27;
		6145: rom = 27;
		6146: rom = 27;
		6147: rom = 27;
		6148: rom = 27;
		6149: rom = 27;
		6150: rom = 27;
		6151: rom = 27;
		6152: rom = 27;
		6153: rom = 27;
		6154: rom = 27;
		6155: rom = 27;
		6156: rom = 27;
		6157: rom = 24;
		6158: rom = 11;
		6159: rom = 16;
		6160: rom = 18;
		6161: rom = 18;
		6162: rom = 18;
		6163: rom = 18;
		6164: rom = 16;
		6165: rom = 10;
		6166: rom = 15;
		6167: rom = 22;
		6168: rom = 21;
		6169: rom = 19;
		6170: rom = 24;
		6171: rom = 24;
		6172: rom = 24;
		6173: rom = 24;
		6174: rom = 24;
		6175: rom = 24;
		6176: rom = 20;
		6177: rom = 4;
		6178: rom = 7;
		6179: rom = 7;
		6180: rom = 7;
		6181: rom = 13;
		6182: rom = 18;
		6183: rom = 18;
		6184: rom = 18;
		6185: rom = 18;
		6186: rom = 16;
		6187: rom = 17;
		6188: rom = 14;
		6189: rom = 20;
		6190: rom = 22;
		6191: rom = 23;
		6192: rom = 24;
		6193: rom = 23;
		6194: rom = 22;
		6195: rom = 12;
		6196: rom = 18;
		6197: rom = 18;
		6198: rom = 18;
		6199: rom = 12;
		6200: rom = 18;
		6201: rom = 18;
		6202: rom = 18;
		6203: rom = 20;
		6204: rom = 25;
		6205: rom = 24;
		6206: rom = 18;
		6207: rom = 18;
		6208: rom = 18;
		6209: rom = 18;
		6210: rom = 23;
		6211: rom = 24;
		6212: rom = 24;
		6213: rom = 14;
		6214: rom = 24;
		6215: rom = 24;
		6216: rom = 24;
		6217: rom = 21;
		6218: rom = 17;
		6219: rom = 24;
		6220: rom = 24;
		6221: rom = 24;
		6222: rom = 24;
		6223: rom = 24;
		6224: rom = 19;
		6225: rom = 24;
		6226: rom = 19;
		6227: rom = 0;
		6228: rom = 0;
		6229: rom = 0;
		6230: rom = 0;
		6231: rom = 18;
		6232: rom = 26;
		6233: rom = 26;
		6234: rom = 27;
		6235: rom = 27;
		6236: rom = 27;
		6237: rom = 27;
		6238: rom = 27;
		6239: rom = 27;
		6240: rom = 27;
		6241: rom = 27;
		6242: rom = 27;
		6243: rom = 27;
		6244: rom = 27;
		6245: rom = 27;
		6246: rom = 27;
		6247: rom = 27;
		6248: rom = 27;
		6249: rom = 27;
		6250: rom = 27;
		6251: rom = 27;
		6252: rom = 27;
		6253: rom = 27;
		6254: rom = 27;
		6255: rom = 27;
		6256: rom = 27;
		6257: rom = 27;
		6258: rom = 27;
		6259: rom = 27;
		6260: rom = 27;
		6261: rom = 27;
		6262: rom = 27;
		6263: rom = 27;
		6264: rom = 27;
		6265: rom = 27;
		6266: rom = 27;
		6272: rom = 27;
		6273: rom = 27;
		6274: rom = 27;
		6275: rom = 27;
		6276: rom = 27;
		6277: rom = 27;
		6278: rom = 27;
		6279: rom = 27;
		6280: rom = 27;
		6281: rom = 27;
		6282: rom = 27;
		6283: rom = 27;
		6284: rom = 27;
		6285: rom = 27;
		6286: rom = 25;
		6287: rom = 12;
		6288: rom = 16;
		6289: rom = 18;
		6290: rom = 18;
		6291: rom = 18;
		6292: rom = 15;
		6293: rom = 9;
		6294: rom = 10;
		6295: rom = 10;
		6296: rom = 19;
		6297: rom = 24;
		6298: rom = 23;
		6299: rom = 21;
		6300: rom = 21;
		6301: rom = 19;
		6302: rom = 18;
		6303: rom = 16;
		6304: rom = 14;
		6305: rom = 7;
		6306: rom = 6;
		6307: rom = 10;
		6308: rom = 18;
		6309: rom = 18;
		6310: rom = 18;
		6311: rom = 18;
		6312: rom = 18;
		6313: rom = 18;
		6314: rom = 11;
		6315: rom = 18;
		6316: rom = 13;
		6317: rom = 18;
		6318: rom = 18;
		6319: rom = 18;
		6320: rom = 18;
		6321: rom = 18;
		6322: rom = 18;
		6323: rom = 14;
		6324: rom = 18;
		6325: rom = 18;
		6326: rom = 18;
		6327: rom = 16;
		6328: rom = 14;
		6329: rom = 18;
		6330: rom = 18;
		6331: rom = 18;
		6332: rom = 23;
		6333: rom = 25;
		6334: rom = 21;
		6335: rom = 18;
		6336: rom = 18;
		6337: rom = 18;
		6338: rom = 21;
		6339: rom = 24;
		6340: rom = 23;
		6341: rom = 16;
		6342: rom = 24;
		6343: rom = 24;
		6344: rom = 24;
		6345: rom = 16;
		6346: rom = 22;
		6347: rom = 24;
		6348: rom = 24;
		6349: rom = 24;
		6350: rom = 24;
		6351: rom = 24;
		6352: rom = 16;
		6353: rom = 26;
		6354: rom = 19;
		6355: rom = 0;
		6356: rom = 0;
		6357: rom = 0;
		6358: rom = 0;
		6359: rom = 0;
		6360: rom = 0;
		6361: rom = 15;
		6362: rom = 27;
		6363: rom = 27;
		6364: rom = 27;
		6365: rom = 27;
		6366: rom = 27;
		6367: rom = 27;
		6368: rom = 27;
		6369: rom = 27;
		6370: rom = 27;
		6371: rom = 27;
		6372: rom = 27;
		6373: rom = 27;
		6374: rom = 27;
		6375: rom = 27;
		6376: rom = 27;
		6377: rom = 27;
		6378: rom = 27;
		6379: rom = 27;
		6380: rom = 27;
		6381: rom = 27;
		6382: rom = 27;
		6383: rom = 27;
		6384: rom = 27;
		6385: rom = 27;
		6386: rom = 27;
		6387: rom = 27;
		6388: rom = 27;
		6389: rom = 27;
		6390: rom = 27;
		6391: rom = 27;
		6392: rom = 27;
		6393: rom = 27;
		6394: rom = 27;
		6400: rom = 27;
		6401: rom = 27;
		6402: rom = 27;
		6403: rom = 27;
		6404: rom = 27;
		6405: rom = 27;
		6406: rom = 27;
		6407: rom = 27;
		6408: rom = 27;
		6409: rom = 27;
		6410: rom = 27;
		6411: rom = 27;
		6412: rom = 27;
		6413: rom = 27;
		6414: rom = 27;
		6415: rom = 26;
		6416: rom = 14;
		6417: rom = 15;
		6418: rom = 18;
		6419: rom = 18;
		6420: rom = 11;
		6421: rom = 20;
		6422: rom = 14;
		6423: rom = 15;
		6424: rom = 12;
		6425: rom = 15;
		6426: rom = 9;
		6427: rom = 12;
		6428: rom = 13;
		6429: rom = 14;
		6430: rom = 15;
		6431: rom = 16;
		6432: rom = 17;
		6433: rom = 17;
		6434: rom = 17;
		6435: rom = 25;
		6436: rom = 24;
		6437: rom = 18;
		6438: rom = 18;
		6439: rom = 18;
		6440: rom = 18;
		6441: rom = 18;
		6442: rom = 11;
		6443: rom = 18;
		6444: rom = 10;
		6445: rom = 18;
		6446: rom = 18;
		6447: rom = 18;
		6448: rom = 18;
		6449: rom = 18;
		6450: rom = 18;
		6451: rom = 17;
		6452: rom = 18;
		6453: rom = 18;
		6454: rom = 18;
		6455: rom = 18;
		6456: rom = 10;
		6457: rom = 18;
		6458: rom = 18;
		6459: rom = 18;
		6460: rom = 19;
		6461: rom = 25;
		6462: rom = 25;
		6463: rom = 19;
		6464: rom = 18;
		6465: rom = 18;
		6466: rom = 19;
		6467: rom = 24;
		6468: rom = 21;
		6469: rom = 18;
		6470: rom = 24;
		6471: rom = 24;
		6472: rom = 23;
		6473: rom = 14;
		6474: rom = 24;
		6475: rom = 24;
		6476: rom = 24;
		6477: rom = 24;
		6478: rom = 24;
		6479: rom = 24;
		6480: rom = 15;
		6481: rom = 27;
		6482: rom = 19;
		6483: rom = 0;
		6484: rom = 0;
		6485: rom = 0;
		6486: rom = 0;
		6487: rom = 0;
		6488: rom = 0;
		6489: rom = 24;
		6490: rom = 27;
		6491: rom = 27;
		6492: rom = 27;
		6493: rom = 27;
		6494: rom = 27;
		6495: rom = 27;
		6496: rom = 27;
		6497: rom = 27;
		6498: rom = 27;
		6499: rom = 27;
		6500: rom = 27;
		6501: rom = 27;
		6502: rom = 27;
		6503: rom = 27;
		6504: rom = 27;
		6505: rom = 27;
		6506: rom = 27;
		6507: rom = 27;
		6508: rom = 27;
		6509: rom = 27;
		6510: rom = 27;
		6511: rom = 27;
		6512: rom = 27;
		6513: rom = 27;
		6514: rom = 27;
		6515: rom = 27;
		6516: rom = 27;
		6517: rom = 27;
		6518: rom = 27;
		6519: rom = 27;
		6520: rom = 27;
		6521: rom = 27;
		6522: rom = 27;
		6528: rom = 27;
		6529: rom = 27;
		6530: rom = 27;
		6531: rom = 27;
		6532: rom = 16;
		6533: rom = 25;
		6534: rom = 27;
		6535: rom = 27;
		6536: rom = 27;
		6537: rom = 27;
		6538: rom = 27;
		6539: rom = 27;
		6540: rom = 27;
		6541: rom = 27;
		6542: rom = 27;
		6543: rom = 27;
		6544: rom = 27;
		6545: rom = 12;
		6546: rom = 10;
		6547: rom = 13;
		6548: rom = 12;
		6549: rom = 17;
		6550: rom = 18;
		6551: rom = 13;
		6552: rom = 17;
		6553: rom = 11;
		6554: rom = 17;
		6555: rom = 18;
		6556: rom = 18;
		6557: rom = 18;
		6558: rom = 18;
		6559: rom = 18;
		6560: rom = 18;
		6561: rom = 18;
		6562: rom = 18;
		6563: rom = 25;
		6564: rom = 24;
		6565: rom = 18;
		6566: rom = 18;
		6567: rom = 18;
		6568: rom = 18;
		6569: rom = 18;
		6570: rom = 15;
		6571: rom = 15;
		6572: rom = 11;
		6573: rom = 18;
		6574: rom = 18;
		6575: rom = 18;
		6576: rom = 18;
		6577: rom = 18;
		6578: rom = 18;
		6579: rom = 18;
		6580: rom = 18;
		6581: rom = 18;
		6582: rom = 18;
		6583: rom = 18;
		6584: rom = 14;
		6585: rom = 16;
		6586: rom = 18;
		6587: rom = 18;
		6588: rom = 18;
		6589: rom = 21;
		6590: rom = 25;
		6591: rom = 24;
		6592: rom = 19;
		6593: rom = 18;
		6594: rom = 18;
		6595: rom = 23;
		6596: rom = 20;
		6597: rom = 20;
		6598: rom = 24;
		6599: rom = 24;
		6600: rom = 21;
		6601: rom = 18;
		6602: rom = 24;
		6603: rom = 24;
		6604: rom = 24;
		6605: rom = 24;
		6606: rom = 24;
		6607: rom = 23;
		6608: rom = 17;
		6609: rom = 27;
		6610: rom = 25;
		6611: rom = 23;
		6612: rom = 23;
		6613: rom = 23;
		6614: rom = 23;
		6615: rom = 23;
		6616: rom = 24;
		6617: rom = 27;
		6618: rom = 27;
		6619: rom = 27;
		6620: rom = 27;
		6621: rom = 27;
		6622: rom = 27;
		6623: rom = 27;
		6624: rom = 27;
		6625: rom = 27;
		6626: rom = 27;
		6627: rom = 27;
		6628: rom = 27;
		6629: rom = 27;
		6630: rom = 27;
		6631: rom = 27;
		6632: rom = 27;
		6633: rom = 27;
		6634: rom = 27;
		6635: rom = 27;
		6636: rom = 27;
		6637: rom = 27;
		6638: rom = 27;
		6639: rom = 27;
		6640: rom = 27;
		6641: rom = 27;
		6642: rom = 27;
		6643: rom = 27;
		6644: rom = 27;
		6645: rom = 27;
		6646: rom = 27;
		6647: rom = 27;
		6648: rom = 27;
		6649: rom = 27;
		6650: rom = 27;
		6656: rom = 27;
		6657: rom = 27;
		6658: rom = 27;
		6659: rom = 27;
		6660: rom = 0;
		6661: rom = 0;
		6662: rom = 27;
		6663: rom = 27;
		6664: rom = 27;
		6665: rom = 27;
		6666: rom = 27;
		6667: rom = 27;
		6668: rom = 27;
		6669: rom = 27;
		6670: rom = 27;
		6671: rom = 27;
		6672: rom = 27;
		6673: rom = 11;
		6674: rom = 19;
		6675: rom = 17;
		6676: rom = 9;
		6677: rom = 8;
		6678: rom = 17;
		6679: rom = 10;
		6680: rom = 10;
		6681: rom = 12;
		6682: rom = 13;
		6683: rom = 18;
		6684: rom = 18;
		6685: rom = 18;
		6686: rom = 18;
		6687: rom = 18;
		6688: rom = 18;
		6689: rom = 18;
		6690: rom = 18;
		6691: rom = 24;
		6692: rom = 24;
		6693: rom = 18;
		6694: rom = 18;
		6695: rom = 18;
		6696: rom = 18;
		6697: rom = 18;
		6698: rom = 17;
		6699: rom = 13;
		6700: rom = 12;
		6701: rom = 18;
		6702: rom = 18;
		6703: rom = 18;
		6704: rom = 18;
		6705: rom = 18;
		6706: rom = 18;
		6707: rom = 18;
		6708: rom = 18;
		6709: rom = 13;
		6710: rom = 18;
		6711: rom = 18;
		6712: rom = 18;
		6713: rom = 11;
		6714: rom = 18;
		6715: rom = 18;
		6716: rom = 18;
		6717: rom = 18;
		6718: rom = 23;
		6719: rom = 25;
		6720: rom = 24;
		6721: rom = 19;
		6722: rom = 18;
		6723: rom = 21;
		6724: rom = 18;
		6725: rom = 21;
		6726: rom = 24;
		6727: rom = 24;
		6728: rom = 16;
		6729: rom = 22;
		6730: rom = 24;
		6731: rom = 24;
		6732: rom = 24;
		6733: rom = 24;
		6734: rom = 24;
		6735: rom = 21;
		6736: rom = 21;
		6737: rom = 27;
		6738: rom = 27;
		6739: rom = 27;
		6740: rom = 27;
		6741: rom = 27;
		6742: rom = 27;
		6743: rom = 27;
		6744: rom = 27;
		6745: rom = 27;
		6746: rom = 27;
		6747: rom = 27;
		6748: rom = 27;
		6749: rom = 27;
		6750: rom = 27;
		6751: rom = 27;
		6752: rom = 27;
		6753: rom = 27;
		6754: rom = 27;
		6755: rom = 27;
		6756: rom = 27;
		6757: rom = 27;
		6758: rom = 27;
		6759: rom = 27;
		6760: rom = 27;
		6761: rom = 27;
		6762: rom = 27;
		6763: rom = 27;
		6764: rom = 27;
		6765: rom = 27;
		6766: rom = 27;
		6767: rom = 27;
		6768: rom = 27;
		6769: rom = 27;
		6770: rom = 27;
		6771: rom = 27;
		6772: rom = 27;
		6773: rom = 27;
		6774: rom = 27;
		6775: rom = 27;
		6776: rom = 27;
		6777: rom = 27;
		6778: rom = 27;
		6784: rom = 27;
		6785: rom = 27;
		6786: rom = 27;
		6787: rom = 27;
		6788: rom = 0;
		6789: rom = 0;
		6790: rom = 27;
		6791: rom = 27;
		6792: rom = 27;
		6793: rom = 27;
		6794: rom = 27;
		6795: rom = 27;
		6796: rom = 27;
		6797: rom = 27;
		6798: rom = 27;
		6799: rom = 27;
		6800: rom = 27;
		6801: rom = 19;
		6802: rom = 16;
		6803: rom = 20;
		6804: rom = 20;
		6805: rom = 12;
		6806: rom = 7;
		6807: rom = 13;
		6808: rom = 20;
		6809: rom = 15;
		6810: rom = 15;
		6811: rom = 18;
		6812: rom = 18;
		6813: rom = 18;
		6814: rom = 18;
		6815: rom = 18;
		6816: rom = 18;
		6817: rom = 18;
		6818: rom = 18;
		6819: rom = 24;
		6820: rom = 24;
		6821: rom = 18;
		6822: rom = 18;
		6823: rom = 18;
		6824: rom = 18;
		6825: rom = 18;
		6826: rom = 18;
		6827: rom = 11;
		6828: rom = 12;
		6829: rom = 18;
		6830: rom = 18;
		6831: rom = 18;
		6832: rom = 18;
		6833: rom = 18;
		6834: rom = 18;
		6835: rom = 18;
		6836: rom = 18;
		6837: rom = 12;
		6838: rom = 18;
		6839: rom = 18;
		6840: rom = 18;
		6841: rom = 12;
		6842: rom = 17;
		6843: rom = 18;
		6844: rom = 18;
		6845: rom = 18;
		6846: rom = 18;
		6847: rom = 23;
		6848: rom = 25;
		6849: rom = 25;
		6850: rom = 21;
		6851: rom = 20;
		6852: rom = 17;
		6853: rom = 22;
		6854: rom = 24;
		6855: rom = 23;
		6856: rom = 14;
		6857: rom = 24;
		6858: rom = 24;
		6859: rom = 24;
		6860: rom = 24;
		6861: rom = 24;
		6862: rom = 24;
		6863: rom = 18;
		6864: rom = 10;
		6865: rom = 10;
		6866: rom = 10;
		6867: rom = 10;
		6868: rom = 10;
		6869: rom = 11;
		6870: rom = 12;
		6871: rom = 15;
		6872: rom = 17;
		6873: rom = 19;
		6874: rom = 23;
		6875: rom = 24;
		6876: rom = 27;
		6877: rom = 27;
		6878: rom = 27;
		6879: rom = 27;
		6880: rom = 27;
		6881: rom = 27;
		6882: rom = 27;
		6883: rom = 27;
		6884: rom = 27;
		6885: rom = 27;
		6886: rom = 27;
		6887: rom = 27;
		6888: rom = 27;
		6889: rom = 27;
		6890: rom = 27;
		6891: rom = 27;
		6892: rom = 27;
		6893: rom = 27;
		6894: rom = 27;
		6895: rom = 27;
		6896: rom = 27;
		6897: rom = 27;
		6898: rom = 27;
		6899: rom = 27;
		6900: rom = 27;
		6901: rom = 27;
		6902: rom = 27;
		6903: rom = 27;
		6904: rom = 27;
		6905: rom = 27;
		6906: rom = 27;
		6912: rom = 27;
		6913: rom = 27;
		6914: rom = 27;
		6915: rom = 27;
		6916: rom = 0;
		6917: rom = 0;
		6918: rom = 27;
		6919: rom = 27;
		6920: rom = 27;
		6921: rom = 27;
		6922: rom = 27;
		6923: rom = 27;
		6924: rom = 27;
		6925: rom = 27;
		6926: rom = 27;
		6927: rom = 27;
		6928: rom = 27;
		6929: rom = 27;
		6930: rom = 20;
		6931: rom = 14;
		6932: rom = 10;
		6933: rom = 5;
		6934: rom = 0;
		6935: rom = 12;
		6936: rom = 12;
		6937: rom = 8;
		6938: rom = 14;
		6939: rom = 16;
		6940: rom = 17;
		6941: rom = 18;
		6942: rom = 18;
		6943: rom = 18;
		6944: rom = 18;
		6945: rom = 18;
		6946: rom = 18;
		6947: rom = 24;
		6948: rom = 24;
		6949: rom = 18;
		6950: rom = 18;
		6951: rom = 18;
		6952: rom = 18;
		6953: rom = 18;
		6954: rom = 18;
		6955: rom = 11;
		6956: rom = 14;
		6957: rom = 12;
		6958: rom = 17;
		6959: rom = 18;
		6960: rom = 18;
		6961: rom = 18;
		6962: rom = 18;
		6963: rom = 17;
		6964: rom = 18;
		6965: rom = 14;
		6966: rom = 18;
		6967: rom = 18;
		6968: rom = 18;
		6969: rom = 17;
		6970: rom = 11;
		6971: rom = 18;
		6972: rom = 18;
		6973: rom = 18;
		6974: rom = 18;
		6975: rom = 18;
		6976: rom = 22;
		6977: rom = 25;
		6978: rom = 25;
		6979: rom = 24;
		6980: rom = 17;
		6981: rom = 23;
		6982: rom = 24;
		6983: rom = 21;
		6984: rom = 18;
		6985: rom = 24;
		6986: rom = 24;
		6987: rom = 24;
		6988: rom = 24;
		6989: rom = 24;
		6990: rom = 24;
		6991: rom = 14;
		6992: rom = 17;
		6993: rom = 18;
		6994: rom = 18;
		6995: rom = 18;
		6996: rom = 18;
		6997: rom = 18;
		6998: rom = 18;
		6999: rom = 17;
		7000: rom = 17;
		7001: rom = 16;
		7002: rom = 14;
		7003: rom = 12;
		7004: rom = 10;
		7005: rom = 13;
		7006: rom = 18;
		7007: rom = 22;
		7008: rom = 25;
		7009: rom = 27;
		7010: rom = 27;
		7011: rom = 27;
		7012: rom = 27;
		7013: rom = 27;
		7014: rom = 27;
		7015: rom = 27;
		7016: rom = 27;
		7017: rom = 27;
		7018: rom = 27;
		7019: rom = 27;
		7020: rom = 27;
		7021: rom = 27;
		7022: rom = 27;
		7023: rom = 27;
		7024: rom = 27;
		7025: rom = 27;
		7026: rom = 27;
		7027: rom = 27;
		7028: rom = 27;
		7029: rom = 27;
		7030: rom = 27;
		7031: rom = 27;
		7032: rom = 27;
		7033: rom = 27;
		7034: rom = 27;
		7040: rom = 27;
		7041: rom = 27;
		7042: rom = 27;
		7043: rom = 27;
		7044: rom = 0;
		7045: rom = 0;
		7046: rom = 27;
		7047: rom = 27;
		7048: rom = 27;
		7049: rom = 27;
		7050: rom = 27;
		7051: rom = 27;
		7052: rom = 27;
		7053: rom = 27;
		7054: rom = 27;
		7055: rom = 27;
		7056: rom = 27;
		7057: rom = 27;
		7058: rom = 27;
		7059: rom = 23;
		7060: rom = 12;
		7061: rom = 9;
		7062: rom = 9;
		7063: rom = 8;
		7064: rom = 11;
		7065: rom = 3;
		7066: rom = 4;
		7067: rom = 7;
		7068: rom = 9;
		7069: rom = 12;
		7070: rom = 17;
		7071: rom = 18;
		7072: rom = 18;
		7073: rom = 18;
		7074: rom = 18;
		7075: rom = 24;
		7076: rom = 24;
		7077: rom = 18;
		7078: rom = 18;
		7079: rom = 18;
		7080: rom = 18;
		7081: rom = 18;
		7082: rom = 18;
		7083: rom = 12;
		7084: rom = 17;
		7085: rom = 26;
		7086: rom = 11;
		7087: rom = 18;
		7088: rom = 18;
		7089: rom = 13;
		7090: rom = 13;
		7091: rom = 20;
		7092: rom = 19;
		7093: rom = 16;
		7094: rom = 18;
		7095: rom = 18;
		7096: rom = 18;
		7097: rom = 18;
		7098: rom = 13;
		7099: rom = 16;
		7100: rom = 18;
		7101: rom = 18;
		7102: rom = 18;
		7103: rom = 18;
		7104: rom = 18;
		7105: rom = 20;
		7106: rom = 24;
		7107: rom = 25;
		7108: rom = 17;
		7109: rom = 23;
		7110: rom = 24;
		7111: rom = 17;
		7112: rom = 22;
		7113: rom = 24;
		7114: rom = 24;
		7115: rom = 24;
		7116: rom = 24;
		7117: rom = 24;
		7118: rom = 24;
		7119: rom = 11;
		7120: rom = 18;
		7121: rom = 18;
		7122: rom = 18;
		7123: rom = 18;
		7124: rom = 18;
		7125: rom = 18;
		7126: rom = 18;
		7127: rom = 18;
		7128: rom = 18;
		7129: rom = 18;
		7130: rom = 18;
		7131: rom = 18;
		7132: rom = 18;
		7133: rom = 18;
		7134: rom = 16;
		7135: rom = 14;
		7136: rom = 11;
		7137: rom = 12;
		7138: rom = 18;
		7139: rom = 24;
		7140: rom = 27;
		7141: rom = 27;
		7142: rom = 27;
		7143: rom = 27;
		7144: rom = 27;
		7145: rom = 27;
		7146: rom = 27;
		7147: rom = 27;
		7148: rom = 27;
		7149: rom = 27;
		7150: rom = 27;
		7151: rom = 27;
		7152: rom = 27;
		7153: rom = 27;
		7154: rom = 27;
		7155: rom = 27;
		7156: rom = 27;
		7157: rom = 27;
		7158: rom = 27;
		7159: rom = 27;
		7160: rom = 27;
		7161: rom = 27;
		7162: rom = 27;
		7168: rom = 27;
		7169: rom = 27;
		7170: rom = 27;
		7171: rom = 27;
		7172: rom = 0;
		7173: rom = 0;
		7174: rom = 0;
		7175: rom = 0;
		7176: rom = 0;
		7177: rom = 0;
		7178: rom = 0;
		7179: rom = 0;
		7180: rom = 0;
		7181: rom = 0;
		7182: rom = 0;
		7183: rom = 16;
		7184: rom = 27;
		7185: rom = 27;
		7186: rom = 27;
		7187: rom = 17;
		7188: rom = 16;
		7189: rom = 9;
		7190: rom = 8;
		7191: rom = 18;
		7192: rom = 9;
		7193: rom = 8;
		7194: rom = 6;
		7195: rom = 5;
		7196: rom = 19;
		7197: rom = 19;
		7198: rom = 10;
		7199: rom = 16;
		7200: rom = 18;
		7201: rom = 18;
		7202: rom = 18;
		7203: rom = 25;
		7204: rom = 24;
		7205: rom = 18;
		7206: rom = 18;
		7207: rom = 18;
		7208: rom = 18;
		7209: rom = 18;
		7210: rom = 15;
		7211: rom = 15;
		7212: rom = 18;
		7213: rom = 27;
		7214: rom = 15;
		7215: rom = 15;
		7216: rom = 18;
		7217: rom = 12;
		7218: rom = 23;
		7219: rom = 24;
		7220: rom = 17;
		7221: rom = 17;
		7222: rom = 18;
		7223: rom = 18;
		7224: rom = 18;
		7225: rom = 18;
		7226: rom = 18;
		7227: rom = 10;
		7228: rom = 18;
		7229: rom = 18;
		7230: rom = 18;
		7231: rom = 18;
		7232: rom = 18;
		7233: rom = 18;
		7234: rom = 19;
		7235: rom = 22;
		7236: rom = 22;
		7237: rom = 24;
		7238: rom = 24;
		7239: rom = 14;
		7240: rom = 24;
		7241: rom = 24;
		7242: rom = 24;
		7243: rom = 24;
		7244: rom = 24;
		7245: rom = 24;
		7246: rom = 21;
		7247: rom = 13;
		7248: rom = 18;
		7249: rom = 18;
		7250: rom = 18;
		7251: rom = 18;
		7252: rom = 18;
		7253: rom = 18;
		7254: rom = 18;
		7255: rom = 18;
		7256: rom = 18;
		7257: rom = 18;
		7258: rom = 18;
		7259: rom = 18;
		7260: rom = 18;
		7261: rom = 18;
		7262: rom = 18;
		7263: rom = 18;
		7264: rom = 18;
		7265: rom = 18;
		7266: rom = 16;
		7267: rom = 13;
		7268: rom = 10;
		7269: rom = 18;
		7270: rom = 25;
		7271: rom = 27;
		7272: rom = 27;
		7273: rom = 27;
		7274: rom = 27;
		7275: rom = 27;
		7276: rom = 27;
		7277: rom = 27;
		7278: rom = 27;
		7279: rom = 27;
		7280: rom = 27;
		7281: rom = 27;
		7282: rom = 27;
		7283: rom = 27;
		7284: rom = 27;
		7285: rom = 27;
		7286: rom = 27;
		7287: rom = 27;
		7288: rom = 27;
		7289: rom = 27;
		7290: rom = 27;
		7296: rom = 27;
		7297: rom = 27;
		7298: rom = 27;
		7299: rom = 27;
		7300: rom = 0;
		7301: rom = 0;
		7302: rom = 0;
		7303: rom = 0;
		7304: rom = 0;
		7305: rom = 0;
		7306: rom = 0;
		7307: rom = 0;
		7308: rom = 0;
		7309: rom = 0;
		7310: rom = 0;
		7311: rom = 16;
		7312: rom = 27;
		7313: rom = 27;
		7314: rom = 27;
		7315: rom = 24;
		7316: rom = 9;
		7317: rom = 22;
		7318: rom = 16;
		7319: rom = 20;
		7320: rom = 10;
		7321: rom = 10;
		7322: rom = 6;
		7323: rom = 4;
		7324: rom = 4;
		7325: rom = 17;
		7326: rom = 22;
		7327: rom = 12;
		7328: rom = 18;
		7329: rom = 18;
		7330: rom = 18;
		7331: rom = 25;
		7332: rom = 24;
		7333: rom = 18;
		7334: rom = 18;
		7335: rom = 18;
		7336: rom = 18;
		7337: rom = 18;
		7338: rom = 11;
		7339: rom = 17;
		7340: rom = 20;
		7341: rom = 27;
		7342: rom = 15;
		7343: rom = 17;
		7344: rom = 18;
		7345: rom = 14;
		7346: rom = 13;
		7347: rom = 20;
		7348: rom = 16;
		7349: rom = 17;
		7350: rom = 18;
		7351: rom = 18;
		7352: rom = 18;
		7353: rom = 18;
		7354: rom = 18;
		7355: rom = 15;
		7356: rom = 13;
		7357: rom = 18;
		7358: rom = 18;
		7359: rom = 18;
		7360: rom = 18;
		7361: rom = 18;
		7362: rom = 18;
		7363: rom = 18;
		7364: rom = 19;
		7365: rom = 23;
		7366: rom = 22;
		7367: rom = 16;
		7368: rom = 24;
		7369: rom = 24;
		7370: rom = 24;
		7371: rom = 24;
		7372: rom = 24;
		7373: rom = 24;
		7374: rom = 17;
		7375: rom = 16;
		7376: rom = 18;
		7377: rom = 18;
		7378: rom = 18;
		7379: rom = 18;
		7380: rom = 18;
		7381: rom = 18;
		7382: rom = 18;
		7383: rom = 18;
		7384: rom = 18;
		7385: rom = 18;
		7386: rom = 18;
		7387: rom = 18;
		7388: rom = 18;
		7389: rom = 18;
		7390: rom = 18;
		7391: rom = 18;
		7392: rom = 18;
		7393: rom = 18;
		7394: rom = 18;
		7395: rom = 18;
		7396: rom = 18;
		7397: rom = 15;
		7398: rom = 10;
		7399: rom = 15;
		7400: rom = 25;
		7401: rom = 27;
		7402: rom = 27;
		7403: rom = 27;
		7404: rom = 27;
		7405: rom = 27;
		7406: rom = 27;
		7407: rom = 27;
		7408: rom = 27;
		7409: rom = 27;
		7410: rom = 27;
		7411: rom = 27;
		7412: rom = 27;
		7413: rom = 27;
		7414: rom = 27;
		7415: rom = 27;
		7416: rom = 27;
		7417: rom = 27;
		7418: rom = 27;
		7424: rom = 27;
		7425: rom = 27;
		7426: rom = 27;
		7427: rom = 27;
		7428: rom = 0;
		7429: rom = 0;
		7430: rom = 20;
		7431: rom = 20;
		7432: rom = 20;
		7433: rom = 20;
		7434: rom = 20;
		7435: rom = 20;
		7436: rom = 20;
		7437: rom = 20;
		7438: rom = 20;
		7439: rom = 20;
		7440: rom = 27;
		7441: rom = 27;
		7442: rom = 27;
		7443: rom = 27;
		7444: rom = 17;
		7445: rom = 25;
		7446: rom = 16;
		7447: rom = 15;
		7448: rom = 21;
		7449: rom = 21;
		7450: rom = 2;
		7451: rom = 12;
		7452: rom = 4;
		7453: rom = 4;
		7454: rom = 9;
		7455: rom = 9;
		7456: rom = 24;
		7457: rom = 21;
		7458: rom = 20;
		7459: rom = 25;
		7460: rom = 23;
		7461: rom = 18;
		7462: rom = 18;
		7463: rom = 18;
		7464: rom = 18;
		7465: rom = 16;
		7466: rom = 12;
		7467: rom = 16;
		7468: rom = 24;
		7469: rom = 26;
		7470: rom = 11;
		7471: rom = 18;
		7472: rom = 13;
		7473: rom = 15;
		7474: rom = 21;
		7475: rom = 22;
		7476: rom = 17;
		7477: rom = 17;
		7478: rom = 18;
		7479: rom = 18;
		7480: rom = 18;
		7481: rom = 18;
		7482: rom = 18;
		7483: rom = 18;
		7484: rom = 10;
		7485: rom = 15;
		7486: rom = 18;
		7487: rom = 18;
		7488: rom = 18;
		7489: rom = 18;
		7490: rom = 18;
		7491: rom = 18;
		7492: rom = 18;
		7493: rom = 23;
		7494: rom = 19;
		7495: rom = 20;
		7496: rom = 24;
		7497: rom = 24;
		7498: rom = 24;
		7499: rom = 24;
		7500: rom = 24;
		7501: rom = 24;
		7502: rom = 13;
		7503: rom = 18;
		7504: rom = 18;
		7505: rom = 18;
		7506: rom = 18;
		7507: rom = 18;
		7508: rom = 18;
		7509: rom = 18;
		7510: rom = 18;
		7511: rom = 18;
		7512: rom = 18;
		7513: rom = 18;
		7514: rom = 18;
		7515: rom = 18;
		7516: rom = 18;
		7517: rom = 18;
		7518: rom = 18;
		7519: rom = 18;
		7520: rom = 18;
		7521: rom = 18;
		7522: rom = 18;
		7523: rom = 18;
		7524: rom = 18;
		7525: rom = 18;
		7526: rom = 18;
		7527: rom = 18;
		7528: rom = 14;
		7529: rom = 20;
		7530: rom = 27;
		7531: rom = 27;
		7532: rom = 27;
		7533: rom = 27;
		7534: rom = 27;
		7535: rom = 27;
		7536: rom = 27;
		7537: rom = 27;
		7538: rom = 27;
		7539: rom = 27;
		7540: rom = 27;
		7541: rom = 27;
		7542: rom = 27;
		7543: rom = 27;
		7544: rom = 27;
		7545: rom = 27;
		7546: rom = 27;
		7552: rom = 27;
		7553: rom = 27;
		7554: rom = 27;
		7555: rom = 27;
		7556: rom = 0;
		7557: rom = 0;
		7558: rom = 27;
		7559: rom = 27;
		7560: rom = 27;
		7561: rom = 27;
		7562: rom = 27;
		7563: rom = 27;
		7564: rom = 27;
		7565: rom = 27;
		7566: rom = 27;
		7567: rom = 27;
		7568: rom = 27;
		7569: rom = 27;
		7570: rom = 27;
		7571: rom = 27;
		7572: rom = 21;
		7573: rom = 22;
		7574: rom = 24;
		7575: rom = 21;
		7576: rom = 23;
		7577: rom = 10;
		7578: rom = 16;
		7579: rom = 18;
		7580: rom = 16;
		7581: rom = 6;
		7582: rom = 8;
		7583: rom = 12;
		7584: rom = 23;
		7585: rom = 25;
		7586: rom = 25;
		7587: rom = 25;
		7588: rom = 22;
		7589: rom = 18;
		7590: rom = 18;
		7591: rom = 18;
		7592: rom = 17;
		7593: rom = 9;
		7594: rom = 18;
		7595: rom = 13;
		7596: rom = 27;
		7597: rom = 19;
		7598: rom = 17;
		7599: rom = 13;
		7600: rom = 18;
		7601: rom = 24;
		7602: rom = 24;
		7603: rom = 24;
		7604: rom = 18;
		7605: rom = 16;
		7606: rom = 18;
		7607: rom = 18;
		7608: rom = 18;
		7609: rom = 18;
		7610: rom = 18;
		7611: rom = 18;
		7612: rom = 15;
		7613: rom = 4;
		7614: rom = 16;
		7615: rom = 18;
		7616: rom = 18;
		7617: rom = 18;
		7618: rom = 18;
		7619: rom = 18;
		7620: rom = 18;
		7621: rom = 22;
		7622: rom = 15;
		7623: rom = 23;
		7624: rom = 24;
		7625: rom = 24;
		7626: rom = 24;
		7627: rom = 24;
		7628: rom = 24;
		7629: rom = 23;
		7630: rom = 16;
		7631: rom = 20;
		7632: rom = 18;
		7633: rom = 18;
		7634: rom = 18;
		7635: rom = 18;
		7636: rom = 18;
		7637: rom = 18;
		7638: rom = 18;
		7639: rom = 18;
		7640: rom = 18;
		7641: rom = 18;
		7642: rom = 18;
		7643: rom = 18;
		7644: rom = 18;
		7645: rom = 18;
		7646: rom = 18;
		7647: rom = 18;
		7648: rom = 18;
		7649: rom = 18;
		7650: rom = 18;
		7651: rom = 18;
		7652: rom = 18;
		7653: rom = 18;
		7654: rom = 18;
		7655: rom = 22;
		7656: rom = 25;
		7657: rom = 20;
		7658: rom = 15;
		7659: rom = 27;
		7660: rom = 27;
		7661: rom = 27;
		7662: rom = 27;
		7663: rom = 27;
		7664: rom = 27;
		7665: rom = 27;
		7666: rom = 27;
		7667: rom = 27;
		7668: rom = 27;
		7669: rom = 27;
		7670: rom = 27;
		7671: rom = 27;
		7672: rom = 27;
		7673: rom = 27;
		7674: rom = 27;
		7680: rom = 27;
		7681: rom = 27;
		7682: rom = 27;
		7683: rom = 27;
		7684: rom = 0;
		7685: rom = 0;
		7686: rom = 27;
		7687: rom = 27;
		7688: rom = 27;
		7689: rom = 27;
		7690: rom = 27;
		7691: rom = 27;
		7692: rom = 27;
		7693: rom = 27;
		7694: rom = 27;
		7695: rom = 27;
		7696: rom = 27;
		7697: rom = 27;
		7698: rom = 27;
		7699: rom = 27;
		7700: rom = 27;
		7701: rom = 27;
		7702: rom = 27;
		7703: rom = 27;
		7704: rom = 11;
		7705: rom = 18;
		7706: rom = 18;
		7707: rom = 18;
		7708: rom = 18;
		7709: rom = 17;
		7710: rom = 17;
		7711: rom = 17;
		7712: rom = 16;
		7713: rom = 23;
		7714: rom = 24;
		7715: rom = 23;
		7716: rom = 19;
		7717: rom = 18;
		7718: rom = 18;
		7719: rom = 18;
		7720: rom = 9;
		7721: rom = 17;
		7722: rom = 17;
		7723: rom = 19;
		7724: rom = 27;
		7725: rom = 14;
		7726: rom = 21;
		7727: rom = 11;
		7728: rom = 23;
		7729: rom = 24;
		7730: rom = 24;
		7731: rom = 18;
		7732: rom = 20;
		7733: rom = 14;
		7734: rom = 18;
		7735: rom = 18;
		7736: rom = 18;
		7737: rom = 18;
		7738: rom = 18;
		7739: rom = 18;
		7740: rom = 18;
		7741: rom = 10;
		7742: rom = 13;
		7743: rom = 15;
		7744: rom = 18;
		7745: rom = 18;
		7746: rom = 18;
		7747: rom = 18;
		7748: rom = 18;
		7749: rom = 20;
		7750: rom = 14;
		7751: rom = 24;
		7752: rom = 24;
		7753: rom = 24;
		7754: rom = 24;
		7755: rom = 24;
		7756: rom = 24;
		7757: rom = 19;
		7758: rom = 21;
		7759: rom = 25;
		7760: rom = 22;
		7761: rom = 18;
		7762: rom = 18;
		7763: rom = 18;
		7764: rom = 18;
		7765: rom = 18;
		7766: rom = 18;
		7767: rom = 18;
		7768: rom = 18;
		7769: rom = 18;
		7770: rom = 18;
		7771: rom = 18;
		7772: rom = 18;
		7773: rom = 18;
		7774: rom = 18;
		7775: rom = 18;
		7776: rom = 18;
		7777: rom = 18;
		7778: rom = 18;
		7779: rom = 18;
		7780: rom = 18;
		7781: rom = 18;
		7782: rom = 18;
		7783: rom = 24;
		7784: rom = 25;
		7785: rom = 25;
		7786: rom = 23;
		7787: rom = 16;
		7788: rom = 27;
		7789: rom = 27;
		7790: rom = 27;
		7791: rom = 27;
		7792: rom = 27;
		7793: rom = 27;
		7794: rom = 27;
		7795: rom = 27;
		7796: rom = 27;
		7797: rom = 27;
		7798: rom = 27;
		7799: rom = 27;
		7800: rom = 27;
		7801: rom = 27;
		7802: rom = 27;
		7808: rom = 27;
		7809: rom = 27;
		7810: rom = 27;
		7811: rom = 27;
		7812: rom = 0;
		7813: rom = 0;
		7814: rom = 27;
		7815: rom = 27;
		7816: rom = 27;
		7817: rom = 27;
		7818: rom = 27;
		7819: rom = 27;
		7820: rom = 27;
		7821: rom = 27;
		7822: rom = 27;
		7823: rom = 27;
		7824: rom = 27;
		7825: rom = 27;
		7826: rom = 27;
		7827: rom = 27;
		7828: rom = 27;
		7829: rom = 27;
		7830: rom = 27;
		7831: rom = 27;
		7832: rom = 11;
		7833: rom = 18;
		7834: rom = 18;
		7835: rom = 18;
		7836: rom = 12;
		7837: rom = 18;
		7838: rom = 15;
		7839: rom = 18;
		7840: rom = 12;
		7841: rom = 18;
		7842: rom = 18;
		7843: rom = 18;
		7844: rom = 18;
		7845: rom = 18;
		7846: rom = 18;
		7847: rom = 15;
		7848: rom = 15;
		7849: rom = 18;
		7850: rom = 12;
		7851: rom = 26;
		7852: rom = 24;
		7853: rom = 19;
		7854: rom = 25;
		7855: rom = 22;
		7856: rom = 12;
		7857: rom = 17;
		7858: rom = 13;
		7859: rom = 13;
		7860: rom = 21;
		7861: rom = 12;
		7862: rom = 18;
		7863: rom = 18;
		7864: rom = 18;
		7865: rom = 18;
		7866: rom = 18;
		7867: rom = 18;
		7868: rom = 18;
		7869: rom = 15;
		7870: rom = 14;
		7871: rom = 18;
		7872: rom = 18;
		7873: rom = 18;
		7874: rom = 18;
		7875: rom = 18;
		7876: rom = 18;
		7877: rom = 19;
		7878: rom = 15;
		7879: rom = 24;
		7880: rom = 24;
		7881: rom = 24;
		7882: rom = 24;
		7883: rom = 24;
		7884: rom = 24;
		7885: rom = 14;
		7886: rom = 21;
		7887: rom = 25;
		7888: rom = 25;
		7889: rom = 20;
		7890: rom = 18;
		7891: rom = 18;
		7892: rom = 18;
		7893: rom = 18;
		7894: rom = 18;
		7895: rom = 18;
		7896: rom = 18;
		7897: rom = 18;
		7898: rom = 18;
		7899: rom = 18;
		7900: rom = 18;
		7901: rom = 18;
		7902: rom = 18;
		7903: rom = 18;
		7904: rom = 18;
		7905: rom = 18;
		7906: rom = 18;
		7907: rom = 18;
		7908: rom = 18;
		7909: rom = 18;
		7910: rom = 18;
		7911: rom = 25;
		7912: rom = 25;
		7913: rom = 25;
		7914: rom = 25;
		7915: rom = 17;
		7916: rom = 23;
		7917: rom = 27;
		7918: rom = 27;
		7919: rom = 27;
		7920: rom = 27;
		7921: rom = 27;
		7922: rom = 27;
		7923: rom = 27;
		7924: rom = 27;
		7925: rom = 27;
		7926: rom = 27;
		7927: rom = 27;
		7928: rom = 27;
		7929: rom = 27;
		7930: rom = 27;
		7936: rom = 27;
		7937: rom = 27;
		7938: rom = 27;
		7939: rom = 27;
		7940: rom = 15;
		7941: rom = 25;
		7942: rom = 27;
		7943: rom = 27;
		7944: rom = 27;
		7945: rom = 27;
		7946: rom = 27;
		7947: rom = 27;
		7948: rom = 27;
		7949: rom = 27;
		7950: rom = 27;
		7951: rom = 27;
		7952: rom = 27;
		7953: rom = 27;
		7954: rom = 27;
		7955: rom = 27;
		7956: rom = 27;
		7957: rom = 27;
		7958: rom = 27;
		7959: rom = 27;
		7960: rom = 20;
		7961: rom = 12;
		7962: rom = 15;
		7963: rom = 11;
		7964: rom = 9;
		7965: rom = 17;
		7966: rom = 5;
		7967: rom = 17;
		7968: rom = 16;
		7969: rom = 15;
		7970: rom = 18;
		7971: rom = 18;
		7972: rom = 18;
		7973: rom = 18;
		7974: rom = 18;
		7975: rom = 11;
		7976: rom = 18;
		7977: rom = 13;
		7978: rom = 22;
		7979: rom = 27;
		7980: rom = 22;
		7981: rom = 17;
		7982: rom = 24;
		7983: rom = 25;
		7984: rom = 24;
		7985: rom = 12;
		7986: rom = 13;
		7987: rom = 20;
		7988: rom = 12;
		7989: rom = 14;
		7990: rom = 18;
		7991: rom = 18;
		7992: rom = 18;
		7993: rom = 18;
		7994: rom = 18;
		7995: rom = 18;
		7996: rom = 18;
		7997: rom = 18;
		7998: rom = 10;
		7999: rom = 18;
		8000: rom = 18;
		8001: rom = 18;
		8002: rom = 18;
		8003: rom = 18;
		8004: rom = 18;
		8005: rom = 17;
		8006: rom = 18;
		8007: rom = 24;
		8008: rom = 24;
		8009: rom = 24;
		8010: rom = 24;
		8011: rom = 24;
		8012: rom = 23;
		8013: rom = 12;
		8014: rom = 18;
		8015: rom = 20;
		8016: rom = 25;
		8017: rom = 23;
		8018: rom = 18;
		8019: rom = 18;
		8020: rom = 18;
		8021: rom = 18;
		8022: rom = 18;
		8023: rom = 18;
		8024: rom = 18;
		8025: rom = 18;
		8026: rom = 18;
		8027: rom = 18;
		8028: rom = 18;
		8029: rom = 18;
		8030: rom = 18;
		8031: rom = 18;
		8032: rom = 18;
		8033: rom = 18;
		8034: rom = 18;
		8035: rom = 18;
		8036: rom = 18;
		8037: rom = 18;
		8038: rom = 20;
		8039: rom = 25;
		8040: rom = 25;
		8041: rom = 25;
		8042: rom = 22;
		8043: rom = 15;
		8044: rom = 27;
		8045: rom = 27;
		8046: rom = 27;
		8047: rom = 27;
		8048: rom = 27;
		8049: rom = 27;
		8050: rom = 27;
		8051: rom = 27;
		8052: rom = 27;
		8053: rom = 27;
		8054: rom = 27;
		8055: rom = 27;
		8056: rom = 27;
		8057: rom = 27;
		8058: rom = 27;
		8064: rom = 27;
		8065: rom = 27;
		8066: rom = 27;
		8067: rom = 27;
		8068: rom = 27;
		8069: rom = 27;
		8070: rom = 27;
		8071: rom = 27;
		8072: rom = 27;
		8073: rom = 27;
		8074: rom = 27;
		8075: rom = 27;
		8076: rom = 27;
		8077: rom = 27;
		8078: rom = 27;
		8079: rom = 27;
		8080: rom = 27;
		8081: rom = 27;
		8082: rom = 27;
		8083: rom = 27;
		8084: rom = 27;
		8085: rom = 27;
		8086: rom = 27;
		8087: rom = 27;
		8088: rom = 27;
		8089: rom = 24;
		8090: rom = 22;
		8091: rom = 25;
		8092: rom = 15;
		8093: rom = 11;
		8094: rom = 12;
		8095: rom = 17;
		8096: rom = 18;
		8097: rom = 12;
		8098: rom = 18;
		8099: rom = 18;
		8100: rom = 18;
		8101: rom = 18;
		8102: rom = 18;
		8103: rom = 10;
		8104: rom = 13;
		8105: rom = 22;
		8106: rom = 27;
		8107: rom = 27;
		8108: rom = 21;
		8109: rom = 16;
		8110: rom = 18;
		8111: rom = 23;
		8112: rom = 25;
		8113: rom = 16;
		8114: rom = 15;
		8115: rom = 9;
		8116: rom = 9;
		8117: rom = 18;
		8118: rom = 14;
		8119: rom = 18;
		8120: rom = 18;
		8121: rom = 18;
		8122: rom = 18;
		8123: rom = 18;
		8124: rom = 18;
		8125: rom = 18;
		8126: rom = 16;
		8127: rom = 14;
		8128: rom = 18;
		8129: rom = 18;
		8130: rom = 18;
		8131: rom = 18;
		8132: rom = 18;
		8133: rom = 18;
		8134: rom = 21;
		8135: rom = 24;
		8136: rom = 24;
		8137: rom = 24;
		8138: rom = 24;
		8139: rom = 24;
		8140: rom = 19;
		8141: rom = 16;
		8142: rom = 18;
		8143: rom = 16;
		8144: rom = 15;
		8145: rom = 13;
		8146: rom = 16;
		8147: rom = 18;
		8148: rom = 18;
		8149: rom = 18;
		8150: rom = 18;
		8151: rom = 18;
		8152: rom = 18;
		8153: rom = 18;
		8154: rom = 18;
		8155: rom = 18;
		8156: rom = 18;
		8157: rom = 18;
		8158: rom = 18;
		8159: rom = 18;
		8160: rom = 18;
		8161: rom = 18;
		8162: rom = 18;
		8163: rom = 18;
		8164: rom = 18;
		8165: rom = 18;
		8166: rom = 21;
		8167: rom = 25;
		8168: rom = 24;
		8169: rom = 17;
		8170: rom = 18;
		8171: rom = 27;
		8172: rom = 27;
		8173: rom = 27;
		8174: rom = 27;
		8175: rom = 27;
		8176: rom = 27;
		8177: rom = 27;
		8178: rom = 27;
		8179: rom = 27;
		8180: rom = 27;
		8181: rom = 27;
		8182: rom = 27;
		8183: rom = 27;
		8184: rom = 27;
		8185: rom = 27;
		8186: rom = 27;
		8192: rom = 27;
		8193: rom = 27;
		8194: rom = 27;
		8195: rom = 27;
		8196: rom = 19;
		8197: rom = 19;
		8198: rom = 19;
		8199: rom = 19;
		8200: rom = 19;
		8201: rom = 19;
		8202: rom = 19;
		8203: rom = 19;
		8204: rom = 19;
		8205: rom = 19;
		8206: rom = 19;
		8207: rom = 22;
		8208: rom = 27;
		8209: rom = 27;
		8210: rom = 27;
		8211: rom = 27;
		8212: rom = 27;
		8213: rom = 27;
		8214: rom = 27;
		8215: rom = 27;
		8216: rom = 27;
		8217: rom = 27;
		8218: rom = 27;
		8219: rom = 27;
		8220: rom = 27;
		8221: rom = 27;
		8222: rom = 13;
		8223: rom = 16;
		8224: rom = 15;
		8225: rom = 12;
		8226: rom = 14;
		8227: rom = 15;
		8228: rom = 16;
		8229: rom = 15;
		8230: rom = 12;
		8231: rom = 16;
		8232: rom = 25;
		8233: rom = 27;
		8234: rom = 27;
		8235: rom = 27;
		8236: rom = 23;
		8237: rom = 15;
		8238: rom = 18;
		8239: rom = 18;
		8240: rom = 23;
		8241: rom = 16;
		8242: rom = 18;
		8243: rom = 18;
		8244: rom = 17;
		8245: rom = 7;
		8246: rom = 10;
		8247: rom = 17;
		8248: rom = 18;
		8249: rom = 18;
		8250: rom = 18;
		8251: rom = 18;
		8252: rom = 18;
		8253: rom = 18;
		8254: rom = 18;
		8255: rom = 10;
		8256: rom = 18;
		8257: rom = 18;
		8258: rom = 18;
		8259: rom = 18;
		8260: rom = 18;
		8261: rom = 18;
		8262: rom = 21;
		8263: rom = 24;
		8264: rom = 24;
		8265: rom = 24;
		8266: rom = 24;
		8267: rom = 24;
		8268: rom = 14;
		8269: rom = 16;
		8270: rom = 10;
		8271: rom = 13;
		8272: rom = 23;
		8273: rom = 24;
		8274: rom = 18;
		8275: rom = 18;
		8276: rom = 18;
		8277: rom = 18;
		8278: rom = 18;
		8279: rom = 18;
		8280: rom = 18;
		8281: rom = 18;
		8282: rom = 18;
		8283: rom = 18;
		8284: rom = 18;
		8285: rom = 18;
		8286: rom = 18;
		8287: rom = 18;
		8288: rom = 18;
		8289: rom = 18;
		8290: rom = 17;
		8291: rom = 13;
		8292: rom = 17;
		8293: rom = 18;
		8294: rom = 19;
		8295: rom = 16;
		8296: rom = 15;
		8297: rom = 24;
		8298: rom = 27;
		8299: rom = 27;
		8300: rom = 27;
		8301: rom = 27;
		8302: rom = 27;
		8303: rom = 27;
		8304: rom = 27;
		8305: rom = 27;
		8306: rom = 27;
		8307: rom = 27;
		8308: rom = 27;
		8309: rom = 27;
		8310: rom = 27;
		8311: rom = 27;
		8312: rom = 27;
		8313: rom = 27;
		8314: rom = 27;
		8320: rom = 27;
		8321: rom = 27;
		8322: rom = 27;
		8323: rom = 27;
		8324: rom = 0;
		8325: rom = 0;
		8326: rom = 0;
		8327: rom = 0;
		8328: rom = 0;
		8329: rom = 0;
		8330: rom = 0;
		8331: rom = 0;
		8332: rom = 0;
		8333: rom = 0;
		8334: rom = 0;
		8335: rom = 14;
		8336: rom = 27;
		8337: rom = 27;
		8338: rom = 27;
		8339: rom = 27;
		8340: rom = 27;
		8341: rom = 27;
		8342: rom = 27;
		8343: rom = 27;
		8344: rom = 27;
		8345: rom = 27;
		8346: rom = 27;
		8347: rom = 27;
		8348: rom = 27;
		8349: rom = 27;
		8350: rom = 23;
		8351: rom = 20;
		8352: rom = 20;
		8353: rom = 26;
		8354: rom = 27;
		8355: rom = 24;
		8356: rom = 23;
		8357: rom = 24;
		8358: rom = 26;
		8359: rom = 27;
		8360: rom = 27;
		8361: rom = 27;
		8362: rom = 27;
		8363: rom = 27;
		8364: rom = 25;
		8365: rom = 12;
		8366: rom = 18;
		8367: rom = 18;
		8368: rom = 18;
		8369: rom = 16;
		8370: rom = 17;
		8371: rom = 18;
		8372: rom = 18;
		8373: rom = 18;
		8374: rom = 18;
		8375: rom = 10;
		8376: rom = 17;
		8377: rom = 18;
		8378: rom = 18;
		8379: rom = 18;
		8380: rom = 18;
		8381: rom = 18;
		8382: rom = 18;
		8383: rom = 16;
		8384: rom = 12;
		8385: rom = 18;
		8386: rom = 18;
		8387: rom = 18;
		8388: rom = 18;
		8389: rom = 18;
		8390: rom = 18;
		8391: rom = 23;
		8392: rom = 24;
		8393: rom = 24;
		8394: rom = 24;
		8395: rom = 23;
		8396: rom = 5;
		8397: rom = 12;
		8398: rom = 18;
		8399: rom = 19;
		8400: rom = 25;
		8401: rom = 23;
		8402: rom = 18;
		8403: rom = 18;
		8404: rom = 18;
		8405: rom = 18;
		8406: rom = 18;
		8407: rom = 18;
		8408: rom = 18;
		8409: rom = 18;
		8410: rom = 18;
		8411: rom = 18;
		8412: rom = 18;
		8413: rom = 18;
		8414: rom = 18;
		8415: rom = 18;
		8416: rom = 18;
		8417: rom = 18;
		8418: rom = 18;
		8419: rom = 15;
		8420: rom = 9;
		8421: rom = 7;
		8422: rom = 19;
		8423: rom = 25;
		8424: rom = 27;
		8425: rom = 27;
		8426: rom = 27;
		8427: rom = 27;
		8428: rom = 27;
		8429: rom = 27;
		8430: rom = 27;
		8431: rom = 27;
		8432: rom = 27;
		8433: rom = 27;
		8434: rom = 27;
		8435: rom = 27;
		8436: rom = 27;
		8437: rom = 27;
		8438: rom = 27;
		8439: rom = 27;
		8440: rom = 27;
		8441: rom = 27;
		8442: rom = 27;
		8448: rom = 27;
		8449: rom = 27;
		8450: rom = 27;
		8451: rom = 27;
		8452: rom = 23;
		8453: rom = 23;
		8454: rom = 23;
		8455: rom = 23;
		8456: rom = 20;
		8457: rom = 0;
		8458: rom = 23;
		8459: rom = 23;
		8460: rom = 23;
		8461: rom = 23;
		8462: rom = 23;
		8463: rom = 24;
		8464: rom = 27;
		8465: rom = 27;
		8466: rom = 27;
		8467: rom = 27;
		8468: rom = 27;
		8469: rom = 27;
		8470: rom = 27;
		8471: rom = 27;
		8472: rom = 27;
		8473: rom = 27;
		8474: rom = 27;
		8475: rom = 27;
		8476: rom = 27;
		8477: rom = 27;
		8478: rom = 27;
		8479: rom = 27;
		8480: rom = 27;
		8481: rom = 27;
		8482: rom = 27;
		8483: rom = 27;
		8484: rom = 27;
		8485: rom = 27;
		8486: rom = 27;
		8487: rom = 27;
		8488: rom = 27;
		8489: rom = 27;
		8490: rom = 27;
		8491: rom = 27;
		8492: rom = 27;
		8493: rom = 14;
		8494: rom = 17;
		8495: rom = 18;
		8496: rom = 18;
		8497: rom = 14;
		8498: rom = 16;
		8499: rom = 18;
		8500: rom = 18;
		8501: rom = 18;
		8502: rom = 18;
		8503: rom = 18;
		8504: rom = 11;
		8505: rom = 11;
		8506: rom = 15;
		8507: rom = 17;
		8508: rom = 17;
		8509: rom = 17;
		8510: rom = 13;
		8511: rom = 9;
		8512: rom = 10;
		8513: rom = 17;
		8514: rom = 18;
		8515: rom = 18;
		8516: rom = 18;
		8517: rom = 18;
		8518: rom = 18;
		8519: rom = 20;
		8520: rom = 24;
		8521: rom = 24;
		8522: rom = 22;
		8523: rom = 12;
		8524: rom = 16;
		8525: rom = 18;
		8526: rom = 18;
		8527: rom = 22;
		8528: rom = 25;
		8529: rom = 21;
		8530: rom = 18;
		8531: rom = 18;
		8532: rom = 18;
		8533: rom = 18;
		8534: rom = 18;
		8535: rom = 18;
		8536: rom = 18;
		8537: rom = 18;
		8538: rom = 18;
		8539: rom = 18;
		8540: rom = 18;
		8541: rom = 18;
		8542: rom = 18;
		8543: rom = 18;
		8544: rom = 18;
		8545: rom = 18;
		8546: rom = 18;
		8547: rom = 18;
		8548: rom = 17;
		8549: rom = 14;
		8550: rom = 18;
		8551: rom = 27;
		8552: rom = 27;
		8553: rom = 27;
		8554: rom = 27;
		8555: rom = 27;
		8556: rom = 27;
		8557: rom = 27;
		8558: rom = 27;
		8559: rom = 27;
		8560: rom = 27;
		8561: rom = 27;
		8562: rom = 27;
		8563: rom = 27;
		8564: rom = 27;
		8565: rom = 27;
		8566: rom = 27;
		8567: rom = 27;
		8568: rom = 27;
		8569: rom = 27;
		8570: rom = 27;
		8576: rom = 27;
		8577: rom = 27;
		8578: rom = 27;
		8579: rom = 27;
		8580: rom = 27;
		8581: rom = 27;
		8582: rom = 27;
		8583: rom = 27;
		8584: rom = 24;
		8585: rom = 0;
		8586: rom = 27;
		8587: rom = 27;
		8588: rom = 27;
		8589: rom = 27;
		8590: rom = 27;
		8591: rom = 27;
		8592: rom = 27;
		8593: rom = 27;
		8594: rom = 27;
		8595: rom = 27;
		8596: rom = 27;
		8597: rom = 27;
		8598: rom = 27;
		8599: rom = 27;
		8600: rom = 27;
		8601: rom = 27;
		8602: rom = 27;
		8603: rom = 27;
		8604: rom = 27;
		8605: rom = 27;
		8606: rom = 27;
		8607: rom = 27;
		8608: rom = 27;
		8609: rom = 27;
		8610: rom = 27;
		8611: rom = 27;
		8612: rom = 27;
		8613: rom = 27;
		8614: rom = 27;
		8615: rom = 27;
		8616: rom = 27;
		8617: rom = 27;
		8618: rom = 27;
		8619: rom = 27;
		8620: rom = 27;
		8621: rom = 23;
		8622: rom = 12;
		8623: rom = 18;
		8624: rom = 18;
		8625: rom = 16;
		8626: rom = 13;
		8627: rom = 18;
		8628: rom = 18;
		8629: rom = 18;
		8630: rom = 18;
		8631: rom = 18;
		8632: rom = 18;
		8633: rom = 17;
		8634: rom = 14;
		8635: rom = 12;
		8636: rom = 12;
		8637: rom = 13;
		8638: rom = 15;
		8639: rom = 18;
		8640: rom = 18;
		8641: rom = 10;
		8642: rom = 18;
		8643: rom = 18;
		8644: rom = 18;
		8645: rom = 18;
		8646: rom = 18;
		8647: rom = 18;
		8648: rom = 23;
		8649: rom = 21;
		8650: rom = 11;
		8651: rom = 17;
		8652: rom = 18;
		8653: rom = 18;
		8654: rom = 20;
		8655: rom = 25;
		8656: rom = 24;
		8657: rom = 18;
		8658: rom = 18;
		8659: rom = 18;
		8660: rom = 18;
		8661: rom = 18;
		8662: rom = 18;
		8663: rom = 18;
		8664: rom = 18;
		8665: rom = 18;
		8666: rom = 18;
		8667: rom = 18;
		8668: rom = 18;
		8669: rom = 18;
		8670: rom = 18;
		8671: rom = 18;
		8672: rom = 18;
		8673: rom = 18;
		8674: rom = 18;
		8675: rom = 18;
		8676: rom = 18;
		8677: rom = 23;
		8678: rom = 21;
		8679: rom = 17;
		8680: rom = 27;
		8681: rom = 27;
		8682: rom = 27;
		8683: rom = 27;
		8684: rom = 27;
		8685: rom = 27;
		8686: rom = 27;
		8687: rom = 27;
		8688: rom = 27;
		8689: rom = 27;
		8690: rom = 27;
		8691: rom = 27;
		8692: rom = 27;
		8693: rom = 27;
		8694: rom = 27;
		8695: rom = 27;
		8696: rom = 27;
		8697: rom = 27;
		8698: rom = 27;
		8704: rom = 27;
		8705: rom = 27;
		8706: rom = 27;
		8707: rom = 27;
		8708: rom = 27;
		8709: rom = 27;
		8710: rom = 27;
		8711: rom = 27;
		8712: rom = 24;
		8713: rom = 0;
		8714: rom = 27;
		8715: rom = 27;
		8716: rom = 27;
		8717: rom = 27;
		8718: rom = 27;
		8719: rom = 27;
		8720: rom = 27;
		8721: rom = 27;
		8722: rom = 27;
		8723: rom = 27;
		8724: rom = 27;
		8725: rom = 27;
		8726: rom = 27;
		8727: rom = 27;
		8728: rom = 27;
		8729: rom = 27;
		8730: rom = 27;
		8731: rom = 27;
		8732: rom = 27;
		8733: rom = 27;
		8734: rom = 27;
		8735: rom = 27;
		8736: rom = 27;
		8737: rom = 27;
		8738: rom = 27;
		8739: rom = 27;
		8740: rom = 27;
		8741: rom = 27;
		8742: rom = 27;
		8743: rom = 27;
		8744: rom = 27;
		8745: rom = 27;
		8746: rom = 27;
		8747: rom = 27;
		8748: rom = 27;
		8749: rom = 27;
		8750: rom = 21;
		8751: rom = 11;
		8752: rom = 17;
		8753: rom = 18;
		8754: rom = 10;
		8755: rom = 18;
		8756: rom = 18;
		8757: rom = 18;
		8758: rom = 18;
		8759: rom = 18;
		8760: rom = 18;
		8761: rom = 18;
		8762: rom = 18;
		8763: rom = 18;
		8764: rom = 18;
		8765: rom = 18;
		8766: rom = 18;
		8767: rom = 15;
		8768: rom = 18;
		8769: rom = 15;
		8770: rom = 13;
		8771: rom = 18;
		8772: rom = 18;
		8773: rom = 18;
		8774: rom = 18;
		8775: rom = 18;
		8776: rom = 19;
		8777: rom = 11;
		8778: rom = 18;
		8779: rom = 18;
		8780: rom = 18;
		8781: rom = 19;
		8782: rom = 25;
		8783: rom = 25;
		8784: rom = 20;
		8785: rom = 18;
		8786: rom = 18;
		8787: rom = 18;
		8788: rom = 18;
		8789: rom = 18;
		8790: rom = 18;
		8791: rom = 18;
		8792: rom = 18;
		8793: rom = 18;
		8794: rom = 18;
		8795: rom = 18;
		8796: rom = 18;
		8797: rom = 18;
		8798: rom = 18;
		8799: rom = 18;
		8800: rom = 16;
		8801: rom = 17;
		8802: rom = 18;
		8803: rom = 18;
		8804: rom = 19;
		8805: rom = 25;
		8806: rom = 25;
		8807: rom = 20;
		8808: rom = 20;
		8809: rom = 27;
		8810: rom = 27;
		8811: rom = 27;
		8812: rom = 27;
		8813: rom = 27;
		8814: rom = 27;
		8815: rom = 27;
		8816: rom = 27;
		8817: rom = 27;
		8818: rom = 27;
		8819: rom = 27;
		8820: rom = 27;
		8821: rom = 27;
		8822: rom = 27;
		8823: rom = 27;
		8824: rom = 27;
		8825: rom = 27;
		8826: rom = 27;
		8832: rom = 27;
		8833: rom = 27;
		8834: rom = 27;
		8835: rom = 27;
		8836: rom = 27;
		8837: rom = 27;
		8838: rom = 27;
		8839: rom = 27;
		8840: rom = 24;
		8841: rom = 0;
		8842: rom = 27;
		8843: rom = 27;
		8844: rom = 27;
		8845: rom = 27;
		8846: rom = 27;
		8847: rom = 27;
		8848: rom = 27;
		8849: rom = 27;
		8850: rom = 27;
		8851: rom = 27;
		8852: rom = 27;
		8853: rom = 27;
		8854: rom = 27;
		8855: rom = 27;
		8856: rom = 27;
		8857: rom = 27;
		8858: rom = 27;
		8859: rom = 27;
		8860: rom = 27;
		8861: rom = 27;
		8862: rom = 27;
		8863: rom = 27;
		8864: rom = 27;
		8865: rom = 27;
		8866: rom = 27;
		8867: rom = 27;
		8868: rom = 27;
		8869: rom = 27;
		8870: rom = 27;
		8871: rom = 27;
		8872: rom = 27;
		8873: rom = 27;
		8874: rom = 27;
		8875: rom = 27;
		8876: rom = 27;
		8877: rom = 27;
		8878: rom = 27;
		8879: rom = 24;
		8880: rom = 14;
		8881: rom = 12;
		8882: rom = 9;
		8883: rom = 17;
		8884: rom = 18;
		8885: rom = 18;
		8886: rom = 18;
		8887: rom = 18;
		8888: rom = 18;
		8889: rom = 18;
		8890: rom = 18;
		8891: rom = 18;
		8892: rom = 18;
		8893: rom = 18;
		8894: rom = 18;
		8895: rom = 9;
		8896: rom = 11;
		8897: rom = 12;
		8898: rom = 10;
		8899: rom = 17;
		8900: rom = 18;
		8901: rom = 18;
		8902: rom = 18;
		8903: rom = 18;
		8904: rom = 10;
		8905: rom = 18;
		8906: rom = 18;
		8907: rom = 18;
		8908: rom = 19;
		8909: rom = 24;
		8910: rom = 25;
		8911: rom = 22;
		8912: rom = 18;
		8913: rom = 18;
		8914: rom = 18;
		8915: rom = 18;
		8916: rom = 18;
		8917: rom = 18;
		8918: rom = 18;
		8919: rom = 18;
		8920: rom = 18;
		8921: rom = 18;
		8922: rom = 18;
		8923: rom = 18;
		8924: rom = 18;
		8925: rom = 18;
		8926: rom = 18;
		8927: rom = 18;
		8928: rom = 14;
		8929: rom = 10;
		8930: rom = 10;
		8931: rom = 16;
		8932: rom = 21;
		8933: rom = 25;
		8934: rom = 25;
		8935: rom = 24;
		8936: rom = 14;
		8937: rom = 26;
		8938: rom = 27;
		8939: rom = 27;
		8940: rom = 27;
		8941: rom = 27;
		8942: rom = 27;
		8943: rom = 27;
		8944: rom = 27;
		8945: rom = 27;
		8946: rom = 27;
		8947: rom = 27;
		8948: rom = 27;
		8949: rom = 27;
		8950: rom = 27;
		8951: rom = 27;
		8952: rom = 27;
		8953: rom = 27;
		8954: rom = 27;
		8960: rom = 27;
		8961: rom = 27;
		8962: rom = 27;
		8963: rom = 27;
		8964: rom = 27;
		8965: rom = 27;
		8966: rom = 27;
		8967: rom = 27;
		8968: rom = 24;
		8969: rom = 0;
		8970: rom = 27;
		8971: rom = 27;
		8972: rom = 27;
		8973: rom = 27;
		8974: rom = 27;
		8975: rom = 27;
		8976: rom = 27;
		8977: rom = 27;
		8978: rom = 27;
		8979: rom = 27;
		8980: rom = 27;
		8981: rom = 27;
		8982: rom = 27;
		8983: rom = 27;
		8984: rom = 27;
		8985: rom = 27;
		8986: rom = 27;
		8987: rom = 27;
		8988: rom = 27;
		8989: rom = 27;
		8990: rom = 27;
		8991: rom = 27;
		8992: rom = 27;
		8993: rom = 27;
		8994: rom = 27;
		8995: rom = 27;
		8996: rom = 27;
		8997: rom = 27;
		8998: rom = 27;
		8999: rom = 27;
		9000: rom = 27;
		9001: rom = 27;
		9002: rom = 27;
		9003: rom = 27;
		9004: rom = 27;
		9005: rom = 27;
		9006: rom = 27;
		9007: rom = 27;
		9008: rom = 27;
		9009: rom = 25;
		9010: rom = 20;
		9011: rom = 12;
		9012: rom = 18;
		9013: rom = 18;
		9014: rom = 18;
		9015: rom = 18;
		9016: rom = 18;
		9017: rom = 18;
		9018: rom = 18;
		9019: rom = 18;
		9020: rom = 18;
		9021: rom = 18;
		9022: rom = 15;
		9023: rom = 14;
		9024: rom = 18;
		9025: rom = 16;
		9026: rom = 8;
		9027: rom = 7;
		9028: rom = 18;
		9029: rom = 18;
		9030: rom = 18;
		9031: rom = 10;
		9032: rom = 17;
		9033: rom = 18;
		9034: rom = 18;
		9035: rom = 20;
		9036: rom = 25;
		9037: rom = 25;
		9038: rom = 23;
		9039: rom = 18;
		9040: rom = 18;
		9041: rom = 18;
		9042: rom = 18;
		9043: rom = 18;
		9044: rom = 18;
		9045: rom = 18;
		9046: rom = 18;
		9047: rom = 18;
		9048: rom = 18;
		9049: rom = 18;
		9050: rom = 18;
		9051: rom = 18;
		9052: rom = 18;
		9053: rom = 18;
		9054: rom = 18;
		9055: rom = 18;
		9056: rom = 18;
		9057: rom = 18;
		9058: rom = 16;
		9059: rom = 10;
		9060: rom = 14;
		9061: rom = 15;
		9062: rom = 14;
		9063: rom = 17;
		9064: rom = 21;
		9065: rom = 26;
		9066: rom = 27;
		9067: rom = 27;
		9068: rom = 27;
		9069: rom = 27;
		9070: rom = 27;
		9071: rom = 27;
		9072: rom = 27;
		9073: rom = 27;
		9074: rom = 27;
		9075: rom = 27;
		9076: rom = 27;
		9077: rom = 27;
		9078: rom = 27;
		9079: rom = 27;
		9080: rom = 27;
		9081: rom = 27;
		9082: rom = 27;
		9088: rom = 27;
		9089: rom = 27;
		9090: rom = 27;
		9091: rom = 27;
		9092: rom = 27;
		9093: rom = 27;
		9094: rom = 27;
		9095: rom = 27;
		9096: rom = 24;
		9097: rom = 0;
		9098: rom = 27;
		9099: rom = 27;
		9100: rom = 27;
		9101: rom = 27;
		9102: rom = 27;
		9103: rom = 27;
		9104: rom = 27;
		9105: rom = 27;
		9106: rom = 27;
		9107: rom = 27;
		9108: rom = 27;
		9109: rom = 27;
		9110: rom = 27;
		9111: rom = 27;
		9112: rom = 27;
		9113: rom = 27;
		9114: rom = 27;
		9115: rom = 27;
		9116: rom = 27;
		9117: rom = 27;
		9118: rom = 27;
		9119: rom = 27;
		9120: rom = 27;
		9121: rom = 27;
		9122: rom = 27;
		9123: rom = 27;
		9124: rom = 27;
		9125: rom = 27;
		9126: rom = 27;
		9127: rom = 27;
		9128: rom = 27;
		9129: rom = 27;
		9130: rom = 27;
		9131: rom = 27;
		9132: rom = 27;
		9133: rom = 24;
		9134: rom = 21;
		9135: rom = 19;
		9136: rom = 17;
		9137: rom = 15;
		9138: rom = 13;
		9139: rom = 10;
		9140: rom = 14;
		9141: rom = 18;
		9142: rom = 18;
		9143: rom = 18;
		9144: rom = 18;
		9145: rom = 18;
		9146: rom = 18;
		9147: rom = 18;
		9148: rom = 18;
		9149: rom = 18;
		9150: rom = 9;
		9151: rom = 18;
		9152: rom = 18;
		9153: rom = 18;
		9154: rom = 18;
		9155: rom = 11;
		9156: rom = 11;
		9157: rom = 18;
		9158: rom = 14;
		9159: rom = 15;
		9160: rom = 18;
		9161: rom = 18;
		9162: rom = 20;
		9163: rom = 25;
		9164: rom = 25;
		9165: rom = 22;
		9166: rom = 18;
		9167: rom = 18;
		9168: rom = 18;
		9169: rom = 18;
		9170: rom = 18;
		9171: rom = 18;
		9172: rom = 18;
		9173: rom = 18;
		9174: rom = 18;
		9175: rom = 18;
		9176: rom = 18;
		9177: rom = 18;
		9178: rom = 18;
		9179: rom = 18;
		9180: rom = 18;
		9181: rom = 18;
		9182: rom = 18;
		9183: rom = 18;
		9184: rom = 18;
		9185: rom = 18;
		9186: rom = 18;
		9187: rom = 21;
		9188: rom = 17;
		9189: rom = 19;
		9190: rom = 27;
		9191: rom = 27;
		9192: rom = 27;
		9193: rom = 27;
		9194: rom = 27;
		9195: rom = 27;
		9196: rom = 27;
		9197: rom = 27;
		9198: rom = 27;
		9199: rom = 27;
		9200: rom = 27;
		9201: rom = 27;
		9202: rom = 27;
		9203: rom = 27;
		9204: rom = 27;
		9205: rom = 27;
		9206: rom = 27;
		9207: rom = 27;
		9208: rom = 27;
		9209: rom = 27;
		9210: rom = 27;
		9216: rom = 27;
		9217: rom = 27;
		9218: rom = 27;
		9219: rom = 27;
		9220: rom = 27;
		9221: rom = 27;
		9222: rom = 27;
		9223: rom = 27;
		9224: rom = 24;
		9225: rom = 0;
		9226: rom = 27;
		9227: rom = 27;
		9228: rom = 27;
		9229: rom = 27;
		9230: rom = 27;
		9231: rom = 27;
		9232: rom = 27;
		9233: rom = 27;
		9234: rom = 27;
		9235: rom = 27;
		9236: rom = 27;
		9237: rom = 27;
		9238: rom = 27;
		9239: rom = 27;
		9240: rom = 27;
		9241: rom = 27;
		9242: rom = 27;
		9243: rom = 27;
		9244: rom = 27;
		9245: rom = 27;
		9246: rom = 27;
		9247: rom = 27;
		9248: rom = 27;
		9249: rom = 27;
		9250: rom = 27;
		9251: rom = 27;
		9252: rom = 27;
		9253: rom = 27;
		9254: rom = 27;
		9255: rom = 27;
		9256: rom = 27;
		9257: rom = 27;
		9258: rom = 27;
		9259: rom = 27;
		9260: rom = 26;
		9261: rom = 9;
		9262: rom = 20;
		9263: rom = 21;
		9264: rom = 23;
		9265: rom = 23;
		9266: rom = 24;
		9267: rom = 24;
		9268: rom = 15;
		9269: rom = 15;
		9270: rom = 18;
		9271: rom = 18;
		9272: rom = 18;
		9273: rom = 18;
		9274: rom = 18;
		9275: rom = 18;
		9276: rom = 18;
		9277: rom = 12;
		9278: rom = 17;
		9279: rom = 18;
		9280: rom = 18;
		9281: rom = 18;
		9282: rom = 18;
		9283: rom = 18;
		9284: rom = 14;
		9285: rom = 13;
		9286: rom = 10;
		9287: rom = 18;
		9288: rom = 18;
		9289: rom = 19;
		9290: rom = 24;
		9291: rom = 25;
		9292: rom = 22;
		9293: rom = 18;
		9294: rom = 18;
		9295: rom = 18;
		9296: rom = 18;
		9297: rom = 18;
		9298: rom = 18;
		9299: rom = 18;
		9300: rom = 18;
		9301: rom = 18;
		9302: rom = 18;
		9303: rom = 18;
		9304: rom = 18;
		9305: rom = 18;
		9306: rom = 18;
		9307: rom = 18;
		9308: rom = 18;
		9309: rom = 18;
		9310: rom = 14;
		9311: rom = 17;
		9312: rom = 18;
		9313: rom = 18;
		9314: rom = 18;
		9315: rom = 25;
		9316: rom = 25;
		9317: rom = 13;
		9318: rom = 26;
		9319: rom = 27;
		9320: rom = 27;
		9321: rom = 27;
		9322: rom = 27;
		9323: rom = 27;
		9324: rom = 27;
		9325: rom = 27;
		9326: rom = 27;
		9327: rom = 27;
		9328: rom = 27;
		9329: rom = 27;
		9330: rom = 27;
		9331: rom = 27;
		9332: rom = 27;
		9333: rom = 27;
		9334: rom = 27;
		9335: rom = 27;
		9336: rom = 27;
		9337: rom = 27;
		9338: rom = 27;
		9344: rom = 27;
		9345: rom = 27;
		9346: rom = 27;
		9347: rom = 27;
		9348: rom = 1;
		9349: rom = 1;
		9350: rom = 1;
		9351: rom = 1;
		9352: rom = 1;
		9353: rom = 0;
		9354: rom = 1;
		9355: rom = 1;
		9356: rom = 1;
		9357: rom = 1;
		9358: rom = 1;
		9359: rom = 14;
		9360: rom = 27;
		9361: rom = 27;
		9362: rom = 27;
		9363: rom = 27;
		9364: rom = 27;
		9365: rom = 27;
		9366: rom = 27;
		9367: rom = 27;
		9368: rom = 27;
		9369: rom = 27;
		9370: rom = 27;
		9371: rom = 27;
		9372: rom = 27;
		9373: rom = 27;
		9374: rom = 27;
		9375: rom = 27;
		9376: rom = 27;
		9377: rom = 27;
		9378: rom = 27;
		9379: rom = 27;
		9380: rom = 27;
		9381: rom = 27;
		9382: rom = 27;
		9383: rom = 27;
		9384: rom = 27;
		9385: rom = 27;
		9386: rom = 27;
		9387: rom = 27;
		9388: rom = 27;
		9389: rom = 22;
		9390: rom = 13;
		9391: rom = 20;
		9392: rom = 23;
		9393: rom = 24;
		9394: rom = 24;
		9395: rom = 24;
		9396: rom = 23;
		9397: rom = 16;
		9398: rom = 12;
		9399: rom = 18;
		9400: rom = 18;
		9401: rom = 18;
		9402: rom = 18;
		9403: rom = 18;
		9404: rom = 13;
		9405: rom = 17;
		9406: rom = 25;
		9407: rom = 21;
		9408: rom = 18;
		9409: rom = 18;
		9410: rom = 18;
		9411: rom = 18;
		9412: rom = 18;
		9413: rom = 10;
		9414: rom = 16;
		9415: rom = 18;
		9416: rom = 18;
		9417: rom = 23;
		9418: rom = 25;
		9419: rom = 22;
		9420: rom = 18;
		9421: rom = 18;
		9422: rom = 18;
		9423: rom = 18;
		9424: rom = 18;
		9425: rom = 18;
		9426: rom = 18;
		9427: rom = 18;
		9428: rom = 18;
		9429: rom = 18;
		9430: rom = 18;
		9431: rom = 18;
		9432: rom = 18;
		9433: rom = 18;
		9434: rom = 18;
		9435: rom = 18;
		9436: rom = 18;
		9437: rom = 18;
		9438: rom = 16;
		9439: rom = 10;
		9440: rom = 12;
		9441: rom = 17;
		9442: rom = 22;
		9443: rom = 25;
		9444: rom = 25;
		9445: rom = 20;
		9446: rom = 16;
		9447: rom = 27;
		9448: rom = 27;
		9449: rom = 27;
		9450: rom = 27;
		9451: rom = 27;
		9452: rom = 27;
		9453: rom = 27;
		9454: rom = 27;
		9455: rom = 27;
		9456: rom = 27;
		9457: rom = 27;
		9458: rom = 27;
		9459: rom = 27;
		9460: rom = 27;
		9461: rom = 27;
		9462: rom = 27;
		9463: rom = 27;
		9464: rom = 27;
		9465: rom = 27;
		9466: rom = 27;
		9472: rom = 27;
		9473: rom = 27;
		9474: rom = 27;
		9475: rom = 27;
		9476: rom = 13;
		9477: rom = 13;
		9478: rom = 13;
		9479: rom = 13;
		9480: rom = 13;
		9481: rom = 13;
		9482: rom = 13;
		9483: rom = 13;
		9484: rom = 13;
		9485: rom = 13;
		9486: rom = 13;
		9487: rom = 18;
		9488: rom = 27;
		9489: rom = 27;
		9490: rom = 27;
		9491: rom = 27;
		9492: rom = 27;
		9493: rom = 27;
		9494: rom = 27;
		9495: rom = 27;
		9496: rom = 27;
		9497: rom = 27;
		9498: rom = 27;
		9499: rom = 27;
		9500: rom = 27;
		9501: rom = 27;
		9502: rom = 27;
		9503: rom = 27;
		9504: rom = 27;
		9505: rom = 27;
		9506: rom = 27;
		9507: rom = 27;
		9508: rom = 27;
		9509: rom = 27;
		9510: rom = 27;
		9511: rom = 27;
		9512: rom = 27;
		9513: rom = 27;
		9514: rom = 27;
		9515: rom = 27;
		9516: rom = 27;
		9517: rom = 27;
		9518: rom = 26;
		9519: rom = 21;
		9520: rom = 14;
		9521: rom = 15;
		9522: rom = 19;
		9523: rom = 22;
		9524: rom = 24;
		9525: rom = 24;
		9526: rom = 20;
		9527: rom = 7;
		9528: rom = 11;
		9529: rom = 13;
		9530: rom = 13;
		9531: rom = 9;
		9532: rom = 8;
		9533: rom = 20;
		9534: rom = 25;
		9535: rom = 25;
		9536: rom = 19;
		9537: rom = 18;
		9538: rom = 18;
		9539: rom = 18;
		9540: rom = 18;
		9541: rom = 11;
		9542: rom = 18;
		9543: rom = 18;
		9544: rom = 20;
		9545: rom = 25;
		9546: rom = 24;
		9547: rom = 18;
		9548: rom = 18;
		9549: rom = 18;
		9550: rom = 18;
		9551: rom = 18;
		9552: rom = 18;
		9553: rom = 18;
		9554: rom = 18;
		9555: rom = 18;
		9556: rom = 18;
		9557: rom = 18;
		9558: rom = 18;
		9559: rom = 18;
		9560: rom = 18;
		9561: rom = 18;
		9562: rom = 18;
		9563: rom = 18;
		9564: rom = 18;
		9565: rom = 18;
		9566: rom = 18;
		9567: rom = 18;
		9568: rom = 14;
		9569: rom = 9;
		9570: rom = 19;
		9571: rom = 20;
		9572: rom = 21;
		9573: rom = 17;
		9574: rom = 6;
		9575: rom = 25;
		9576: rom = 27;
		9577: rom = 27;
		9578: rom = 27;
		9579: rom = 27;
		9580: rom = 27;
		9581: rom = 27;
		9582: rom = 27;
		9583: rom = 27;
		9584: rom = 27;
		9585: rom = 27;
		9586: rom = 27;
		9587: rom = 27;
		9588: rom = 27;
		9589: rom = 27;
		9590: rom = 27;
		9591: rom = 27;
		9592: rom = 27;
		9593: rom = 27;
		9594: rom = 27;
		9600: rom = 27;
		9601: rom = 27;
		9602: rom = 27;
		9603: rom = 27;
		9604: rom = 27;
		9605: rom = 27;
		9606: rom = 27;
		9607: rom = 27;
		9608: rom = 27;
		9609: rom = 27;
		9610: rom = 27;
		9611: rom = 27;
		9612: rom = 27;
		9613: rom = 27;
		9614: rom = 27;
		9615: rom = 27;
		9616: rom = 27;
		9617: rom = 27;
		9618: rom = 27;
		9619: rom = 27;
		9620: rom = 27;
		9621: rom = 27;
		9622: rom = 27;
		9623: rom = 27;
		9624: rom = 27;
		9625: rom = 27;
		9626: rom = 27;
		9627: rom = 27;
		9628: rom = 27;
		9629: rom = 27;
		9630: rom = 27;
		9631: rom = 27;
		9632: rom = 27;
		9633: rom = 27;
		9634: rom = 27;
		9635: rom = 27;
		9636: rom = 27;
		9637: rom = 27;
		9638: rom = 27;
		9639: rom = 27;
		9640: rom = 27;
		9641: rom = 27;
		9642: rom = 27;
		9643: rom = 27;
		9644: rom = 27;
		9645: rom = 27;
		9646: rom = 27;
		9647: rom = 27;
		9648: rom = 27;
		9649: rom = 26;
		9650: rom = 21;
		9651: rom = 16;
		9652: rom = 10;
		9653: rom = 12;
		9654: rom = 13;
		9655: rom = 17;
		9656: rom = 21;
		9657: rom = 21;
		9658: rom = 21;
		9659: rom = 23;
		9660: rom = 19;
		9661: rom = 11;
		9662: rom = 16;
		9663: rom = 22;
		9664: rom = 23;
		9665: rom = 18;
		9666: rom = 18;
		9667: rom = 18;
		9668: rom = 14;
		9669: rom = 16;
		9670: rom = 18;
		9671: rom = 18;
		9672: rom = 23;
		9673: rom = 25;
		9674: rom = 20;
		9675: rom = 18;
		9676: rom = 18;
		9677: rom = 18;
		9678: rom = 18;
		9679: rom = 18;
		9680: rom = 18;
		9681: rom = 18;
		9682: rom = 18;
		9683: rom = 18;
		9684: rom = 18;
		9685: rom = 18;
		9686: rom = 18;
		9687: rom = 18;
		9688: rom = 18;
		9689: rom = 18;
		9690: rom = 18;
		9691: rom = 18;
		9692: rom = 18;
		9693: rom = 18;
		9694: rom = 18;
		9695: rom = 18;
		9696: rom = 18;
		9697: rom = 21;
		9698: rom = 11;
		9699: rom = 11;
		9700: rom = 13;
		9701: rom = 14;
		9702: rom = 16;
		9703: rom = 16;
		9704: rom = 27;
		9705: rom = 27;
		9706: rom = 27;
		9707: rom = 27;
		9708: rom = 27;
		9709: rom = 27;
		9710: rom = 27;
		9711: rom = 27;
		9712: rom = 27;
		9713: rom = 27;
		9714: rom = 27;
		9715: rom = 27;
		9716: rom = 27;
		9717: rom = 27;
		9718: rom = 27;
		9719: rom = 27;
		9720: rom = 27;
		9721: rom = 27;
		9722: rom = 27;
		9728: rom = 27;
		9729: rom = 27;
		9730: rom = 27;
		9731: rom = 27;
		9732: rom = 27;
		9733: rom = 27;
		9734: rom = 27;
		9735: rom = 27;
		9736: rom = 27;
		9737: rom = 27;
		9738: rom = 27;
		9739: rom = 27;
		9740: rom = 27;
		9741: rom = 27;
		9742: rom = 27;
		9743: rom = 27;
		9744: rom = 27;
		9745: rom = 27;
		9746: rom = 27;
		9747: rom = 27;
		9748: rom = 27;
		9749: rom = 27;
		9750: rom = 27;
		9751: rom = 27;
		9752: rom = 27;
		9753: rom = 27;
		9754: rom = 27;
		9755: rom = 27;
		9756: rom = 27;
		9757: rom = 27;
		9758: rom = 27;
		9759: rom = 27;
		9760: rom = 27;
		9761: rom = 27;
		9762: rom = 27;
		9763: rom = 27;
		9764: rom = 27;
		9765: rom = 27;
		9766: rom = 27;
		9767: rom = 27;
		9768: rom = 27;
		9769: rom = 27;
		9770: rom = 27;
		9771: rom = 27;
		9772: rom = 27;
		9773: rom = 27;
		9774: rom = 27;
		9775: rom = 27;
		9776: rom = 27;
		9777: rom = 27;
		9778: rom = 21;
		9779: rom = 13;
		9780: rom = 19;
		9781: rom = 23;
		9782: rom = 24;
		9783: rom = 24;
		9784: rom = 24;
		9785: rom = 24;
		9786: rom = 24;
		9787: rom = 24;
		9788: rom = 24;
		9789: rom = 24;
		9790: rom = 21;
		9791: rom = 13;
		9792: rom = 7;
		9793: rom = 10;
		9794: rom = 14;
		9795: rom = 14;
		9796: rom = 10;
		9797: rom = 18;
		9798: rom = 18;
		9799: rom = 19;
		9800: rom = 25;
		9801: rom = 24;
		9802: rom = 18;
		9803: rom = 18;
		9804: rom = 18;
		9805: rom = 18;
		9806: rom = 18;
		9807: rom = 18;
		9808: rom = 18;
		9809: rom = 18;
		9810: rom = 18;
		9811: rom = 18;
		9812: rom = 18;
		9813: rom = 18;
		9814: rom = 18;
		9815: rom = 18;
		9816: rom = 18;
		9817: rom = 18;
		9818: rom = 18;
		9819: rom = 18;
		9820: rom = 18;
		9821: rom = 18;
		9822: rom = 18;
		9823: rom = 18;
		9824: rom = 18;
		9825: rom = 25;
		9826: rom = 24;
		9827: rom = 13;
		9828: rom = 16;
		9829: rom = 18;
		9830: rom = 18;
		9831: rom = 12;
		9832: rom = 24;
		9833: rom = 27;
		9834: rom = 27;
		9835: rom = 27;
		9836: rom = 27;
		9837: rom = 27;
		9838: rom = 27;
		9839: rom = 27;
		9840: rom = 27;
		9841: rom = 27;
		9842: rom = 27;
		9843: rom = 27;
		9844: rom = 27;
		9845: rom = 27;
		9846: rom = 27;
		9847: rom = 27;
		9848: rom = 27;
		9849: rom = 27;
		9850: rom = 27;
		9856: rom = 27;
		9857: rom = 27;
		9858: rom = 27;
		9859: rom = 27;
		9860: rom = 27;
		9861: rom = 27;
		9862: rom = 27;
		9863: rom = 27;
		9864: rom = 24;
		9865: rom = 22;
		9866: rom = 23;
		9867: rom = 25;
		9868: rom = 27;
		9869: rom = 27;
		9870: rom = 27;
		9871: rom = 27;
		9872: rom = 27;
		9873: rom = 27;
		9874: rom = 27;
		9875: rom = 27;
		9876: rom = 27;
		9877: rom = 27;
		9878: rom = 27;
		9879: rom = 27;
		9880: rom = 27;
		9881: rom = 27;
		9882: rom = 27;
		9883: rom = 27;
		9884: rom = 27;
		9885: rom = 27;
		9886: rom = 27;
		9887: rom = 27;
		9888: rom = 27;
		9889: rom = 27;
		9890: rom = 27;
		9891: rom = 27;
		9892: rom = 27;
		9893: rom = 27;
		9894: rom = 27;
		9895: rom = 27;
		9896: rom = 27;
		9897: rom = 27;
		9898: rom = 27;
		9899: rom = 27;
		9900: rom = 27;
		9901: rom = 27;
		9902: rom = 27;
		9903: rom = 27;
		9904: rom = 27;
		9905: rom = 24;
		9906: rom = 12;
		9907: rom = 23;
		9908: rom = 24;
		9909: rom = 24;
		9910: rom = 24;
		9911: rom = 24;
		9912: rom = 24;
		9913: rom = 24;
		9914: rom = 24;
		9915: rom = 24;
		9916: rom = 23;
		9917: rom = 20;
		9918: rom = 13;
		9919: rom = 15;
		9920: rom = 21;
		9921: rom = 23;
		9922: rom = 21;
		9923: rom = 18;
		9924: rom = 12;
		9925: rom = 18;
		9926: rom = 18;
		9927: rom = 21;
		9928: rom = 25;
		9929: rom = 22;
		9930: rom = 18;
		9931: rom = 18;
		9932: rom = 18;
		9933: rom = 18;
		9934: rom = 18;
		9935: rom = 18;
		9936: rom = 18;
		9937: rom = 18;
		9938: rom = 18;
		9939: rom = 18;
		9940: rom = 18;
		9941: rom = 18;
		9942: rom = 18;
		9943: rom = 18;
		9944: rom = 18;
		9945: rom = 18;
		9946: rom = 18;
		9947: rom = 18;
		9948: rom = 18;
		9949: rom = 18;
		9950: rom = 18;
		9951: rom = 18;
		9952: rom = 20;
		9953: rom = 25;
		9954: rom = 25;
		9955: rom = 24;
		9956: rom = 10;
		9957: rom = 18;
		9958: rom = 18;
		9959: rom = 17;
		9960: rom = 16;
		9961: rom = 27;
		9962: rom = 27;
		9963: rom = 27;
		9964: rom = 27;
		9965: rom = 27;
		9966: rom = 27;
		9967: rom = 27;
		9968: rom = 27;
		9969: rom = 27;
		9970: rom = 27;
		9971: rom = 27;
		9972: rom = 27;
		9973: rom = 27;
		9974: rom = 27;
		9975: rom = 27;
		9976: rom = 27;
		9977: rom = 27;
		9978: rom = 27;
		9984: rom = 27;
		9985: rom = 27;
		9986: rom = 27;
		9987: rom = 27;
		9988: rom = 27;
		9989: rom = 27;
		9990: rom = 19;
		9991: rom = 0;
		9992: rom = 0;
		9993: rom = 0;
		9994: rom = 0;
		9995: rom = 0;
		9996: rom = 11;
		9997: rom = 23;
		9998: rom = 27;
		9999: rom = 27;
		10000: rom = 27;
		10001: rom = 27;
		10002: rom = 27;
		10003: rom = 27;
		10004: rom = 27;
		10005: rom = 27;
		10006: rom = 27;
		10007: rom = 27;
		10008: rom = 27;
		10009: rom = 27;
		10010: rom = 27;
		10011: rom = 27;
		10012: rom = 27;
		10013: rom = 27;
		10014: rom = 27;
		10015: rom = 27;
		10016: rom = 27;
		10017: rom = 27;
		10018: rom = 27;
		10019: rom = 27;
		10020: rom = 27;
		10021: rom = 27;
		10022: rom = 27;
		10023: rom = 27;
		10024: rom = 27;
		10025: rom = 27;
		10026: rom = 27;
		10027: rom = 27;
		10028: rom = 27;
		10029: rom = 27;
		10030: rom = 27;
		10031: rom = 27;
		10032: rom = 27;
		10033: rom = 27;
		10034: rom = 22;
		10035: rom = 15;
		10036: rom = 14;
		10037: rom = 17;
		10038: rom = 19;
		10039: rom = 21;
		10040: rom = 22;
		10041: rom = 23;
		10042: rom = 23;
		10043: rom = 19;
		10044: rom = 12;
		10045: rom = 17;
		10046: rom = 23;
		10047: rom = 24;
		10048: rom = 24;
		10049: rom = 24;
		10050: rom = 24;
		10051: rom = 19;
		10052: rom = 16;
		10053: rom = 18;
		10054: rom = 18;
		10055: rom = 22;
		10056: rom = 25;
		10057: rom = 20;
		10058: rom = 18;
		10059: rom = 18;
		10060: rom = 18;
		10061: rom = 18;
		10062: rom = 18;
		10063: rom = 18;
		10064: rom = 18;
		10065: rom = 18;
		10066: rom = 18;
		10067: rom = 18;
		10068: rom = 18;
		10069: rom = 18;
		10070: rom = 18;
		10071: rom = 18;
		10072: rom = 18;
		10073: rom = 18;
		10074: rom = 18;
		10075: rom = 18;
		10076: rom = 18;
		10077: rom = 18;
		10078: rom = 18;
		10079: rom = 18;
		10080: rom = 22;
		10081: rom = 25;
		10082: rom = 25;
		10083: rom = 17;
		10084: rom = 14;
		10085: rom = 18;
		10086: rom = 18;
		10087: rom = 18;
		10088: rom = 12;
		10089: rom = 25;
		10090: rom = 27;
		10091: rom = 27;
		10092: rom = 27;
		10093: rom = 27;
		10094: rom = 27;
		10095: rom = 27;
		10096: rom = 27;
		10097: rom = 27;
		10098: rom = 27;
		10099: rom = 27;
		10100: rom = 27;
		10101: rom = 27;
		10102: rom = 27;
		10103: rom = 27;
		10104: rom = 27;
		10105: rom = 27;
		10106: rom = 27;
		10112: rom = 27;
		10113: rom = 27;
		10114: rom = 27;
		10115: rom = 27;
		10116: rom = 27;
		10117: rom = 14;
		10118: rom = 0;
		10119: rom = 0;
		10120: rom = 16;
		10121: rom = 18;
		10122: rom = 18;
		10123: rom = 14;
		10124: rom = 0;
		10125: rom = 0;
		10126: rom = 22;
		10127: rom = 27;
		10128: rom = 27;
		10129: rom = 27;
		10130: rom = 27;
		10131: rom = 27;
		10132: rom = 27;
		10133: rom = 27;
		10134: rom = 27;
		10135: rom = 27;
		10136: rom = 27;
		10137: rom = 27;
		10138: rom = 27;
		10139: rom = 27;
		10140: rom = 27;
		10141: rom = 27;
		10142: rom = 27;
		10143: rom = 27;
		10144: rom = 27;
		10145: rom = 27;
		10146: rom = 27;
		10147: rom = 27;
		10148: rom = 27;
		10149: rom = 27;
		10150: rom = 27;
		10151: rom = 27;
		10152: rom = 27;
		10153: rom = 27;
		10154: rom = 27;
		10155: rom = 27;
		10156: rom = 27;
		10157: rom = 27;
		10158: rom = 27;
		10159: rom = 27;
		10160: rom = 27;
		10161: rom = 27;
		10162: rom = 27;
		10163: rom = 27;
		10164: rom = 27;
		10165: rom = 24;
		10166: rom = 22;
		10167: rom = 20;
		10168: rom = 18;
		10169: rom = 10;
		10170: rom = 7;
		10171: rom = 18;
		10172: rom = 23;
		10173: rom = 24;
		10174: rom = 24;
		10175: rom = 24;
		10176: rom = 24;
		10177: rom = 24;
		10178: rom = 24;
		10179: rom = 14;
		10180: rom = 18;
		10181: rom = 18;
		10182: rom = 18;
		10183: rom = 22;
		10184: rom = 25;
		10185: rom = 20;
		10186: rom = 18;
		10187: rom = 18;
		10188: rom = 18;
		10189: rom = 18;
		10190: rom = 18;
		10191: rom = 18;
		10192: rom = 18;
		10193: rom = 18;
		10194: rom = 18;
		10195: rom = 18;
		10196: rom = 18;
		10197: rom = 18;
		10198: rom = 18;
		10199: rom = 18;
		10200: rom = 18;
		10201: rom = 18;
		10202: rom = 18;
		10203: rom = 18;
		10204: rom = 18;
		10205: rom = 18;
		10206: rom = 18;
		10207: rom = 18;
		10208: rom = 23;
		10209: rom = 24;
		10210: rom = 15;
		10211: rom = 14;
		10212: rom = 18;
		10213: rom = 18;
		10214: rom = 18;
		10215: rom = 18;
		10216: rom = 17;
		10217: rom = 18;
		10218: rom = 27;
		10219: rom = 27;
		10220: rom = 27;
		10221: rom = 27;
		10222: rom = 27;
		10223: rom = 27;
		10224: rom = 27;
		10225: rom = 27;
		10226: rom = 27;
		10227: rom = 27;
		10228: rom = 27;
		10229: rom = 27;
		10230: rom = 27;
		10231: rom = 27;
		10232: rom = 27;
		10233: rom = 27;
		10234: rom = 27;
		10240: rom = 27;
		10241: rom = 27;
		10242: rom = 27;
		10243: rom = 27;
		10244: rom = 20;
		10245: rom = 0;
		10246: rom = 19;
		10247: rom = 27;
		10248: rom = 27;
		10249: rom = 27;
		10250: rom = 27;
		10251: rom = 27;
		10252: rom = 25;
		10253: rom = 12;
		10254: rom = 0;
		10255: rom = 25;
		10256: rom = 27;
		10257: rom = 27;
		10258: rom = 27;
		10259: rom = 27;
		10260: rom = 27;
		10261: rom = 27;
		10262: rom = 27;
		10263: rom = 27;
		10264: rom = 27;
		10265: rom = 27;
		10266: rom = 27;
		10267: rom = 27;
		10268: rom = 27;
		10269: rom = 27;
		10270: rom = 27;
		10271: rom = 27;
		10272: rom = 27;
		10273: rom = 27;
		10274: rom = 27;
		10275: rom = 27;
		10276: rom = 27;
		10277: rom = 27;
		10278: rom = 27;
		10279: rom = 27;
		10280: rom = 27;
		10281: rom = 27;
		10282: rom = 27;
		10283: rom = 27;
		10284: rom = 27;
		10285: rom = 27;
		10286: rom = 27;
		10287: rom = 27;
		10288: rom = 27;
		10289: rom = 27;
		10290: rom = 27;
		10291: rom = 27;
		10292: rom = 27;
		10293: rom = 27;
		10294: rom = 27;
		10295: rom = 26;
		10296: rom = 16;
		10297: rom = 16;
		10298: rom = 23;
		10299: rom = 24;
		10300: rom = 24;
		10301: rom = 24;
		10302: rom = 24;
		10303: rom = 24;
		10304: rom = 24;
		10305: rom = 24;
		10306: rom = 24;
		10307: rom = 11;
		10308: rom = 18;
		10309: rom = 18;
		10310: rom = 18;
		10311: rom = 21;
		10312: rom = 25;
		10313: rom = 21;
		10314: rom = 18;
		10315: rom = 18;
		10316: rom = 18;
		10317: rom = 18;
		10318: rom = 18;
		10319: rom = 18;
		10320: rom = 18;
		10321: rom = 18;
		10322: rom = 18;
		10323: rom = 18;
		10324: rom = 18;
		10325: rom = 18;
		10326: rom = 18;
		10327: rom = 18;
		10328: rom = 18;
		10329: rom = 18;
		10330: rom = 18;
		10331: rom = 18;
		10332: rom = 17;
		10333: rom = 18;
		10334: rom = 18;
		10335: rom = 17;
		10336: rom = 17;
		10337: rom = 10;
		10338: rom = 16;
		10339: rom = 18;
		10340: rom = 18;
		10341: rom = 18;
		10342: rom = 18;
		10343: rom = 18;
		10344: rom = 18;
		10345: rom = 11;
		10346: rom = 26;
		10347: rom = 27;
		10348: rom = 27;
		10349: rom = 27;
		10350: rom = 27;
		10351: rom = 27;
		10352: rom = 27;
		10353: rom = 27;
		10354: rom = 27;
		10355: rom = 27;
		10356: rom = 27;
		10357: rom = 27;
		10358: rom = 27;
		10359: rom = 27;
		10360: rom = 27;
		10361: rom = 27;
		10362: rom = 27;
		10368: rom = 27;
		10369: rom = 27;
		10370: rom = 27;
		10371: rom = 27;
		10372: rom = 0;
		10373: rom = 18;
		10374: rom = 27;
		10375: rom = 27;
		10376: rom = 27;
		10377: rom = 27;
		10378: rom = 27;
		10379: rom = 27;
		10380: rom = 27;
		10381: rom = 26;
		10382: rom = 0;
		10383: rom = 18;
		10384: rom = 27;
		10385: rom = 27;
		10386: rom = 27;
		10387: rom = 27;
		10388: rom = 27;
		10389: rom = 27;
		10390: rom = 27;
		10391: rom = 27;
		10392: rom = 27;
		10393: rom = 27;
		10394: rom = 27;
		10395: rom = 27;
		10396: rom = 27;
		10397: rom = 27;
		10398: rom = 27;
		10399: rom = 27;
		10400: rom = 27;
		10401: rom = 27;
		10402: rom = 27;
		10403: rom = 27;
		10404: rom = 27;
		10405: rom = 27;
		10406: rom = 27;
		10407: rom = 27;
		10408: rom = 27;
		10409: rom = 27;
		10410: rom = 27;
		10411: rom = 27;
		10412: rom = 27;
		10413: rom = 27;
		10414: rom = 27;
		10415: rom = 27;
		10416: rom = 27;
		10417: rom = 27;
		10418: rom = 27;
		10419: rom = 27;
		10420: rom = 27;
		10421: rom = 27;
		10422: rom = 22;
		10423: rom = 14;
		10424: rom = 22;
		10425: rom = 24;
		10426: rom = 24;
		10427: rom = 24;
		10428: rom = 24;
		10429: rom = 24;
		10430: rom = 24;
		10431: rom = 24;
		10432: rom = 24;
		10433: rom = 24;
		10434: rom = 21;
		10435: rom = 13;
		10436: rom = 18;
		10437: rom = 18;
		10438: rom = 18;
		10439: rom = 19;
		10440: rom = 25;
		10441: rom = 24;
		10442: rom = 18;
		10443: rom = 18;
		10444: rom = 18;
		10445: rom = 18;
		10446: rom = 18;
		10447: rom = 18;
		10448: rom = 18;
		10449: rom = 18;
		10450: rom = 18;
		10451: rom = 18;
		10452: rom = 18;
		10453: rom = 18;
		10454: rom = 18;
		10455: rom = 18;
		10456: rom = 18;
		10457: rom = 18;
		10458: rom = 18;
		10459: rom = 14;
		10460: rom = 15;
		10461: rom = 16;
		10462: rom = 12;
		10463: rom = 9;
		10464: rom = 15;
		10465: rom = 17;
		10466: rom = 18;
		10467: rom = 18;
		10468: rom = 18;
		10469: rom = 18;
		10470: rom = 18;
		10471: rom = 18;
		10472: rom = 18;
		10473: rom = 15;
		10474: rom = 21;
		10475: rom = 27;
		10476: rom = 27;
		10477: rom = 27;
		10478: rom = 27;
		10479: rom = 27;
		10480: rom = 27;
		10481: rom = 27;
		10482: rom = 27;
		10483: rom = 27;
		10484: rom = 27;
		10485: rom = 27;
		10486: rom = 27;
		10487: rom = 27;
		10488: rom = 27;
		10489: rom = 27;
		10490: rom = 27;
		10496: rom = 27;
		10497: rom = 27;
		10498: rom = 27;
		10499: rom = 24;
		10500: rom = 0;
		10501: rom = 26;
		10502: rom = 27;
		10503: rom = 27;
		10504: rom = 27;
		10505: rom = 27;
		10506: rom = 27;
		10507: rom = 27;
		10508: rom = 27;
		10509: rom = 27;
		10510: rom = 19;
		10511: rom = 0;
		10512: rom = 27;
		10513: rom = 27;
		10514: rom = 27;
		10515: rom = 27;
		10516: rom = 27;
		10517: rom = 27;
		10518: rom = 27;
		10519: rom = 27;
		10520: rom = 27;
		10521: rom = 27;
		10522: rom = 27;
		10523: rom = 27;
		10524: rom = 27;
		10525: rom = 27;
		10526: rom = 27;
		10527: rom = 27;
		10528: rom = 27;
		10529: rom = 27;
		10530: rom = 27;
		10531: rom = 27;
		10532: rom = 27;
		10533: rom = 27;
		10534: rom = 27;
		10535: rom = 27;
		10536: rom = 27;
		10537: rom = 27;
		10538: rom = 27;
		10539: rom = 27;
		10540: rom = 27;
		10541: rom = 27;
		10542: rom = 27;
		10543: rom = 27;
		10544: rom = 27;
		10545: rom = 27;
		10546: rom = 27;
		10547: rom = 27;
		10548: rom = 27;
		10549: rom = 25;
		10550: rom = 14;
		10551: rom = 23;
		10552: rom = 24;
		10553: rom = 24;
		10554: rom = 24;
		10555: rom = 24;
		10556: rom = 24;
		10557: rom = 24;
		10558: rom = 24;
		10559: rom = 22;
		10560: rom = 18;
		10561: rom = 13;
		10562: rom = 12;
		10563: rom = 16;
		10564: rom = 18;
		10565: rom = 18;
		10566: rom = 18;
		10567: rom = 18;
		10568: rom = 23;
		10569: rom = 25;
		10570: rom = 24;
		10571: rom = 19;
		10572: rom = 18;
		10573: rom = 18;
		10574: rom = 18;
		10575: rom = 18;
		10576: rom = 18;
		10577: rom = 18;
		10578: rom = 18;
		10579: rom = 18;
		10580: rom = 18;
		10581: rom = 18;
		10582: rom = 18;
		10583: rom = 18;
		10584: rom = 18;
		10585: rom = 18;
		10586: rom = 17;
		10587: rom = 5;
		10588: rom = 9;
		10589: rom = 11;
		10590: rom = 16;
		10591: rom = 18;
		10592: rom = 18;
		10593: rom = 18;
		10594: rom = 18;
		10595: rom = 18;
		10596: rom = 18;
		10597: rom = 18;
		10598: rom = 18;
		10599: rom = 18;
		10600: rom = 18;
		10601: rom = 18;
		10602: rom = 13;
		10603: rom = 27;
		10604: rom = 27;
		10605: rom = 27;
		10606: rom = 27;
		10607: rom = 27;
		10608: rom = 27;
		10609: rom = 27;
		10610: rom = 27;
		10611: rom = 27;
		10612: rom = 27;
		10613: rom = 27;
		10614: rom = 27;
		10615: rom = 27;
		10616: rom = 27;
		10617: rom = 27;
		10618: rom = 27;
		10624: rom = 27;
		10625: rom = 27;
		10626: rom = 27;
		10627: rom = 0;
		10628: rom = 1;
		10629: rom = 27;
		10630: rom = 27;
		10631: rom = 27;
		10632: rom = 27;
		10633: rom = 27;
		10634: rom = 27;
		10635: rom = 27;
		10636: rom = 27;
		10637: rom = 27;
		10638: rom = 23;
		10639: rom = 5;
		10640: rom = 0;
		10641: rom = 27;
		10642: rom = 27;
		10643: rom = 27;
		10644: rom = 27;
		10645: rom = 27;
		10646: rom = 27;
		10647: rom = 27;
		10648: rom = 27;
		10649: rom = 27;
		10650: rom = 27;
		10651: rom = 27;
		10652: rom = 27;
		10653: rom = 27;
		10654: rom = 27;
		10655: rom = 27;
		10656: rom = 27;
		10657: rom = 27;
		10658: rom = 27;
		10659: rom = 27;
		10660: rom = 27;
		10661: rom = 27;
		10662: rom = 27;
		10663: rom = 27;
		10664: rom = 27;
		10665: rom = 27;
		10666: rom = 27;
		10667: rom = 27;
		10668: rom = 27;
		10669: rom = 27;
		10670: rom = 27;
		10671: rom = 27;
		10672: rom = 27;
		10673: rom = 27;
		10674: rom = 27;
		10675: rom = 27;
		10676: rom = 27;
		10677: rom = 27;
		10678: rom = 16;
		10679: rom = 15;
		10680: rom = 19;
		10681: rom = 21;
		10682: rom = 21;
		10683: rom = 20;
		10684: rom = 17;
		10685: rom = 15;
		10686: rom = 13;
		10687: rom = 18;
		10688: rom = 23;
		10689: rom = 27;
		10690: rom = 20;
		10691: rom = 17;
		10692: rom = 18;
		10693: rom = 18;
		10694: rom = 18;
		10695: rom = 18;
		10696: rom = 19;
		10697: rom = 24;
		10698: rom = 25;
		10699: rom = 25;
		10700: rom = 23;
		10701: rom = 20;
		10702: rom = 18;
		10703: rom = 18;
		10704: rom = 18;
		10705: rom = 18;
		10706: rom = 18;
		10707: rom = 18;
		10708: rom = 18;
		10709: rom = 18;
		10710: rom = 19;
		10711: rom = 21;
		10712: rom = 23;
		10713: rom = 24;
		10714: rom = 13;
		10715: rom = 16;
		10716: rom = 18;
		10717: rom = 18;
		10718: rom = 18;
		10719: rom = 18;
		10720: rom = 18;
		10721: rom = 18;
		10722: rom = 18;
		10723: rom = 18;
		10724: rom = 18;
		10725: rom = 18;
		10726: rom = 18;
		10727: rom = 18;
		10728: rom = 18;
		10729: rom = 18;
		10730: rom = 13;
		10731: rom = 24;
		10732: rom = 27;
		10733: rom = 27;
		10734: rom = 27;
		10735: rom = 27;
		10736: rom = 27;
		10737: rom = 27;
		10738: rom = 27;
		10739: rom = 27;
		10740: rom = 27;
		10741: rom = 27;
		10742: rom = 27;
		10743: rom = 27;
		10744: rom = 27;
		10745: rom = 27;
		10746: rom = 27;
		10752: rom = 27;
		10753: rom = 27;
		10754: rom = 27;
		10755: rom = 0;
		10756: rom = 1;
		10757: rom = 27;
		10758: rom = 27;
		10759: rom = 27;
		10760: rom = 27;
		10761: rom = 27;
		10762: rom = 27;
		10763: rom = 27;
		10764: rom = 27;
		10765: rom = 27;
		10766: rom = 23;
		10767: rom = 6;
		10768: rom = 0;
		10769: rom = 27;
		10770: rom = 27;
		10771: rom = 27;
		10772: rom = 27;
		10773: rom = 27;
		10774: rom = 27;
		10775: rom = 27;
		10776: rom = 27;
		10777: rom = 27;
		10778: rom = 27;
		10779: rom = 27;
		10780: rom = 27;
		10781: rom = 27;
		10782: rom = 27;
		10783: rom = 27;
		10784: rom = 27;
		10785: rom = 27;
		10786: rom = 27;
		10787: rom = 27;
		10788: rom = 27;
		10789: rom = 27;
		10790: rom = 27;
		10791: rom = 27;
		10792: rom = 27;
		10793: rom = 27;
		10794: rom = 27;
		10795: rom = 27;
		10796: rom = 27;
		10797: rom = 27;
		10798: rom = 27;
		10799: rom = 27;
		10800: rom = 27;
		10801: rom = 27;
		10802: rom = 27;
		10803: rom = 27;
		10804: rom = 27;
		10805: rom = 27;
		10806: rom = 27;
		10807: rom = 26;
		10808: rom = 22;
		10809: rom = 20;
		10810: rom = 20;
		10811: rom = 21;
		10812: rom = 24;
		10813: rom = 26;
		10814: rom = 27;
		10815: rom = 27;
		10816: rom = 27;
		10817: rom = 27;
		10818: rom = 19;
		10819: rom = 18;
		10820: rom = 18;
		10821: rom = 18;
		10822: rom = 18;
		10823: rom = 18;
		10824: rom = 18;
		10825: rom = 18;
		10826: rom = 22;
		10827: rom = 25;
		10828: rom = 25;
		10829: rom = 25;
		10830: rom = 25;
		10831: rom = 24;
		10832: rom = 23;
		10833: rom = 23;
		10834: rom = 23;
		10835: rom = 23;
		10836: rom = 24;
		10837: rom = 25;
		10838: rom = 25;
		10839: rom = 25;
		10840: rom = 24;
		10841: rom = 13;
		10842: rom = 16;
		10843: rom = 18;
		10844: rom = 18;
		10845: rom = 18;
		10846: rom = 18;
		10847: rom = 18;
		10848: rom = 18;
		10849: rom = 18;
		10850: rom = 18;
		10851: rom = 18;
		10852: rom = 18;
		10853: rom = 18;
		10854: rom = 18;
		10855: rom = 18;
		10856: rom = 18;
		10857: rom = 18;
		10858: rom = 17;
		10859: rom = 18;
		10860: rom = 27;
		10861: rom = 27;
		10862: rom = 27;
		10863: rom = 27;
		10864: rom = 27;
		10865: rom = 27;
		10866: rom = 27;
		10867: rom = 27;
		10868: rom = 27;
		10869: rom = 27;
		10870: rom = 27;
		10871: rom = 27;
		10872: rom = 27;
		10873: rom = 27;
		10874: rom = 27;
		10880: rom = 27;
		10881: rom = 27;
		10882: rom = 27;
		10883: rom = 25;
		10884: rom = 0;
		10885: rom = 25;
		10886: rom = 27;
		10887: rom = 27;
		10888: rom = 27;
		10889: rom = 27;
		10890: rom = 27;
		10891: rom = 27;
		10892: rom = 27;
		10893: rom = 27;
		10894: rom = 18;
		10895: rom = 0;
		10896: rom = 27;
		10897: rom = 27;
		10898: rom = 27;
		10899: rom = 27;
		10900: rom = 27;
		10901: rom = 27;
		10902: rom = 27;
		10903: rom = 27;
		10904: rom = 27;
		10905: rom = 27;
		10906: rom = 27;
		10907: rom = 27;
		10908: rom = 27;
		10909: rom = 27;
		10910: rom = 27;
		10911: rom = 27;
		10912: rom = 27;
		10913: rom = 27;
		10914: rom = 27;
		10915: rom = 27;
		10916: rom = 27;
		10917: rom = 27;
		10918: rom = 27;
		10919: rom = 27;
		10920: rom = 27;
		10921: rom = 27;
		10922: rom = 27;
		10923: rom = 27;
		10924: rom = 27;
		10925: rom = 27;
		10926: rom = 27;
		10927: rom = 27;
		10928: rom = 27;
		10929: rom = 27;
		10930: rom = 27;
		10931: rom = 27;
		10932: rom = 27;
		10933: rom = 27;
		10934: rom = 27;
		10935: rom = 27;
		10936: rom = 27;
		10937: rom = 27;
		10938: rom = 27;
		10939: rom = 27;
		10940: rom = 27;
		10941: rom = 27;
		10942: rom = 27;
		10943: rom = 27;
		10944: rom = 27;
		10945: rom = 27;
		10946: rom = 15;
		10947: rom = 18;
		10948: rom = 18;
		10949: rom = 18;
		10950: rom = 18;
		10951: rom = 18;
		10952: rom = 18;
		10953: rom = 18;
		10954: rom = 18;
		10955: rom = 19;
		10956: rom = 22;
		10957: rom = 24;
		10958: rom = 25;
		10959: rom = 25;
		10960: rom = 25;
		10961: rom = 25;
		10962: rom = 25;
		10963: rom = 25;
		10964: rom = 25;
		10965: rom = 25;
		10966: rom = 24;
		10967: rom = 21;
		10968: rom = 11;
		10969: rom = 16;
		10970: rom = 18;
		10971: rom = 18;
		10972: rom = 18;
		10973: rom = 18;
		10974: rom = 18;
		10975: rom = 18;
		10976: rom = 18;
		10977: rom = 18;
		10978: rom = 18;
		10979: rom = 18;
		10980: rom = 18;
		10981: rom = 18;
		10982: rom = 18;
		10983: rom = 18;
		10984: rom = 18;
		10985: rom = 18;
		10986: rom = 18;
		10987: rom = 12;
		10988: rom = 27;
		10989: rom = 27;
		10990: rom = 27;
		10991: rom = 27;
		10992: rom = 27;
		10993: rom = 27;
		10994: rom = 27;
		10995: rom = 27;
		10996: rom = 27;
		10997: rom = 27;
		10998: rom = 27;
		10999: rom = 27;
		11000: rom = 27;
		11001: rom = 27;
		11002: rom = 27;
		11008: rom = 27;
		11009: rom = 27;
		11010: rom = 27;
		11011: rom = 27;
		11012: rom = 0;
		11013: rom = 15;
		11014: rom = 27;
		11015: rom = 27;
		11016: rom = 27;
		11017: rom = 27;
		11018: rom = 27;
		11019: rom = 27;
		11020: rom = 27;
		11021: rom = 25;
		11022: rom = 0;
		11023: rom = 20;
		11024: rom = 27;
		11025: rom = 27;
		11026: rom = 27;
		11027: rom = 27;
		11028: rom = 27;
		11029: rom = 27;
		11030: rom = 27;
		11031: rom = 27;
		11032: rom = 27;
		11033: rom = 27;
		11034: rom = 27;
		11035: rom = 27;
		11036: rom = 27;
		11037: rom = 27;
		11038: rom = 27;
		11039: rom = 27;
		11040: rom = 27;
		11041: rom = 27;
		11042: rom = 27;
		11043: rom = 27;
		11044: rom = 27;
		11045: rom = 27;
		11046: rom = 27;
		11047: rom = 27;
		11048: rom = 27;
		11049: rom = 27;
		11050: rom = 27;
		11051: rom = 27;
		11052: rom = 27;
		11053: rom = 27;
		11054: rom = 27;
		11055: rom = 27;
		11056: rom = 27;
		11057: rom = 27;
		11058: rom = 27;
		11059: rom = 27;
		11060: rom = 27;
		11061: rom = 27;
		11062: rom = 27;
		11063: rom = 27;
		11064: rom = 27;
		11065: rom = 27;
		11066: rom = 27;
		11067: rom = 27;
		11068: rom = 27;
		11069: rom = 27;
		11070: rom = 27;
		11071: rom = 27;
		11072: rom = 27;
		11073: rom = 27;
		11074: rom = 15;
		11075: rom = 18;
		11076: rom = 18;
		11077: rom = 18;
		11078: rom = 18;
		11079: rom = 18;
		11080: rom = 18;
		11081: rom = 18;
		11082: rom = 18;
		11083: rom = 18;
		11084: rom = 18;
		11085: rom = 18;
		11086: rom = 18;
		11087: rom = 20;
		11088: rom = 20;
		11089: rom = 20;
		11090: rom = 20;
		11091: rom = 20;
		11092: rom = 20;
		11093: rom = 18;
		11094: rom = 12;
		11095: rom = 12;
		11096: rom = 10;
		11097: rom = 16;
		11098: rom = 18;
		11099: rom = 18;
		11100: rom = 18;
		11101: rom = 18;
		11102: rom = 18;
		11103: rom = 18;
		11104: rom = 18;
		11105: rom = 18;
		11106: rom = 18;
		11107: rom = 18;
		11108: rom = 18;
		11109: rom = 18;
		11110: rom = 18;
		11111: rom = 18;
		11112: rom = 18;
		11113: rom = 18;
		11114: rom = 18;
		11115: rom = 14;
		11116: rom = 23;
		11117: rom = 27;
		11118: rom = 27;
		11119: rom = 27;
		11120: rom = 27;
		11121: rom = 27;
		11122: rom = 27;
		11123: rom = 27;
		11124: rom = 27;
		11125: rom = 27;
		11126: rom = 27;
		11127: rom = 27;
		11128: rom = 27;
		11129: rom = 27;
		11130: rom = 27;
		11136: rom = 27;
		11137: rom = 27;
		11138: rom = 27;
		11139: rom = 27;
		11140: rom = 22;
		11141: rom = 0;
		11142: rom = 15;
		11143: rom = 25;
		11144: rom = 27;
		11145: rom = 27;
		11146: rom = 27;
		11147: rom = 27;
		11148: rom = 22;
		11149: rom = 0;
		11150: rom = 0;
		11151: rom = 26;
		11152: rom = 27;
		11153: rom = 27;
		11154: rom = 27;
		11155: rom = 27;
		11156: rom = 27;
		11157: rom = 27;
		11158: rom = 27;
		11159: rom = 27;
		11160: rom = 27;
		11161: rom = 27;
		11162: rom = 27;
		11163: rom = 27;
		11164: rom = 27;
		11165: rom = 27;
		11166: rom = 27;
		11167: rom = 27;
		11168: rom = 27;
		11169: rom = 27;
		11170: rom = 27;
		11171: rom = 27;
		11172: rom = 27;
		11173: rom = 27;
		11174: rom = 27;
		11175: rom = 27;
		11176: rom = 27;
		11177: rom = 27;
		11178: rom = 27;
		11179: rom = 27;
		11180: rom = 27;
		11181: rom = 27;
		11182: rom = 27;
		11183: rom = 27;
		11184: rom = 27;
		11185: rom = 27;
		11186: rom = 27;
		11187: rom = 27;
		11188: rom = 27;
		11189: rom = 27;
		11190: rom = 27;
		11191: rom = 27;
		11192: rom = 27;
		11193: rom = 27;
		11194: rom = 27;
		11195: rom = 27;
		11196: rom = 27;
		11197: rom = 27;
		11198: rom = 27;
		11199: rom = 27;
		11200: rom = 27;
		11201: rom = 27;
		11202: rom = 15;
		11203: rom = 18;
		11204: rom = 18;
		11205: rom = 18;
		11206: rom = 18;
		11207: rom = 18;
		11208: rom = 18;
		11209: rom = 18;
		11210: rom = 18;
		11211: rom = 18;
		11212: rom = 18;
		11213: rom = 18;
		11214: rom = 18;
		11215: rom = 18;
		11216: rom = 18;
		11217: rom = 18;
		11218: rom = 18;
		11219: rom = 17;
		11220: rom = 12;
		11221: rom = 10;
		11222: rom = 16;
		11223: rom = 18;
		11224: rom = 17;
		11225: rom = 10;
		11226: rom = 17;
		11227: rom = 18;
		11228: rom = 18;
		11229: rom = 18;
		11230: rom = 18;
		11231: rom = 18;
		11232: rom = 18;
		11233: rom = 18;
		11234: rom = 18;
		11235: rom = 18;
		11236: rom = 18;
		11237: rom = 18;
		11238: rom = 18;
		11239: rom = 18;
		11240: rom = 18;
		11241: rom = 18;
		11242: rom = 18;
		11243: rom = 17;
		11244: rom = 18;
		11245: rom = 27;
		11246: rom = 27;
		11247: rom = 27;
		11248: rom = 27;
		11249: rom = 27;
		11250: rom = 27;
		11251: rom = 27;
		11252: rom = 27;
		11253: rom = 27;
		11254: rom = 27;
		11255: rom = 27;
		11256: rom = 27;
		11257: rom = 27;
		11258: rom = 27;
		11264: rom = 27;
		11265: rom = 27;
		11266: rom = 27;
		11267: rom = 27;
		11268: rom = 27;
		11269: rom = 18;
		11270: rom = 0;
		11271: rom = 0;
		11272: rom = 9;
		11273: rom = 15;
		11274: rom = 14;
		11275: rom = 0;
		11276: rom = 0;
		11277: rom = 0;
		11278: rom = 24;
		11279: rom = 27;
		11280: rom = 27;
		11281: rom = 27;
		11282: rom = 27;
		11283: rom = 27;
		11284: rom = 27;
		11285: rom = 27;
		11286: rom = 27;
		11287: rom = 27;
		11288: rom = 27;
		11289: rom = 27;
		11290: rom = 27;
		11291: rom = 27;
		11292: rom = 27;
		11293: rom = 27;
		11294: rom = 27;
		11295: rom = 27;
		11296: rom = 27;
		11297: rom = 27;
		11298: rom = 27;
		11299: rom = 27;
		11300: rom = 27;
		11301: rom = 27;
		11302: rom = 27;
		11303: rom = 27;
		11304: rom = 27;
		11305: rom = 27;
		11306: rom = 27;
		11307: rom = 27;
		11308: rom = 27;
		11309: rom = 27;
		11310: rom = 27;
		11311: rom = 27;
		11312: rom = 27;
		11313: rom = 27;
		11314: rom = 27;
		11315: rom = 27;
		11316: rom = 27;
		11317: rom = 27;
		11318: rom = 27;
		11319: rom = 27;
		11320: rom = 27;
		11321: rom = 27;
		11322: rom = 27;
		11323: rom = 27;
		11324: rom = 27;
		11325: rom = 27;
		11326: rom = 27;
		11327: rom = 27;
		11328: rom = 27;
		11329: rom = 27;
		11330: rom = 18;
		11331: rom = 18;
		11332: rom = 18;
		11333: rom = 18;
		11334: rom = 18;
		11335: rom = 18;
		11336: rom = 18;
		11337: rom = 18;
		11338: rom = 18;
		11339: rom = 18;
		11340: rom = 18;
		11341: rom = 18;
		11342: rom = 18;
		11343: rom = 18;
		11344: rom = 17;
		11345: rom = 14;
		11346: rom = 10;
		11347: rom = 12;
		11348: rom = 16;
		11349: rom = 18;
		11350: rom = 18;
		11351: rom = 18;
		11352: rom = 18;
		11353: rom = 16;
		11354: rom = 11;
		11355: rom = 18;
		11356: rom = 18;
		11357: rom = 18;
		11358: rom = 18;
		11359: rom = 18;
		11360: rom = 18;
		11361: rom = 18;
		11362: rom = 18;
		11363: rom = 18;
		11364: rom = 18;
		11365: rom = 18;
		11366: rom = 18;
		11367: rom = 18;
		11368: rom = 18;
		11369: rom = 18;
		11370: rom = 18;
		11371: rom = 18;
		11372: rom = 12;
		11373: rom = 27;
		11374: rom = 27;
		11375: rom = 27;
		11376: rom = 27;
		11377: rom = 27;
		11378: rom = 27;
		11379: rom = 27;
		11380: rom = 27;
		11381: rom = 27;
		11382: rom = 27;
		11383: rom = 27;
		11384: rom = 27;
		11385: rom = 27;
		11386: rom = 27;
		11392: rom = 27;
		11393: rom = 27;
		11394: rom = 27;
		11395: rom = 27;
		11396: rom = 27;
		11397: rom = 27;
		11398: rom = 23;
		11399: rom = 13;
		11400: rom = 1;
		11401: rom = 0;
		11402: rom = 0;
		11403: rom = 0;
		11404: rom = 17;
		11405: rom = 25;
		11406: rom = 27;
		11407: rom = 27;
		11408: rom = 27;
		11409: rom = 27;
		11410: rom = 27;
		11411: rom = 27;
		11412: rom = 27;
		11413: rom = 27;
		11414: rom = 27;
		11415: rom = 27;
		11416: rom = 27;
		11417: rom = 27;
		11418: rom = 27;
		11419: rom = 27;
		11420: rom = 27;
		11421: rom = 27;
		11422: rom = 27;
		11423: rom = 27;
		11424: rom = 27;
		11425: rom = 27;
		11426: rom = 27;
		11427: rom = 27;
		11428: rom = 27;
		11429: rom = 27;
		11430: rom = 27;
		11431: rom = 27;
		11432: rom = 27;
		11433: rom = 27;
		11434: rom = 27;
		11435: rom = 27;
		11436: rom = 27;
		11437: rom = 27;
		11438: rom = 27;
		11439: rom = 27;
		11440: rom = 27;
		11441: rom = 27;
		11442: rom = 27;
		11443: rom = 27;
		11444: rom = 27;
		11445: rom = 27;
		11446: rom = 27;
		11447: rom = 27;
		11448: rom = 27;
		11449: rom = 27;
		11450: rom = 27;
		11451: rom = 27;
		11452: rom = 27;
		11453: rom = 27;
		11454: rom = 27;
		11455: rom = 27;
		11456: rom = 27;
		11457: rom = 27;
		11458: rom = 20;
		11459: rom = 16;
		11460: rom = 18;
		11461: rom = 18;
		11462: rom = 18;
		11463: rom = 18;
		11464: rom = 18;
		11465: rom = 18;
		11466: rom = 18;
		11467: rom = 17;
		11468: rom = 15;
		11469: rom = 13;
		11470: rom = 10;
		11471: rom = 10;
		11472: rom = 12;
		11473: rom = 8;
		11474: rom = 17;
		11475: rom = 18;
		11476: rom = 18;
		11477: rom = 18;
		11478: rom = 18;
		11479: rom = 18;
		11480: rom = 18;
		11481: rom = 18;
		11482: rom = 14;
		11483: rom = 14;
		11484: rom = 18;
		11485: rom = 18;
		11486: rom = 18;
		11487: rom = 18;
		11488: rom = 18;
		11489: rom = 18;
		11490: rom = 18;
		11491: rom = 18;
		11492: rom = 18;
		11493: rom = 18;
		11494: rom = 18;
		11495: rom = 18;
		11496: rom = 18;
		11497: rom = 18;
		11498: rom = 18;
		11499: rom = 18;
		11500: rom = 13;
		11501: rom = 25;
		11502: rom = 27;
		11503: rom = 27;
		11504: rom = 27;
		11505: rom = 27;
		11506: rom = 27;
		11507: rom = 27;
		11508: rom = 27;
		11509: rom = 27;
		11510: rom = 27;
		11511: rom = 27;
		11512: rom = 27;
		11513: rom = 27;
		11514: rom = 27;
		11520: rom = 27;
		11521: rom = 27;
		11522: rom = 27;
		11523: rom = 27;
		11524: rom = 27;
		11525: rom = 27;
		11526: rom = 27;
		11527: rom = 27;
		11528: rom = 27;
		11529: rom = 25;
		11530: rom = 26;
		11531: rom = 27;
		11532: rom = 27;
		11533: rom = 27;
		11534: rom = 27;
		11535: rom = 27;
		11536: rom = 27;
		11537: rom = 27;
		11538: rom = 27;
		11539: rom = 27;
		11540: rom = 27;
		11541: rom = 27;
		11542: rom = 27;
		11543: rom = 27;
		11544: rom = 27;
		11545: rom = 27;
		11546: rom = 27;
		11547: rom = 27;
		11548: rom = 27;
		11549: rom = 27;
		11550: rom = 27;
		11551: rom = 27;
		11552: rom = 27;
		11553: rom = 27;
		11554: rom = 27;
		11555: rom = 27;
		11556: rom = 27;
		11557: rom = 27;
		11558: rom = 27;
		11559: rom = 27;
		11560: rom = 27;
		11561: rom = 27;
		11562: rom = 27;
		11563: rom = 27;
		11564: rom = 27;
		11565: rom = 27;
		11566: rom = 27;
		11567: rom = 27;
		11568: rom = 27;
		11569: rom = 27;
		11570: rom = 27;
		11571: rom = 27;
		11572: rom = 27;
		11573: rom = 27;
		11574: rom = 27;
		11575: rom = 27;
		11576: rom = 27;
		11577: rom = 27;
		11578: rom = 27;
		11579: rom = 27;
		11580: rom = 27;
		11581: rom = 27;
		11582: rom = 27;
		11583: rom = 27;
		11584: rom = 27;
		11585: rom = 27;
		11586: rom = 24;
		11587: rom = 14;
		11588: rom = 18;
		11589: rom = 18;
		11590: rom = 18;
		11591: rom = 18;
		11592: rom = 18;
		11593: rom = 18;
		11594: rom = 18;
		11595: rom = 18;
		11596: rom = 18;
		11597: rom = 18;
		11598: rom = 18;
		11599: rom = 18;
		11600: rom = 18;
		11601: rom = 17;
		11602: rom = 10;
		11603: rom = 18;
		11604: rom = 18;
		11605: rom = 18;
		11606: rom = 18;
		11607: rom = 18;
		11608: rom = 18;
		11609: rom = 18;
		11610: rom = 18;
		11611: rom = 10;
		11612: rom = 17;
		11613: rom = 18;
		11614: rom = 18;
		11615: rom = 18;
		11616: rom = 18;
		11617: rom = 18;
		11618: rom = 18;
		11619: rom = 18;
		11620: rom = 18;
		11621: rom = 18;
		11622: rom = 18;
		11623: rom = 18;
		11624: rom = 18;
		11625: rom = 18;
		11626: rom = 18;
		11627: rom = 18;
		11628: rom = 16;
		11629: rom = 20;
		11630: rom = 27;
		11631: rom = 27;
		11632: rom = 27;
		11633: rom = 27;
		11634: rom = 27;
		11635: rom = 27;
		11636: rom = 27;
		11637: rom = 27;
		11638: rom = 27;
		11639: rom = 27;
		11640: rom = 27;
		11641: rom = 27;
		11642: rom = 27;
		11648: rom = 27;
		11649: rom = 27;
		11650: rom = 27;
		11651: rom = 27;
		11652: rom = 27;
		11653: rom = 27;
		11654: rom = 27;
		11655: rom = 27;
		11656: rom = 27;
		11657: rom = 27;
		11658: rom = 27;
		11659: rom = 27;
		11660: rom = 27;
		11661: rom = 27;
		11662: rom = 27;
		11663: rom = 27;
		11664: rom = 27;
		11665: rom = 27;
		11666: rom = 27;
		11667: rom = 27;
		11668: rom = 27;
		11669: rom = 27;
		11670: rom = 27;
		11671: rom = 27;
		11672: rom = 27;
		11673: rom = 27;
		11674: rom = 27;
		11675: rom = 27;
		11676: rom = 27;
		11677: rom = 27;
		11678: rom = 27;
		11679: rom = 27;
		11680: rom = 27;
		11681: rom = 27;
		11682: rom = 27;
		11683: rom = 27;
		11684: rom = 27;
		11685: rom = 27;
		11686: rom = 27;
		11687: rom = 27;
		11688: rom = 27;
		11689: rom = 27;
		11690: rom = 27;
		11691: rom = 27;
		11692: rom = 27;
		11693: rom = 27;
		11694: rom = 27;
		11695: rom = 27;
		11696: rom = 27;
		11697: rom = 27;
		11698: rom = 27;
		11699: rom = 27;
		11700: rom = 27;
		11701: rom = 27;
		11702: rom = 27;
		11703: rom = 27;
		11704: rom = 27;
		11705: rom = 27;
		11706: rom = 27;
		11707: rom = 27;
		11708: rom = 27;
		11709: rom = 27;
		11710: rom = 27;
		11711: rom = 27;
		11712: rom = 27;
		11713: rom = 27;
		11714: rom = 27;
		11715: rom = 12;
		11716: rom = 18;
		11717: rom = 18;
		11718: rom = 18;
		11719: rom = 18;
		11720: rom = 18;
		11721: rom = 18;
		11722: rom = 18;
		11723: rom = 18;
		11724: rom = 18;
		11725: rom = 18;
		11726: rom = 18;
		11727: rom = 18;
		11728: rom = 18;
		11729: rom = 18;
		11730: rom = 16;
		11731: rom = 13;
		11732: rom = 18;
		11733: rom = 18;
		11734: rom = 18;
		11735: rom = 18;
		11736: rom = 18;
		11737: rom = 18;
		11738: rom = 18;
		11739: rom = 17;
		11740: rom = 11;
		11741: rom = 18;
		11742: rom = 18;
		11743: rom = 18;
		11744: rom = 18;
		11745: rom = 18;
		11746: rom = 18;
		11747: rom = 18;
		11748: rom = 18;
		11749: rom = 18;
		11750: rom = 18;
		11751: rom = 18;
		11752: rom = 18;
		11753: rom = 18;
		11754: rom = 18;
		11755: rom = 18;
		11756: rom = 18;
		11757: rom = 15;
		11758: rom = 27;
		11759: rom = 27;
		11760: rom = 27;
		11761: rom = 27;
		11762: rom = 27;
		11763: rom = 27;
		11764: rom = 27;
		11765: rom = 27;
		11766: rom = 27;
		11767: rom = 27;
		11768: rom = 27;
		11769: rom = 27;
		11770: rom = 27;
		11776: rom = 27;
		11777: rom = 27;
		11778: rom = 27;
		11779: rom = 27;
		11780: rom = 27;
		11781: rom = 27;
		11782: rom = 27;
		11783: rom = 27;
		11784: rom = 27;
		11785: rom = 27;
		11786: rom = 27;
		11787: rom = 27;
		11788: rom = 27;
		11789: rom = 27;
		11790: rom = 27;
		11791: rom = 27;
		11792: rom = 27;
		11793: rom = 27;
		11794: rom = 27;
		11795: rom = 27;
		11796: rom = 27;
		11797: rom = 27;
		11798: rom = 27;
		11799: rom = 27;
		11800: rom = 27;
		11801: rom = 27;
		11802: rom = 27;
		11803: rom = 27;
		11804: rom = 27;
		11805: rom = 27;
		11806: rom = 27;
		11807: rom = 27;
		11808: rom = 27;
		11809: rom = 27;
		11810: rom = 27;
		11811: rom = 27;
		11812: rom = 27;
		11813: rom = 27;
		11814: rom = 27;
		11815: rom = 27;
		11816: rom = 27;
		11817: rom = 27;
		11818: rom = 27;
		11819: rom = 27;
		11820: rom = 27;
		11821: rom = 27;
		11822: rom = 27;
		11823: rom = 27;
		11824: rom = 27;
		11825: rom = 27;
		11826: rom = 27;
		11827: rom = 27;
		11828: rom = 27;
		11829: rom = 27;
		11830: rom = 27;
		11831: rom = 27;
		11832: rom = 27;
		11833: rom = 27;
		11834: rom = 27;
		11835: rom = 27;
		11836: rom = 27;
		11837: rom = 27;
		11838: rom = 27;
		11839: rom = 27;
		11840: rom = 27;
		11841: rom = 27;
		11842: rom = 27;
		11843: rom = 17;
		11844: rom = 18;
		11845: rom = 18;
		11846: rom = 18;
		11847: rom = 18;
		11848: rom = 18;
		11849: rom = 18;
		11850: rom = 18;
		11851: rom = 18;
		11852: rom = 18;
		11853: rom = 18;
		11854: rom = 18;
		11855: rom = 18;
		11856: rom = 18;
		11857: rom = 18;
		11858: rom = 18;
		11859: rom = 11;
		11860: rom = 18;
		11861: rom = 18;
		11862: rom = 18;
		11863: rom = 18;
		11864: rom = 18;
		11865: rom = 18;
		11866: rom = 18;
		11867: rom = 18;
		11868: rom = 13;
		11869: rom = 15;
		11870: rom = 18;
		11871: rom = 18;
		11872: rom = 18;
		11873: rom = 18;
		11874: rom = 18;
		11875: rom = 18;
		11876: rom = 18;
		11877: rom = 18;
		11878: rom = 18;
		11879: rom = 18;
		11880: rom = 18;
		11881: rom = 18;
		11882: rom = 18;
		11883: rom = 18;
		11884: rom = 18;
		11885: rom = 11;
		11886: rom = 27;
		11887: rom = 27;
		11888: rom = 27;
		11889: rom = 27;
		11890: rom = 27;
		11891: rom = 27;
		11892: rom = 27;
		11893: rom = 27;
		11894: rom = 27;
		11895: rom = 27;
		11896: rom = 27;
		11897: rom = 27;
		11898: rom = 27;
		11904: rom = 27;
		11905: rom = 27;
		11906: rom = 27;
		11907: rom = 27;
		11908: rom = 0;
		11909: rom = 0;
		11910: rom = 0;
		11911: rom = 0;
		11912: rom = 0;
		11913: rom = 0;
		11914: rom = 0;
		11915: rom = 0;
		11916: rom = 0;
		11917: rom = 0;
		11918: rom = 0;
		11919: rom = 0;
		11920: rom = 27;
		11921: rom = 27;
		11922: rom = 27;
		11923: rom = 27;
		11924: rom = 27;
		11925: rom = 27;
		11926: rom = 27;
		11927: rom = 27;
		11928: rom = 27;
		11929: rom = 27;
		11930: rom = 27;
		11931: rom = 27;
		11932: rom = 27;
		11933: rom = 27;
		11934: rom = 27;
		11935: rom = 27;
		11936: rom = 27;
		11937: rom = 27;
		11938: rom = 27;
		11939: rom = 27;
		11940: rom = 27;
		11941: rom = 27;
		11942: rom = 27;
		11943: rom = 27;
		11944: rom = 27;
		11945: rom = 27;
		11946: rom = 27;
		11947: rom = 27;
		11948: rom = 27;
		11949: rom = 27;
		11950: rom = 27;
		11951: rom = 27;
		11952: rom = 27;
		11953: rom = 27;
		11954: rom = 27;
		11955: rom = 27;
		11956: rom = 27;
		11957: rom = 27;
		11958: rom = 27;
		11959: rom = 27;
		11960: rom = 27;
		11961: rom = 27;
		11962: rom = 27;
		11963: rom = 27;
		11964: rom = 27;
		11965: rom = 27;
		11966: rom = 27;
		11967: rom = 27;
		11968: rom = 27;
		11969: rom = 27;
		11970: rom = 27;
		11971: rom = 23;
		11972: rom = 14;
		11973: rom = 18;
		11974: rom = 18;
		11975: rom = 18;
		11976: rom = 18;
		11977: rom = 18;
		11978: rom = 18;
		11979: rom = 18;
		11980: rom = 18;
		11981: rom = 18;
		11982: rom = 18;
		11983: rom = 18;
		11984: rom = 18;
		11985: rom = 18;
		11986: rom = 18;
		11987: rom = 16;
		11988: rom = 14;
		11989: rom = 18;
		11990: rom = 18;
		11991: rom = 18;
		11992: rom = 18;
		11993: rom = 18;
		11994: rom = 18;
		11995: rom = 18;
		11996: rom = 18;
		11997: rom = 10;
		11998: rom = 17;
		11999: rom = 18;
		12000: rom = 18;
		12001: rom = 18;
		12002: rom = 18;
		12003: rom = 18;
		12004: rom = 18;
		12005: rom = 18;
		12006: rom = 18;
		12007: rom = 18;
		12008: rom = 18;
		12009: rom = 18;
		12010: rom = 18;
		12011: rom = 18;
		12012: rom = 18;
		12013: rom = 13;
		12014: rom = 25;
		12015: rom = 27;
		12016: rom = 27;
		12017: rom = 27;
		12018: rom = 27;
		12019: rom = 27;
		12020: rom = 27;
		12021: rom = 27;
		12022: rom = 27;
		12023: rom = 27;
		12024: rom = 27;
		12025: rom = 27;
		12026: rom = 27;
		12032: rom = 27;
		12033: rom = 27;
		12034: rom = 27;
		12035: rom = 27;
		12036: rom = 0;
		12037: rom = 0;
		12038: rom = 0;
		12039: rom = 0;
		12040: rom = 0;
		12041: rom = 0;
		12042: rom = 0;
		12043: rom = 0;
		12044: rom = 0;
		12045: rom = 0;
		12046: rom = 0;
		12047: rom = 0;
		12048: rom = 27;
		12049: rom = 27;
		12050: rom = 27;
		12051: rom = 27;
		12052: rom = 27;
		12053: rom = 27;
		12054: rom = 27;
		12055: rom = 27;
		12056: rom = 27;
		12057: rom = 27;
		12058: rom = 27;
		12059: rom = 27;
		12060: rom = 27;
		12061: rom = 27;
		12062: rom = 27;
		12063: rom = 27;
		12064: rom = 27;
		12065: rom = 27;
		12066: rom = 27;
		12067: rom = 27;
		12068: rom = 27;
		12069: rom = 27;
		12070: rom = 27;
		12071: rom = 27;
		12072: rom = 27;
		12073: rom = 27;
		12074: rom = 27;
		12075: rom = 27;
		12076: rom = 27;
		12077: rom = 27;
		12078: rom = 27;
		12079: rom = 27;
		12080: rom = 27;
		12081: rom = 27;
		12082: rom = 27;
		12083: rom = 27;
		12084: rom = 27;
		12085: rom = 27;
		12086: rom = 27;
		12087: rom = 27;
		12088: rom = 27;
		12089: rom = 27;
		12090: rom = 27;
		12091: rom = 27;
		12092: rom = 27;
		12093: rom = 27;
		12094: rom = 27;
		12095: rom = 27;
		12096: rom = 27;
		12097: rom = 27;
		12098: rom = 27;
		12099: rom = 27;
		12100: rom = 13;
		12101: rom = 18;
		12102: rom = 18;
		12103: rom = 18;
		12104: rom = 18;
		12105: rom = 18;
		12106: rom = 18;
		12107: rom = 18;
		12108: rom = 18;
		12109: rom = 18;
		12110: rom = 18;
		12111: rom = 18;
		12112: rom = 18;
		12113: rom = 18;
		12114: rom = 18;
		12115: rom = 18;
		12116: rom = 12;
		12117: rom = 17;
		12118: rom = 18;
		12119: rom = 18;
		12120: rom = 18;
		12121: rom = 18;
		12122: rom = 18;
		12123: rom = 18;
		12124: rom = 18;
		12125: rom = 14;
		12126: rom = 14;
		12127: rom = 18;
		12128: rom = 18;
		12129: rom = 18;
		12130: rom = 18;
		12131: rom = 18;
		12132: rom = 18;
		12133: rom = 18;
		12134: rom = 18;
		12135: rom = 18;
		12136: rom = 18;
		12137: rom = 18;
		12138: rom = 18;
		12139: rom = 18;
		12140: rom = 18;
		12141: rom = 15;
		12142: rom = 21;
		12143: rom = 27;
		12144: rom = 27;
		12145: rom = 27;
		12146: rom = 27;
		12147: rom = 27;
		12148: rom = 27;
		12149: rom = 27;
		12150: rom = 27;
		12151: rom = 27;
		12152: rom = 27;
		12153: rom = 27;
		12154: rom = 27;
		12160: rom = 27;
		12161: rom = 27;
		12162: rom = 27;
		12163: rom = 27;
		12164: rom = 27;
		12165: rom = 27;
		12166: rom = 27;
		12167: rom = 27;
		12168: rom = 27;
		12169: rom = 27;
		12170: rom = 27;
		12171: rom = 27;
		12172: rom = 27;
		12173: rom = 27;
		12174: rom = 8;
		12175: rom = 0;
		12176: rom = 27;
		12177: rom = 27;
		12178: rom = 27;
		12179: rom = 27;
		12180: rom = 27;
		12181: rom = 27;
		12182: rom = 27;
		12183: rom = 27;
		12184: rom = 27;
		12185: rom = 27;
		12186: rom = 27;
		12187: rom = 27;
		12188: rom = 27;
		12189: rom = 27;
		12190: rom = 27;
		12191: rom = 27;
		12192: rom = 27;
		12193: rom = 27;
		12194: rom = 27;
		12195: rom = 27;
		12196: rom = 27;
		12197: rom = 27;
		12198: rom = 27;
		12199: rom = 27;
		12200: rom = 27;
		12201: rom = 27;
		12202: rom = 27;
		12203: rom = 27;
		12204: rom = 27;
		12205: rom = 27;
		12206: rom = 27;
		12207: rom = 27;
		12208: rom = 27;
		12209: rom = 27;
		12210: rom = 27;
		12211: rom = 27;
		12212: rom = 27;
		12213: rom = 27;
		12214: rom = 27;
		12215: rom = 27;
		12216: rom = 27;
		12217: rom = 27;
		12218: rom = 27;
		12219: rom = 27;
		12220: rom = 27;
		12221: rom = 27;
		12222: rom = 27;
		12223: rom = 27;
		12224: rom = 27;
		12225: rom = 27;
		12226: rom = 27;
		12227: rom = 27;
		12228: rom = 24;
		12229: rom = 11;
		12230: rom = 18;
		12231: rom = 18;
		12232: rom = 18;
		12233: rom = 18;
		12234: rom = 18;
		12235: rom = 18;
		12236: rom = 18;
		12237: rom = 18;
		12238: rom = 18;
		12239: rom = 18;
		12240: rom = 18;
		12241: rom = 18;
		12242: rom = 18;
		12243: rom = 18;
		12244: rom = 16;
		12245: rom = 12;
		12246: rom = 9;
		12247: rom = 14;
		12248: rom = 18;
		12249: rom = 18;
		12250: rom = 18;
		12251: rom = 18;
		12252: rom = 18;
		12253: rom = 18;
		12254: rom = 10;
		12255: rom = 18;
		12256: rom = 18;
		12257: rom = 18;
		12258: rom = 18;
		12259: rom = 18;
		12260: rom = 18;
		12261: rom = 18;
		12262: rom = 18;
		12263: rom = 18;
		12264: rom = 18;
		12265: rom = 18;
		12266: rom = 18;
		12267: rom = 18;
		12268: rom = 18;
		12269: rom = 17;
		12270: rom = 18;
		12271: rom = 27;
		12272: rom = 27;
		12273: rom = 27;
		12274: rom = 27;
		12275: rom = 27;
		12276: rom = 27;
		12277: rom = 27;
		12278: rom = 27;
		12279: rom = 27;
		12280: rom = 27;
		12281: rom = 27;
		12282: rom = 27;
		12288: rom = 27;
		12289: rom = 27;
		12290: rom = 27;
		12291: rom = 27;
		12292: rom = 27;
		12293: rom = 27;
		12294: rom = 27;
		12295: rom = 27;
		12296: rom = 27;
		12297: rom = 27;
		12298: rom = 27;
		12299: rom = 27;
		12300: rom = 27;
		12301: rom = 27;
		12302: rom = 8;
		12303: rom = 0;
		12304: rom = 27;
		12305: rom = 27;
		12306: rom = 27;
		12307: rom = 27;
		12308: rom = 27;
		12309: rom = 27;
		12310: rom = 27;
		12311: rom = 27;
		12312: rom = 27;
		12313: rom = 27;
		12314: rom = 27;
		12315: rom = 27;
		12316: rom = 27;
		12317: rom = 27;
		12318: rom = 27;
		12319: rom = 27;
		12320: rom = 27;
		12321: rom = 27;
		12322: rom = 27;
		12323: rom = 27;
		12324: rom = 27;
		12325: rom = 27;
		12326: rom = 27;
		12327: rom = 27;
		12328: rom = 27;
		12329: rom = 27;
		12330: rom = 27;
		12331: rom = 27;
		12332: rom = 27;
		12333: rom = 27;
		12334: rom = 27;
		12335: rom = 27;
		12336: rom = 27;
		12337: rom = 27;
		12338: rom = 27;
		12339: rom = 27;
		12340: rom = 27;
		12341: rom = 27;
		12342: rom = 27;
		12343: rom = 27;
		12344: rom = 27;
		12345: rom = 27;
		12346: rom = 27;
		12347: rom = 27;
		12348: rom = 27;
		12349: rom = 27;
		12350: rom = 27;
		12351: rom = 27;
		12352: rom = 27;
		12353: rom = 27;
		12354: rom = 27;
		12355: rom = 27;
		12356: rom = 27;
		12357: rom = 22;
		12358: rom = 12;
		12359: rom = 15;
		12360: rom = 18;
		12361: rom = 18;
		12362: rom = 18;
		12363: rom = 18;
		12364: rom = 18;
		12365: rom = 18;
		12366: rom = 18;
		12367: rom = 18;
		12368: rom = 18;
		12369: rom = 18;
		12370: rom = 18;
		12371: rom = 18;
		12372: rom = 18;
		12373: rom = 18;
		12374: rom = 18;
		12375: rom = 14;
		12376: rom = 12;
		12377: rom = 18;
		12378: rom = 18;
		12379: rom = 18;
		12380: rom = 18;
		12381: rom = 18;
		12382: rom = 14;
		12383: rom = 15;
		12384: rom = 18;
		12385: rom = 18;
		12386: rom = 18;
		12387: rom = 18;
		12388: rom = 18;
		12389: rom = 18;
		12390: rom = 18;
		12391: rom = 18;
		12392: rom = 18;
		12393: rom = 18;
		12394: rom = 18;
		12395: rom = 18;
		12396: rom = 18;
		12397: rom = 18;
		12398: rom = 15;
		12399: rom = 27;
		12400: rom = 27;
		12401: rom = 27;
		12402: rom = 27;
		12403: rom = 27;
		12404: rom = 27;
		12405: rom = 27;
		12406: rom = 27;
		12407: rom = 27;
		12408: rom = 27;
		12409: rom = 27;
		12410: rom = 27;
		12416: rom = 27;
		12417: rom = 27;
		12418: rom = 27;
		12419: rom = 27;
		12420: rom = 27;
		12421: rom = 27;
		12422: rom = 27;
		12423: rom = 27;
		12424: rom = 27;
		12425: rom = 27;
		12426: rom = 27;
		12427: rom = 27;
		12428: rom = 27;
		12429: rom = 27;
		12430: rom = 8;
		12431: rom = 0;
		12432: rom = 27;
		12433: rom = 27;
		12434: rom = 27;
		12435: rom = 27;
		12436: rom = 27;
		12437: rom = 27;
		12438: rom = 27;
		12439: rom = 27;
		12440: rom = 27;
		12441: rom = 27;
		12442: rom = 27;
		12443: rom = 27;
		12444: rom = 27;
		12445: rom = 27;
		12446: rom = 27;
		12447: rom = 27;
		12448: rom = 27;
		12449: rom = 27;
		12450: rom = 27;
		12451: rom = 27;
		12452: rom = 27;
		12453: rom = 27;
		12454: rom = 27;
		12455: rom = 27;
		12456: rom = 27;
		12457: rom = 27;
		12458: rom = 27;
		12459: rom = 27;
		12460: rom = 27;
		12461: rom = 27;
		12462: rom = 27;
		12463: rom = 27;
		12464: rom = 27;
		12465: rom = 27;
		12466: rom = 27;
		12467: rom = 27;
		12468: rom = 27;
		12469: rom = 27;
		12470: rom = 27;
		12471: rom = 27;
		12472: rom = 27;
		12473: rom = 27;
		12474: rom = 27;
		12475: rom = 27;
		12476: rom = 27;
		12477: rom = 27;
		12478: rom = 27;
		12479: rom = 27;
		12480: rom = 27;
		12481: rom = 27;
		12482: rom = 27;
		12483: rom = 27;
		12484: rom = 27;
		12485: rom = 27;
		12486: rom = 27;
		12487: rom = 21;
		12488: rom = 13;
		12489: rom = 12;
		12490: rom = 15;
		12491: rom = 17;
		12492: rom = 18;
		12493: rom = 18;
		12494: rom = 18;
		12495: rom = 18;
		12496: rom = 18;
		12497: rom = 18;
		12498: rom = 18;
		12499: rom = 18;
		12500: rom = 18;
		12501: rom = 18;
		12502: rom = 18;
		12503: rom = 18;
		12504: rom = 13;
		12505: rom = 16;
		12506: rom = 18;
		12507: rom = 18;
		12508: rom = 18;
		12509: rom = 18;
		12510: rom = 18;
		12511: rom = 11;
		12512: rom = 18;
		12513: rom = 18;
		12514: rom = 18;
		12515: rom = 18;
		12516: rom = 18;
		12517: rom = 18;
		12518: rom = 18;
		12519: rom = 18;
		12520: rom = 18;
		12521: rom = 18;
		12522: rom = 18;
		12523: rom = 18;
		12524: rom = 18;
		12525: rom = 18;
		12526: rom = 11;
		12527: rom = 27;
		12528: rom = 27;
		12529: rom = 27;
		12530: rom = 27;
		12531: rom = 27;
		12532: rom = 27;
		12533: rom = 27;
		12534: rom = 27;
		12535: rom = 27;
		12536: rom = 27;
		12537: rom = 27;
		12538: rom = 27;
		12544: rom = 27;
		12545: rom = 27;
		12546: rom = 27;
		12547: rom = 27;
		12548: rom = 27;
		12549: rom = 27;
		12550: rom = 27;
		12551: rom = 27;
		12552: rom = 27;
		12553: rom = 27;
		12554: rom = 27;
		12555: rom = 27;
		12556: rom = 27;
		12557: rom = 27;
		12558: rom = 8;
		12559: rom = 0;
		12560: rom = 27;
		12561: rom = 27;
		12562: rom = 27;
		12563: rom = 27;
		12564: rom = 27;
		12565: rom = 27;
		12566: rom = 27;
		12567: rom = 27;
		12568: rom = 27;
		12569: rom = 27;
		12570: rom = 27;
		12571: rom = 27;
		12572: rom = 27;
		12573: rom = 27;
		12574: rom = 27;
		12575: rom = 27;
		12576: rom = 27;
		12577: rom = 27;
		12578: rom = 27;
		12579: rom = 27;
		12580: rom = 27;
		12581: rom = 27;
		12582: rom = 27;
		12583: rom = 27;
		12584: rom = 27;
		12585: rom = 27;
		12586: rom = 27;
		12587: rom = 27;
		12588: rom = 27;
		12589: rom = 27;
		12590: rom = 27;
		12591: rom = 27;
		12592: rom = 27;
		12593: rom = 27;
		12594: rom = 27;
		12595: rom = 27;
		12596: rom = 27;
		12597: rom = 27;
		12598: rom = 27;
		12599: rom = 27;
		12600: rom = 27;
		12601: rom = 27;
		12602: rom = 27;
		12603: rom = 27;
		12604: rom = 27;
		12605: rom = 27;
		12606: rom = 27;
		12607: rom = 27;
		12608: rom = 27;
		12609: rom = 27;
		12610: rom = 27;
		12611: rom = 27;
		12612: rom = 27;
		12613: rom = 27;
		12614: rom = 27;
		12615: rom = 27;
		12616: rom = 27;
		12617: rom = 25;
		12618: rom = 21;
		12619: rom = 17;
		12620: rom = 13;
		12621: rom = 11;
		12622: rom = 12;
		12623: rom = 13;
		12624: rom = 14;
		12625: rom = 18;
		12626: rom = 18;
		12627: rom = 18;
		12628: rom = 18;
		12629: rom = 18;
		12630: rom = 18;
		12631: rom = 18;
		12632: rom = 18;
		12633: rom = 12;
		12634: rom = 18;
		12635: rom = 18;
		12636: rom = 18;
		12637: rom = 18;
		12638: rom = 18;
		12639: rom = 11;
		12640: rom = 17;
		12641: rom = 18;
		12642: rom = 18;
		12643: rom = 18;
		12644: rom = 18;
		12645: rom = 18;
		12646: rom = 18;
		12647: rom = 18;
		12648: rom = 18;
		12649: rom = 18;
		12650: rom = 18;
		12651: rom = 18;
		12652: rom = 18;
		12653: rom = 18;
		12654: rom = 12;
		12655: rom = 26;
		12656: rom = 27;
		12657: rom = 27;
		12658: rom = 27;
		12659: rom = 27;
		12660: rom = 27;
		12661: rom = 27;
		12662: rom = 27;
		12663: rom = 27;
		12664: rom = 27;
		12665: rom = 27;
		12666: rom = 27;
		12672: rom = 27;
		12673: rom = 27;
		12674: rom = 27;
		12675: rom = 27;
		12676: rom = 27;
		12677: rom = 27;
		12678: rom = 27;
		12679: rom = 27;
		12680: rom = 27;
		12681: rom = 27;
		12682: rom = 27;
		12683: rom = 27;
		12684: rom = 27;
		12685: rom = 27;
		12686: rom = 8;
		12687: rom = 0;
		12688: rom = 27;
		12689: rom = 27;
		12690: rom = 27;
		12691: rom = 27;
		12692: rom = 27;
		12693: rom = 27;
		12694: rom = 27;
		12695: rom = 27;
		12696: rom = 27;
		12697: rom = 27;
		12698: rom = 27;
		12699: rom = 27;
		12700: rom = 27;
		12701: rom = 27;
		12702: rom = 27;
		12703: rom = 27;
		12704: rom = 27;
		12705: rom = 27;
		12706: rom = 27;
		12707: rom = 27;
		12708: rom = 27;
		12709: rom = 27;
		12710: rom = 27;
		12711: rom = 27;
		12712: rom = 27;
		12713: rom = 27;
		12714: rom = 27;
		12715: rom = 27;
		12716: rom = 27;
		12717: rom = 27;
		12718: rom = 27;
		12719: rom = 27;
		12720: rom = 27;
		12721: rom = 27;
		12722: rom = 27;
		12723: rom = 27;
		12724: rom = 27;
		12725: rom = 27;
		12726: rom = 27;
		12727: rom = 27;
		12728: rom = 27;
		12729: rom = 27;
		12730: rom = 27;
		12731: rom = 27;
		12732: rom = 27;
		12733: rom = 27;
		12734: rom = 27;
		12735: rom = 27;
		12736: rom = 27;
		12737: rom = 27;
		12738: rom = 27;
		12739: rom = 27;
		12740: rom = 27;
		12741: rom = 27;
		12742: rom = 27;
		12743: rom = 27;
		12744: rom = 27;
		12745: rom = 27;
		12746: rom = 27;
		12747: rom = 27;
		12748: rom = 27;
		12749: rom = 27;
		12750: rom = 25;
		12751: rom = 23;
		12752: rom = 17;
		12753: rom = 16;
		12754: rom = 18;
		12755: rom = 18;
		12756: rom = 18;
		12757: rom = 18;
		12758: rom = 18;
		12759: rom = 18;
		12760: rom = 18;
		12761: rom = 11;
		12762: rom = 18;
		12763: rom = 18;
		12764: rom = 18;
		12765: rom = 18;
		12766: rom = 18;
		12767: rom = 15;
		12768: rom = 14;
		12769: rom = 18;
		12770: rom = 18;
		12771: rom = 18;
		12772: rom = 18;
		12773: rom = 18;
		12774: rom = 18;
		12775: rom = 18;
		12776: rom = 18;
		12777: rom = 18;
		12778: rom = 18;
		12779: rom = 18;
		12780: rom = 18;
		12781: rom = 18;
		12782: rom = 14;
		12783: rom = 24;
		12784: rom = 27;
		12785: rom = 27;
		12786: rom = 27;
		12787: rom = 27;
		12788: rom = 27;
		12789: rom = 27;
		12790: rom = 27;
		12791: rom = 27;
		12792: rom = 27;
		12793: rom = 27;
		12794: rom = 27;
		12800: rom = 27;
		12801: rom = 27;
		12802: rom = 27;
		12803: rom = 27;
		12804: rom = 27;
		12805: rom = 27;
		12806: rom = 27;
		12807: rom = 27;
		12808: rom = 27;
		12809: rom = 27;
		12810: rom = 27;
		12811: rom = 27;
		12812: rom = 27;
		12813: rom = 27;
		12814: rom = 8;
		12815: rom = 0;
		12816: rom = 27;
		12817: rom = 27;
		12818: rom = 27;
		12819: rom = 27;
		12820: rom = 27;
		12821: rom = 27;
		12822: rom = 27;
		12823: rom = 27;
		12824: rom = 27;
		12825: rom = 27;
		12826: rom = 27;
		12827: rom = 27;
		12828: rom = 27;
		12829: rom = 27;
		12830: rom = 27;
		12831: rom = 27;
		12832: rom = 27;
		12833: rom = 27;
		12834: rom = 27;
		12835: rom = 27;
		12836: rom = 27;
		12837: rom = 27;
		12838: rom = 27;
		12839: rom = 27;
		12840: rom = 27;
		12841: rom = 27;
		12842: rom = 27;
		12843: rom = 27;
		12844: rom = 27;
		12845: rom = 27;
		12846: rom = 27;
		12847: rom = 27;
		12848: rom = 27;
		12849: rom = 27;
		12850: rom = 27;
		12851: rom = 27;
		12852: rom = 27;
		12853: rom = 27;
		12854: rom = 27;
		12855: rom = 27;
		12856: rom = 27;
		12857: rom = 27;
		12858: rom = 27;
		12859: rom = 27;
		12860: rom = 27;
		12861: rom = 27;
		12862: rom = 27;
		12863: rom = 27;
		12864: rom = 27;
		12865: rom = 27;
		12866: rom = 27;
		12867: rom = 27;
		12868: rom = 27;
		12869: rom = 27;
		12870: rom = 27;
		12871: rom = 27;
		12872: rom = 27;
		12873: rom = 27;
		12874: rom = 27;
		12875: rom = 27;
		12876: rom = 27;
		12877: rom = 27;
		12878: rom = 27;
		12879: rom = 27;
		12880: rom = 22;
		12881: rom = 15;
		12882: rom = 18;
		12883: rom = 18;
		12884: rom = 18;
		12885: rom = 18;
		12886: rom = 18;
		12887: rom = 18;
		12888: rom = 18;
		12889: rom = 13;
		12890: rom = 17;
		12891: rom = 18;
		12892: rom = 18;
		12893: rom = 18;
		12894: rom = 18;
		12895: rom = 18;
		12896: rom = 11;
		12897: rom = 18;
		12898: rom = 18;
		12899: rom = 18;
		12900: rom = 18;
		12901: rom = 18;
		12902: rom = 18;
		12903: rom = 18;
		12904: rom = 18;
		12905: rom = 18;
		12906: rom = 18;
		12907: rom = 18;
		12908: rom = 18;
		12909: rom = 18;
		12910: rom = 15;
		12911: rom = 22;
		12912: rom = 27;
		12913: rom = 27;
		12914: rom = 27;
		12915: rom = 27;
		12916: rom = 27;
		12917: rom = 27;
		12918: rom = 27;
		12919: rom = 27;
		12920: rom = 27;
		12921: rom = 27;
		12922: rom = 27;
		12928: rom = 27;
		12929: rom = 27;
		12930: rom = 27;
		12931: rom = 27;
		12932: rom = 27;
		12933: rom = 27;
		12934: rom = 27;
		12935: rom = 27;
		12936: rom = 27;
		12937: rom = 27;
		12938: rom = 27;
		12939: rom = 27;
		12940: rom = 27;
		12941: rom = 27;
		12942: rom = 24;
		12943: rom = 22;
		12944: rom = 27;
		12945: rom = 27;
		12946: rom = 27;
		12947: rom = 27;
		12948: rom = 27;
		12949: rom = 27;
		12950: rom = 27;
		12951: rom = 27;
		12952: rom = 27;
		12953: rom = 27;
		12954: rom = 27;
		12955: rom = 27;
		12956: rom = 27;
		12957: rom = 27;
		12958: rom = 27;
		12959: rom = 27;
		12960: rom = 27;
		12961: rom = 27;
		12962: rom = 27;
		12963: rom = 27;
		12964: rom = 27;
		12965: rom = 27;
		12966: rom = 27;
		12967: rom = 27;
		12968: rom = 27;
		12969: rom = 27;
		12970: rom = 27;
		12971: rom = 27;
		12972: rom = 27;
		12973: rom = 27;
		12974: rom = 27;
		12975: rom = 27;
		12976: rom = 27;
		12977: rom = 27;
		12978: rom = 27;
		12979: rom = 27;
		12980: rom = 27;
		12981: rom = 27;
		12982: rom = 27;
		12983: rom = 27;
		12984: rom = 27;
		12985: rom = 27;
		12986: rom = 27;
		12987: rom = 27;
		12988: rom = 27;
		12989: rom = 27;
		12990: rom = 27;
		12991: rom = 27;
		12992: rom = 27;
		12993: rom = 27;
		12994: rom = 27;
		12995: rom = 27;
		12996: rom = 27;
		12997: rom = 27;
		12998: rom = 27;
		12999: rom = 27;
		13000: rom = 27;
		13001: rom = 27;
		13002: rom = 27;
		13003: rom = 27;
		13004: rom = 27;
		13005: rom = 27;
		13006: rom = 27;
		13007: rom = 27;
		13008: rom = 23;
		13009: rom = 14;
		13010: rom = 18;
		13011: rom = 18;
		13012: rom = 18;
		13013: rom = 18;
		13014: rom = 18;
		13015: rom = 18;
		13016: rom = 18;
		13017: rom = 15;
		13018: rom = 15;
		13019: rom = 18;
		13020: rom = 18;
		13021: rom = 18;
		13022: rom = 18;
		13023: rom = 18;
		13024: rom = 11;
		13025: rom = 18;
		13026: rom = 18;
		13027: rom = 18;
		13028: rom = 18;
		13029: rom = 18;
		13030: rom = 18;
		13031: rom = 18;
		13032: rom = 18;
		13033: rom = 18;
		13034: rom = 18;
		13035: rom = 18;
		13036: rom = 18;
		13037: rom = 18;
		13038: rom = 16;
		13039: rom = 20;
		13040: rom = 27;
		13041: rom = 27;
		13042: rom = 27;
		13043: rom = 27;
		13044: rom = 27;
		13045: rom = 27;
		13046: rom = 27;
		13047: rom = 27;
		13048: rom = 27;
		13049: rom = 27;
		13050: rom = 27;
		13056: rom = 27;
		13057: rom = 27;
		13058: rom = 27;
		13059: rom = 27;
		13060: rom = 27;
		13061: rom = 27;
		13062: rom = 27;
		13063: rom = 27;
		13064: rom = 27;
		13065: rom = 27;
		13066: rom = 27;
		13067: rom = 27;
		13068: rom = 27;
		13069: rom = 27;
		13070: rom = 27;
		13071: rom = 27;
		13072: rom = 27;
		13073: rom = 27;
		13074: rom = 27;
		13075: rom = 27;
		13076: rom = 27;
		13077: rom = 27;
		13078: rom = 27;
		13079: rom = 27;
		13080: rom = 27;
		13081: rom = 27;
		13082: rom = 27;
		13083: rom = 27;
		13084: rom = 27;
		13085: rom = 27;
		13086: rom = 27;
		13087: rom = 27;
		13088: rom = 27;
		13089: rom = 27;
		13090: rom = 27;
		13091: rom = 27;
		13092: rom = 27;
		13093: rom = 27;
		13094: rom = 27;
		13095: rom = 27;
		13096: rom = 27;
		13097: rom = 27;
		13098: rom = 27;
		13099: rom = 27;
		13100: rom = 27;
		13101: rom = 27;
		13102: rom = 27;
		13103: rom = 27;
		13104: rom = 27;
		13105: rom = 27;
		13106: rom = 27;
		13107: rom = 27;
		13108: rom = 27;
		13109: rom = 27;
		13110: rom = 27;
		13111: rom = 27;
		13112: rom = 27;
		13113: rom = 27;
		13114: rom = 27;
		13115: rom = 27;
		13116: rom = 27;
		13117: rom = 27;
		13118: rom = 27;
		13119: rom = 27;
		13120: rom = 27;
		13121: rom = 27;
		13122: rom = 27;
		13123: rom = 27;
		13124: rom = 27;
		13125: rom = 27;
		13126: rom = 27;
		13127: rom = 27;
		13128: rom = 27;
		13129: rom = 27;
		13130: rom = 27;
		13131: rom = 27;
		13132: rom = 27;
		13133: rom = 27;
		13134: rom = 27;
		13135: rom = 27;
		13136: rom = 22;
		13137: rom = 16;
		13138: rom = 18;
		13139: rom = 18;
		13140: rom = 18;
		13141: rom = 18;
		13142: rom = 18;
		13143: rom = 18;
		13144: rom = 18;
		13145: rom = 17;
		13146: rom = 13;
		13147: rom = 18;
		13148: rom = 18;
		13149: rom = 18;
		13150: rom = 18;
		13151: rom = 18;
		13152: rom = 13;
		13153: rom = 16;
		13154: rom = 18;
		13155: rom = 18;
		13156: rom = 18;
		13157: rom = 18;
		13158: rom = 18;
		13159: rom = 18;
		13160: rom = 18;
		13161: rom = 18;
		13162: rom = 18;
		13163: rom = 18;
		13164: rom = 18;
		13165: rom = 18;
		13166: rom = 17;
		13167: rom = 18;
		13168: rom = 27;
		13169: rom = 27;
		13170: rom = 27;
		13171: rom = 27;
		13172: rom = 27;
		13173: rom = 27;
		13174: rom = 27;
		13175: rom = 27;
		13176: rom = 27;
		13177: rom = 27;
		13178: rom = 27;
		13184: rom = 27;
		13185: rom = 27;
		13186: rom = 27;
		13187: rom = 27;
		13188: rom = 17;
		13189: rom = 17;
		13190: rom = 17;
		13191: rom = 17;
		13192: rom = 17;
		13193: rom = 17;
		13194: rom = 17;
		13195: rom = 17;
		13196: rom = 17;
		13197: rom = 17;
		13198: rom = 17;
		13199: rom = 20;
		13200: rom = 27;
		13201: rom = 27;
		13202: rom = 27;
		13203: rom = 27;
		13204: rom = 27;
		13205: rom = 27;
		13206: rom = 27;
		13207: rom = 27;
		13208: rom = 27;
		13209: rom = 27;
		13210: rom = 27;
		13211: rom = 27;
		13212: rom = 27;
		13213: rom = 27;
		13214: rom = 27;
		13215: rom = 27;
		13216: rom = 27;
		13217: rom = 27;
		13218: rom = 27;
		13219: rom = 27;
		13220: rom = 27;
		13221: rom = 27;
		13222: rom = 27;
		13223: rom = 27;
		13224: rom = 27;
		13225: rom = 27;
		13226: rom = 27;
		13227: rom = 27;
		13228: rom = 27;
		13229: rom = 27;
		13230: rom = 27;
		13231: rom = 27;
		13232: rom = 27;
		13233: rom = 27;
		13234: rom = 27;
		13235: rom = 27;
		13236: rom = 27;
		13237: rom = 27;
		13238: rom = 27;
		13239: rom = 27;
		13240: rom = 27;
		13241: rom = 27;
		13242: rom = 27;
		13243: rom = 27;
		13244: rom = 27;
		13245: rom = 27;
		13246: rom = 27;
		13247: rom = 27;
		13248: rom = 27;
		13249: rom = 27;
		13250: rom = 27;
		13251: rom = 27;
		13252: rom = 27;
		13253: rom = 27;
		13254: rom = 27;
		13255: rom = 27;
		13256: rom = 27;
		13257: rom = 27;
		13258: rom = 27;
		13259: rom = 27;
		13260: rom = 27;
		13261: rom = 27;
		13262: rom = 27;
		13263: rom = 27;
		13264: rom = 21;
		13265: rom = 16;
		13266: rom = 18;
		13267: rom = 18;
		13268: rom = 18;
		13269: rom = 18;
		13270: rom = 18;
		13271: rom = 18;
		13272: rom = 18;
		13273: rom = 18;
		13274: rom = 12;
		13275: rom = 18;
		13276: rom = 18;
		13277: rom = 18;
		13278: rom = 18;
		13279: rom = 18;
		13280: rom = 16;
		13281: rom = 14;
		13282: rom = 18;
		13283: rom = 18;
		13284: rom = 18;
		13285: rom = 18;
		13286: rom = 18;
		13287: rom = 18;
		13288: rom = 18;
		13289: rom = 18;
		13290: rom = 18;
		13291: rom = 18;
		13292: rom = 18;
		13293: rom = 18;
		13294: rom = 18;
		13295: rom = 17;
		13296: rom = 27;
		13297: rom = 27;
		13298: rom = 27;
		13299: rom = 27;
		13300: rom = 27;
		13301: rom = 27;
		13302: rom = 27;
		13303: rom = 27;
		13304: rom = 27;
		13305: rom = 27;
		13306: rom = 27;
		13312: rom = 27;
		13313: rom = 27;
		13314: rom = 27;
		13315: rom = 27;
		13316: rom = 0;
		13317: rom = 0;
		13318: rom = 0;
		13319: rom = 0;
		13320: rom = 0;
		13321: rom = 0;
		13322: rom = 0;
		13323: rom = 0;
		13324: rom = 0;
		13325: rom = 0;
		13326: rom = 0;
		13327: rom = 14;
		13328: rom = 27;
		13329: rom = 27;
		13330: rom = 27;
		13331: rom = 27;
		13332: rom = 27;
		13333: rom = 27;
		13334: rom = 27;
		13335: rom = 27;
		13336: rom = 27;
		13337: rom = 27;
		13338: rom = 27;
		13339: rom = 27;
		13340: rom = 27;
		13341: rom = 27;
		13342: rom = 27;
		13343: rom = 27;
		13344: rom = 27;
		13345: rom = 27;
		13346: rom = 27;
		13347: rom = 27;
		13348: rom = 27;
		13349: rom = 27;
		13350: rom = 27;
		13351: rom = 27;
		13352: rom = 27;
		13353: rom = 27;
		13354: rom = 27;
		13355: rom = 27;
		13356: rom = 27;
		13357: rom = 27;
		13358: rom = 27;
		13359: rom = 27;
		13360: rom = 27;
		13361: rom = 27;
		13362: rom = 27;
		13363: rom = 27;
		13364: rom = 27;
		13365: rom = 27;
		13366: rom = 27;
		13367: rom = 27;
		13368: rom = 27;
		13369: rom = 27;
		13370: rom = 27;
		13371: rom = 27;
		13372: rom = 27;
		13373: rom = 27;
		13374: rom = 27;
		13375: rom = 27;
		13376: rom = 27;
		13377: rom = 27;
		13378: rom = 27;
		13379: rom = 27;
		13380: rom = 27;
		13381: rom = 27;
		13382: rom = 27;
		13383: rom = 27;
		13384: rom = 27;
		13385: rom = 27;
		13386: rom = 27;
		13387: rom = 27;
		13388: rom = 27;
		13389: rom = 27;
		13390: rom = 27;
		13391: rom = 27;
		13392: rom = 20;
		13393: rom = 17;
		13394: rom = 18;
		13395: rom = 18;
		13396: rom = 18;
		13397: rom = 18;
		13398: rom = 18;
		13399: rom = 18;
		13400: rom = 18;
		13401: rom = 18;
		13402: rom = 11;
		13403: rom = 18;
		13404: rom = 18;
		13405: rom = 18;
		13406: rom = 18;
		13407: rom = 18;
		13408: rom = 18;
		13409: rom = 12;
		13410: rom = 18;
		13411: rom = 18;
		13412: rom = 18;
		13413: rom = 18;
		13414: rom = 18;
		13415: rom = 18;
		13416: rom = 18;
		13417: rom = 18;
		13418: rom = 18;
		13419: rom = 18;
		13420: rom = 18;
		13421: rom = 18;
		13422: rom = 18;
		13423: rom = 15;
		13424: rom = 27;
		13425: rom = 27;
		13426: rom = 27;
		13427: rom = 27;
		13428: rom = 27;
		13429: rom = 27;
		13430: rom = 27;
		13431: rom = 27;
		13432: rom = 27;
		13433: rom = 27;
		13434: rom = 27;
		13440: rom = 27;
		13441: rom = 27;
		13442: rom = 27;
		13443: rom = 27;
		13444: rom = 24;
		13445: rom = 24;
		13446: rom = 24;
		13447: rom = 24;
		13448: rom = 24;
		13449: rom = 24;
		13450: rom = 24;
		13451: rom = 24;
		13452: rom = 24;
		13453: rom = 24;
		13454: rom = 24;
		13455: rom = 25;
		13456: rom = 27;
		13457: rom = 27;
		13458: rom = 27;
		13459: rom = 27;
		13460: rom = 27;
		13461: rom = 27;
		13462: rom = 27;
		13463: rom = 27;
		13464: rom = 27;
		13465: rom = 27;
		13466: rom = 27;
		13467: rom = 27;
		13468: rom = 27;
		13469: rom = 27;
		13470: rom = 27;
		13471: rom = 27;
		13472: rom = 27;
		13473: rom = 27;
		13474: rom = 27;
		13475: rom = 27;
		13476: rom = 27;
		13477: rom = 27;
		13478: rom = 27;
		13479: rom = 27;
		13480: rom = 27;
		13481: rom = 27;
		13482: rom = 27;
		13483: rom = 27;
		13484: rom = 27;
		13485: rom = 27;
		13486: rom = 27;
		13487: rom = 27;
		13488: rom = 27;
		13489: rom = 27;
		13490: rom = 27;
		13491: rom = 27;
		13492: rom = 27;
		13493: rom = 27;
		13494: rom = 27;
		13495: rom = 27;
		13496: rom = 27;
		13497: rom = 27;
		13498: rom = 27;
		13499: rom = 27;
		13500: rom = 27;
		13501: rom = 27;
		13502: rom = 27;
		13503: rom = 27;
		13504: rom = 27;
		13505: rom = 27;
		13506: rom = 27;
		13507: rom = 27;
		13508: rom = 27;
		13509: rom = 27;
		13510: rom = 27;
		13511: rom = 27;
		13512: rom = 27;
		13513: rom = 27;
		13514: rom = 27;
		13515: rom = 27;
		13516: rom = 27;
		13517: rom = 27;
		13518: rom = 27;
		13519: rom = 27;
		13520: rom = 19;
		13521: rom = 18;
		13522: rom = 18;
		13523: rom = 18;
		13524: rom = 18;
		13525: rom = 18;
		13526: rom = 18;
		13527: rom = 18;
		13528: rom = 18;
		13529: rom = 18;
		13530: rom = 11;
		13531: rom = 18;
		13532: rom = 18;
		13533: rom = 18;
		13534: rom = 18;
		13535: rom = 18;
		13536: rom = 18;
		13537: rom = 10;
		13538: rom = 18;
		13539: rom = 18;
		13540: rom = 18;
		13541: rom = 18;
		13542: rom = 18;
		13543: rom = 18;
		13544: rom = 18;
		13545: rom = 18;
		13546: rom = 18;
		13547: rom = 18;
		13548: rom = 18;
		13549: rom = 18;
		13550: rom = 18;
		13551: rom = 14;
		13552: rom = 27;
		13553: rom = 27;
		13554: rom = 27;
		13555: rom = 27;
		13556: rom = 27;
		13557: rom = 27;
		13558: rom = 27;
		13559: rom = 27;
		13560: rom = 27;
		13561: rom = 27;
		13562: rom = 27;
		13568: rom = 27;
		13569: rom = 27;
		13570: rom = 27;
		13571: rom = 27;
		13572: rom = 27;
		13573: rom = 27;
		13574: rom = 27;
		13575: rom = 27;
		13576: rom = 27;
		13577: rom = 27;
		13578: rom = 27;
		13579: rom = 27;
		13580: rom = 27;
		13581: rom = 27;
		13582: rom = 27;
		13583: rom = 27;
		13584: rom = 27;
		13585: rom = 27;
		13586: rom = 27;
		13587: rom = 27;
		13588: rom = 27;
		13589: rom = 27;
		13590: rom = 27;
		13591: rom = 27;
		13592: rom = 27;
		13593: rom = 27;
		13594: rom = 27;
		13595: rom = 27;
		13596: rom = 27;
		13597: rom = 27;
		13598: rom = 27;
		13599: rom = 27;
		13600: rom = 27;
		13601: rom = 27;
		13602: rom = 27;
		13603: rom = 27;
		13604: rom = 27;
		13605: rom = 27;
		13606: rom = 27;
		13607: rom = 27;
		13608: rom = 27;
		13609: rom = 27;
		13610: rom = 27;
		13611: rom = 27;
		13612: rom = 27;
		13613: rom = 27;
		13614: rom = 27;
		13615: rom = 27;
		13616: rom = 27;
		13617: rom = 27;
		13618: rom = 27;
		13619: rom = 27;
		13620: rom = 27;
		13621: rom = 27;
		13622: rom = 27;
		13623: rom = 27;
		13624: rom = 27;
		13625: rom = 27;
		13626: rom = 27;
		13627: rom = 27;
		13628: rom = 27;
		13629: rom = 27;
		13630: rom = 27;
		13631: rom = 27;
		13632: rom = 27;
		13633: rom = 27;
		13634: rom = 27;
		13635: rom = 27;
		13636: rom = 27;
		13637: rom = 27;
		13638: rom = 27;
		13639: rom = 27;
		13640: rom = 27;
		13641: rom = 27;
		13642: rom = 27;
		13643: rom = 27;
		13644: rom = 27;
		13645: rom = 27;
		13646: rom = 27;
		13647: rom = 27;
		13648: rom = 17;
		13649: rom = 17;
		13650: rom = 18;
		13651: rom = 18;
		13652: rom = 18;
		13653: rom = 18;
		13654: rom = 18;
		13655: rom = 18;
		13656: rom = 18;
		13657: rom = 18;
		13658: rom = 14;
		13659: rom = 13;
		13660: rom = 18;
		13661: rom = 18;
		13662: rom = 18;
		13663: rom = 18;
		13664: rom = 18;
		13665: rom = 12;
		13666: rom = 18;
		13667: rom = 18;
		13668: rom = 18;
		13669: rom = 18;
		13670: rom = 18;
		13671: rom = 18;
		13672: rom = 18;
		13673: rom = 18;
		13674: rom = 18;
		13675: rom = 18;
		13676: rom = 18;
		13677: rom = 18;
		13678: rom = 18;
		13679: rom = 14;
		13680: rom = 27;
		13681: rom = 27;
		13682: rom = 27;
		13683: rom = 27;
		13684: rom = 27;
		13685: rom = 27;
		13686: rom = 27;
		13687: rom = 27;
		13688: rom = 27;
		13689: rom = 27;
		13690: rom = 27;
		13696: rom = 27;
		13697: rom = 27;
		13698: rom = 27;
		13699: rom = 27;
		13700: rom = 27;
		13701: rom = 27;
		13702: rom = 27;
		13703: rom = 27;
		13704: rom = 27;
		13705: rom = 27;
		13706: rom = 27;
		13707: rom = 27;
		13708: rom = 27;
		13709: rom = 27;
		13710: rom = 27;
		13711: rom = 27;
		13712: rom = 27;
		13713: rom = 27;
		13714: rom = 27;
		13715: rom = 27;
		13716: rom = 27;
		13717: rom = 27;
		13718: rom = 27;
		13719: rom = 27;
		13720: rom = 27;
		13721: rom = 27;
		13722: rom = 27;
		13723: rom = 27;
		13724: rom = 27;
		13725: rom = 27;
		13726: rom = 27;
		13727: rom = 27;
		13728: rom = 27;
		13729: rom = 27;
		13730: rom = 27;
		13731: rom = 27;
		13732: rom = 27;
		13733: rom = 27;
		13734: rom = 27;
		13735: rom = 27;
		13736: rom = 27;
		13737: rom = 27;
		13738: rom = 27;
		13739: rom = 27;
		13740: rom = 27;
		13741: rom = 27;
		13742: rom = 27;
		13743: rom = 27;
		13744: rom = 27;
		13745: rom = 27;
		13746: rom = 27;
		13747: rom = 27;
		13748: rom = 27;
		13749: rom = 27;
		13750: rom = 27;
		13751: rom = 27;
		13752: rom = 27;
		13753: rom = 27;
		13754: rom = 27;
		13755: rom = 27;
		13756: rom = 27;
		13757: rom = 27;
		13758: rom = 27;
		13759: rom = 27;
		13760: rom = 27;
		13761: rom = 27;
		13762: rom = 27;
		13763: rom = 27;
		13764: rom = 27;
		13765: rom = 27;
		13766: rom = 27;
		13767: rom = 27;
		13768: rom = 27;
		13769: rom = 27;
		13770: rom = 27;
		13771: rom = 27;
		13772: rom = 27;
		13773: rom = 27;
		13774: rom = 27;
		13775: rom = 27;
		13776: rom = 17;
		13777: rom = 15;
		13778: rom = 16;
		13779: rom = 18;
		13780: rom = 18;
		13781: rom = 18;
		13782: rom = 18;
		13783: rom = 18;
		13784: rom = 18;
		13785: rom = 18;
		13786: rom = 17;
		13787: rom = 2;
		13788: rom = 17;
		13789: rom = 18;
		13790: rom = 18;
		13791: rom = 18;
		13792: rom = 18;
		13793: rom = 10;
		13794: rom = 18;
		13795: rom = 18;
		13796: rom = 18;
		13797: rom = 18;
		13798: rom = 18;
		13799: rom = 18;
		13800: rom = 18;
		13801: rom = 18;
		13802: rom = 18;
		13803: rom = 18;
		13804: rom = 18;
		13805: rom = 18;
		13806: rom = 18;
		13807: rom = 14;
		13808: rom = 27;
		13809: rom = 27;
		13810: rom = 27;
		13811: rom = 27;
		13812: rom = 27;
		13813: rom = 27;
		13814: rom = 27;
		13815: rom = 27;
		13816: rom = 27;
		13817: rom = 27;
		13818: rom = 27;
		13824: rom = 27;
		13825: rom = 27;
		13826: rom = 27;
		13827: rom = 27;
		13828: rom = 26;
		13829: rom = 26;
		13830: rom = 26;
		13831: rom = 26;
		13832: rom = 26;
		13833: rom = 26;
		13834: rom = 26;
		13835: rom = 26;
		13836: rom = 26;
		13837: rom = 26;
		13838: rom = 26;
		13839: rom = 26;
		13840: rom = 27;
		13841: rom = 27;
		13842: rom = 27;
		13843: rom = 27;
		13844: rom = 27;
		13845: rom = 27;
		13846: rom = 27;
		13847: rom = 27;
		13848: rom = 27;
		13849: rom = 27;
		13850: rom = 27;
		13851: rom = 27;
		13852: rom = 27;
		13853: rom = 27;
		13854: rom = 27;
		13855: rom = 27;
		13856: rom = 27;
		13857: rom = 27;
		13858: rom = 27;
		13859: rom = 27;
		13860: rom = 27;
		13861: rom = 27;
		13862: rom = 27;
		13863: rom = 27;
		13864: rom = 27;
		13865: rom = 27;
		13866: rom = 27;
		13867: rom = 27;
		13868: rom = 27;
		13869: rom = 27;
		13870: rom = 27;
		13871: rom = 27;
		13872: rom = 27;
		13873: rom = 27;
		13874: rom = 27;
		13875: rom = 27;
		13876: rom = 27;
		13877: rom = 27;
		13878: rom = 27;
		13879: rom = 27;
		13880: rom = 27;
		13881: rom = 27;
		13882: rom = 27;
		13883: rom = 27;
		13884: rom = 27;
		13885: rom = 27;
		13886: rom = 27;
		13887: rom = 27;
		13888: rom = 27;
		13889: rom = 27;
		13890: rom = 27;
		13891: rom = 27;
		13892: rom = 27;
		13893: rom = 27;
		13894: rom = 27;
		13895: rom = 27;
		13896: rom = 27;
		13897: rom = 27;
		13898: rom = 27;
		13899: rom = 27;
		13900: rom = 27;
		13901: rom = 27;
		13902: rom = 27;
		13903: rom = 27;
		13904: rom = 17;
		13905: rom = 15;
		13906: rom = 15;
		13907: rom = 18;
		13908: rom = 18;
		13909: rom = 18;
		13910: rom = 18;
		13911: rom = 18;
		13912: rom = 18;
		13913: rom = 18;
		13914: rom = 18;
		13915: rom = 10;
		13916: rom = 12;
		13917: rom = 18;
		13918: rom = 18;
		13919: rom = 18;
		13920: rom = 18;
		13921: rom = 10;
		13922: rom = 17;
		13923: rom = 18;
		13924: rom = 18;
		13925: rom = 18;
		13926: rom = 18;
		13927: rom = 18;
		13928: rom = 18;
		13929: rom = 18;
		13930: rom = 18;
		13931: rom = 18;
		13932: rom = 18;
		13933: rom = 18;
		13934: rom = 18;
		13935: rom = 11;
		13936: rom = 25;
		13937: rom = 27;
		13938: rom = 27;
		13939: rom = 27;
		13940: rom = 27;
		13941: rom = 27;
		13942: rom = 27;
		13943: rom = 27;
		13944: rom = 27;
		13945: rom = 27;
		13946: rom = 27;
		13952: rom = 27;
		13953: rom = 27;
		13954: rom = 27;
		13955: rom = 27;
		13956: rom = 0;
		13957: rom = 0;
		13958: rom = 0;
		13959: rom = 0;
		13960: rom = 0;
		13961: rom = 0;
		13962: rom = 0;
		13963: rom = 0;
		13964: rom = 0;
		13965: rom = 0;
		13966: rom = 0;
		13967: rom = 14;
		13968: rom = 27;
		13969: rom = 27;
		13970: rom = 27;
		13971: rom = 27;
		13972: rom = 27;
		13973: rom = 27;
		13974: rom = 27;
		13975: rom = 27;
		13976: rom = 27;
		13977: rom = 27;
		13978: rom = 27;
		13979: rom = 27;
		13980: rom = 27;
		13981: rom = 27;
		13982: rom = 27;
		13983: rom = 27;
		13984: rom = 27;
		13985: rom = 27;
		13986: rom = 27;
		13987: rom = 27;
		13988: rom = 27;
		13989: rom = 27;
		13990: rom = 27;
		13991: rom = 27;
		13992: rom = 27;
		13993: rom = 27;
		13994: rom = 27;
		13995: rom = 27;
		13996: rom = 27;
		13997: rom = 27;
		13998: rom = 27;
		13999: rom = 27;
		14000: rom = 27;
		14001: rom = 27;
		14002: rom = 27;
		14003: rom = 27;
		14004: rom = 27;
		14005: rom = 27;
		14006: rom = 27;
		14007: rom = 27;
		14008: rom = 27;
		14009: rom = 27;
		14010: rom = 27;
		14011: rom = 27;
		14012: rom = 27;
		14013: rom = 27;
		14014: rom = 27;
		14015: rom = 27;
		14016: rom = 27;
		14017: rom = 27;
		14018: rom = 27;
		14019: rom = 27;
		14020: rom = 27;
		14021: rom = 27;
		14022: rom = 27;
		14023: rom = 27;
		14024: rom = 27;
		14025: rom = 27;
		14026: rom = 27;
		14027: rom = 27;
		14028: rom = 27;
		14029: rom = 27;
		14030: rom = 27;
		14031: rom = 27;
		14032: rom = 19;
		14033: rom = 11;
		14034: rom = 13;
		14035: rom = 18;
		14036: rom = 18;
		14037: rom = 18;
		14038: rom = 18;
		14039: rom = 18;
		14040: rom = 18;
		14041: rom = 18;
		14042: rom = 18;
		14043: rom = 13;
		14044: rom = 18;
		14045: rom = 14;
		14046: rom = 18;
		14047: rom = 18;
		14048: rom = 18;
		14049: rom = 12;
		14050: rom = 17;
		14051: rom = 18;
		14052: rom = 18;
		14053: rom = 18;
		14054: rom = 18;
		14055: rom = 18;
		14056: rom = 18;
		14057: rom = 18;
		14058: rom = 18;
		14059: rom = 18;
		14060: rom = 18;
		14061: rom = 18;
		14062: rom = 18;
		14063: rom = 11;
		14064: rom = 11;
		14065: rom = 23;
		14066: rom = 27;
		14067: rom = 27;
		14068: rom = 27;
		14069: rom = 27;
		14070: rom = 27;
		14071: rom = 27;
		14072: rom = 27;
		14073: rom = 27;
		14074: rom = 27;
		14080: rom = 27;
		14081: rom = 27;
		14082: rom = 27;
		14083: rom = 27;
		14084: rom = 0;
		14085: rom = 0;
		14086: rom = 15;
		14087: rom = 16;
		14088: rom = 16;
		14089: rom = 16;
		14090: rom = 16;
		14091: rom = 16;
		14092: rom = 16;
		14093: rom = 16;
		14094: rom = 16;
		14095: rom = 20;
		14096: rom = 27;
		14097: rom = 27;
		14098: rom = 27;
		14099: rom = 27;
		14100: rom = 27;
		14101: rom = 27;
		14102: rom = 27;
		14103: rom = 27;
		14104: rom = 27;
		14105: rom = 27;
		14106: rom = 27;
		14107: rom = 27;
		14108: rom = 27;
		14109: rom = 27;
		14110: rom = 27;
		14111: rom = 27;
		14112: rom = 27;
		14113: rom = 27;
		14114: rom = 27;
		14115: rom = 27;
		14116: rom = 27;
		14117: rom = 27;
		14118: rom = 27;
		14119: rom = 27;
		14120: rom = 27;
		14121: rom = 27;
		14122: rom = 27;
		14123: rom = 27;
		14124: rom = 27;
		14125: rom = 27;
		14126: rom = 27;
		14127: rom = 27;
		14128: rom = 27;
		14129: rom = 27;
		14130: rom = 27;
		14131: rom = 27;
		14132: rom = 27;
		14133: rom = 27;
		14134: rom = 27;
		14135: rom = 27;
		14136: rom = 27;
		14137: rom = 27;
		14138: rom = 27;
		14139: rom = 27;
		14140: rom = 27;
		14141: rom = 27;
		14142: rom = 27;
		14143: rom = 27;
		14144: rom = 27;
		14145: rom = 27;
		14146: rom = 27;
		14147: rom = 27;
		14148: rom = 27;
		14149: rom = 27;
		14150: rom = 27;
		14151: rom = 27;
		14152: rom = 27;
		14153: rom = 27;
		14154: rom = 27;
		14155: rom = 27;
		14156: rom = 27;
		14157: rom = 27;
		14158: rom = 27;
		14159: rom = 27;
		14160: rom = 27;
		14161: rom = 11;
		14162: rom = 11;
		14163: rom = 18;
		14164: rom = 18;
		14165: rom = 18;
		14166: rom = 18;
		14167: rom = 18;
		14168: rom = 18;
		14169: rom = 18;
		14170: rom = 18;
		14171: rom = 18;
		14172: rom = 11;
		14173: rom = 7;
		14174: rom = 17;
		14175: rom = 18;
		14176: rom = 18;
		14177: rom = 12;
		14178: rom = 17;
		14179: rom = 18;
		14180: rom = 18;
		14181: rom = 18;
		14182: rom = 18;
		14183: rom = 18;
		14184: rom = 18;
		14185: rom = 18;
		14186: rom = 18;
		14187: rom = 18;
		14188: rom = 18;
		14189: rom = 18;
		14190: rom = 18;
		14191: rom = 12;
		14192: rom = 18;
		14193: rom = 12;
		14194: rom = 23;
		14195: rom = 27;
		14196: rom = 27;
		14197: rom = 27;
		14198: rom = 27;
		14199: rom = 27;
		14200: rom = 27;
		14201: rom = 27;
		14202: rom = 27;
		14208: rom = 27;
		14209: rom = 27;
		14210: rom = 27;
		14211: rom = 27;
		14212: rom = 16;
		14213: rom = 0;
		14214: rom = 0;
		14215: rom = 23;
		14216: rom = 27;
		14217: rom = 27;
		14218: rom = 27;
		14219: rom = 27;
		14220: rom = 27;
		14221: rom = 27;
		14222: rom = 27;
		14223: rom = 27;
		14224: rom = 27;
		14225: rom = 27;
		14226: rom = 27;
		14227: rom = 27;
		14228: rom = 27;
		14229: rom = 27;
		14230: rom = 27;
		14231: rom = 27;
		14232: rom = 27;
		14233: rom = 27;
		14234: rom = 27;
		14235: rom = 27;
		14236: rom = 27;
		14237: rom = 27;
		14238: rom = 27;
		14239: rom = 27;
		14240: rom = 27;
		14241: rom = 27;
		14242: rom = 27;
		14243: rom = 27;
		14244: rom = 27;
		14245: rom = 27;
		14246: rom = 27;
		14247: rom = 27;
		14248: rom = 27;
		14249: rom = 27;
		14250: rom = 27;
		14251: rom = 27;
		14252: rom = 27;
		14253: rom = 27;
		14254: rom = 27;
		14255: rom = 27;
		14256: rom = 27;
		14257: rom = 27;
		14258: rom = 27;
		14259: rom = 27;
		14260: rom = 27;
		14261: rom = 27;
		14262: rom = 27;
		14263: rom = 27;
		14264: rom = 27;
		14265: rom = 27;
		14266: rom = 27;
		14267: rom = 27;
		14268: rom = 27;
		14269: rom = 27;
		14270: rom = 27;
		14271: rom = 27;
		14272: rom = 27;
		14273: rom = 27;
		14274: rom = 27;
		14275: rom = 27;
		14276: rom = 27;
		14277: rom = 27;
		14278: rom = 27;
		14279: rom = 27;
		14280: rom = 27;
		14281: rom = 27;
		14282: rom = 27;
		14283: rom = 27;
		14284: rom = 27;
		14285: rom = 27;
		14286: rom = 27;
		14287: rom = 27;
		14288: rom = 27;
		14289: rom = 21;
		14290: rom = 8;
		14291: rom = 18;
		14292: rom = 18;
		14293: rom = 18;
		14294: rom = 18;
		14295: rom = 18;
		14296: rom = 18;
		14297: rom = 18;
		14298: rom = 18;
		14299: rom = 18;
		14300: rom = 18;
		14301: rom = 12;
		14302: rom = 6;
		14303: rom = 17;
		14304: rom = 18;
		14305: rom = 12;
		14306: rom = 17;
		14307: rom = 18;
		14308: rom = 18;
		14309: rom = 18;
		14310: rom = 18;
		14311: rom = 18;
		14312: rom = 18;
		14313: rom = 18;
		14314: rom = 18;
		14315: rom = 18;
		14316: rom = 18;
		14317: rom = 18;
		14318: rom = 18;
		14319: rom = 11;
		14320: rom = 18;
		14321: rom = 18;
		14322: rom = 12;
		14323: rom = 26;
		14324: rom = 27;
		14325: rom = 27;
		14326: rom = 27;
		14327: rom = 27;
		14328: rom = 27;
		14329: rom = 27;
		14330: rom = 27;
		14336: rom = 27;
		14337: rom = 27;
		14338: rom = 27;
		14339: rom = 27;
		14340: rom = 27;
		14341: rom = 23;
		14342: rom = 0;
		14343: rom = 0;
		14344: rom = 15;
		14345: rom = 25;
		14346: rom = 27;
		14347: rom = 27;
		14348: rom = 27;
		14349: rom = 27;
		14350: rom = 27;
		14351: rom = 27;
		14352: rom = 27;
		14353: rom = 27;
		14354: rom = 27;
		14355: rom = 27;
		14356: rom = 27;
		14357: rom = 27;
		14358: rom = 27;
		14359: rom = 27;
		14360: rom = 27;
		14361: rom = 27;
		14362: rom = 27;
		14363: rom = 27;
		14364: rom = 27;
		14365: rom = 27;
		14366: rom = 27;
		14367: rom = 27;
		14368: rom = 27;
		14369: rom = 27;
		14370: rom = 27;
		14371: rom = 27;
		14372: rom = 27;
		14373: rom = 27;
		14374: rom = 27;
		14375: rom = 27;
		14376: rom = 27;
		14377: rom = 27;
		14378: rom = 27;
		14379: rom = 27;
		14380: rom = 27;
		14381: rom = 27;
		14382: rom = 27;
		14383: rom = 27;
		14384: rom = 27;
		14385: rom = 27;
		14386: rom = 27;
		14387: rom = 27;
		14388: rom = 27;
		14389: rom = 27;
		14390: rom = 27;
		14391: rom = 27;
		14392: rom = 27;
		14393: rom = 27;
		14394: rom = 27;
		14395: rom = 27;
		14396: rom = 27;
		14397: rom = 27;
		14398: rom = 27;
		14399: rom = 27;
		14400: rom = 27;
		14401: rom = 27;
		14402: rom = 27;
		14403: rom = 27;
		14404: rom = 27;
		14405: rom = 27;
		14406: rom = 27;
		14407: rom = 27;
		14408: rom = 27;
		14409: rom = 27;
		14410: rom = 27;
		14411: rom = 27;
		14412: rom = 27;
		14413: rom = 27;
		14414: rom = 27;
		14415: rom = 27;
		14416: rom = 27;
		14417: rom = 27;
		14418: rom = 16;
		14419: rom = 18;
		14420: rom = 18;
		14421: rom = 18;
		14422: rom = 18;
		14423: rom = 18;
		14424: rom = 18;
		14425: rom = 18;
		14426: rom = 18;
		14427: rom = 18;
		14428: rom = 18;
		14429: rom = 18;
		14430: rom = 10;
		14431: rom = 8;
		14432: rom = 15;
		14433: rom = 10;
		14434: rom = 17;
		14435: rom = 18;
		14436: rom = 18;
		14437: rom = 18;
		14438: rom = 18;
		14439: rom = 18;
		14440: rom = 18;
		14441: rom = 18;
		14442: rom = 18;
		14443: rom = 18;
		14444: rom = 18;
		14445: rom = 18;
		14446: rom = 18;
		14447: rom = 7;
		14448: rom = 17;
		14449: rom = 18;
		14450: rom = 17;
		14451: rom = 18;
		14452: rom = 27;
		14453: rom = 27;
		14454: rom = 27;
		14455: rom = 27;
		14456: rom = 27;
		14457: rom = 27;
		14458: rom = 27;
		14464: rom = 27;
		14465: rom = 27;
		14466: rom = 27;
		14467: rom = 27;
		14468: rom = 27;
		14469: rom = 27;
		14470: rom = 27;
		14471: rom = 19;
		14472: rom = 0;
		14473: rom = 0;
		14474: rom = 20;
		14475: rom = 27;
		14476: rom = 27;
		14477: rom = 27;
		14478: rom = 27;
		14479: rom = 27;
		14480: rom = 27;
		14481: rom = 27;
		14482: rom = 27;
		14483: rom = 27;
		14484: rom = 27;
		14485: rom = 27;
		14486: rom = 27;
		14487: rom = 27;
		14488: rom = 27;
		14489: rom = 27;
		14490: rom = 27;
		14491: rom = 27;
		14492: rom = 27;
		14493: rom = 27;
		14494: rom = 27;
		14495: rom = 27;
		14496: rom = 27;
		14497: rom = 27;
		14498: rom = 27;
		14499: rom = 27;
		14500: rom = 27;
		14501: rom = 27;
		14502: rom = 27;
		14503: rom = 27;
		14504: rom = 27;
		14505: rom = 27;
		14506: rom = 27;
		14507: rom = 27;
		14508: rom = 27;
		14509: rom = 27;
		14510: rom = 27;
		14511: rom = 27;
		14512: rom = 27;
		14513: rom = 27;
		14514: rom = 27;
		14515: rom = 27;
		14516: rom = 27;
		14517: rom = 27;
		14518: rom = 27;
		14519: rom = 27;
		14520: rom = 27;
		14521: rom = 27;
		14522: rom = 27;
		14523: rom = 27;
		14524: rom = 27;
		14525: rom = 27;
		14526: rom = 27;
		14527: rom = 27;
		14528: rom = 27;
		14529: rom = 27;
		14530: rom = 27;
		14531: rom = 27;
		14532: rom = 27;
		14533: rom = 27;
		14534: rom = 27;
		14535: rom = 27;
		14536: rom = 27;
		14537: rom = 27;
		14538: rom = 27;
		14539: rom = 27;
		14540: rom = 27;
		14541: rom = 27;
		14542: rom = 27;
		14543: rom = 27;
		14544: rom = 27;
		14545: rom = 27;
		14546: rom = 21;
		14547: rom = 16;
		14548: rom = 18;
		14549: rom = 18;
		14550: rom = 18;
		14551: rom = 18;
		14552: rom = 18;
		14553: rom = 18;
		14554: rom = 18;
		14555: rom = 18;
		14556: rom = 18;
		14557: rom = 18;
		14558: rom = 15;
		14559: rom = 22;
		14560: rom = 19;
		14561: rom = 8;
		14562: rom = 18;
		14563: rom = 18;
		14564: rom = 18;
		14565: rom = 18;
		14566: rom = 18;
		14567: rom = 18;
		14568: rom = 18;
		14569: rom = 18;
		14570: rom = 18;
		14571: rom = 18;
		14572: rom = 18;
		14573: rom = 18;
		14574: rom = 18;
		14575: rom = 6;
		14576: rom = 12;
		14577: rom = 18;
		14578: rom = 18;
		14579: rom = 12;
		14580: rom = 27;
		14581: rom = 27;
		14582: rom = 27;
		14583: rom = 27;
		14584: rom = 27;
		14585: rom = 27;
		14586: rom = 27;
		14592: rom = 27;
		14593: rom = 27;
		14594: rom = 27;
		14595: rom = 27;
		14596: rom = 27;
		14597: rom = 27;
		14598: rom = 27;
		14599: rom = 27;
		14600: rom = 25;
		14601: rom = 15;
		14602: rom = 0;
		14603: rom = 0;
		14604: rom = 23;
		14605: rom = 27;
		14606: rom = 27;
		14607: rom = 27;
		14608: rom = 27;
		14609: rom = 27;
		14610: rom = 27;
		14611: rom = 27;
		14612: rom = 27;
		14613: rom = 27;
		14614: rom = 27;
		14615: rom = 27;
		14616: rom = 27;
		14617: rom = 27;
		14618: rom = 27;
		14619: rom = 27;
		14620: rom = 27;
		14621: rom = 27;
		14622: rom = 27;
		14623: rom = 27;
		14624: rom = 27;
		14625: rom = 27;
		14626: rom = 27;
		14627: rom = 27;
		14628: rom = 27;
		14629: rom = 27;
		14630: rom = 27;
		14631: rom = 27;
		14632: rom = 27;
		14633: rom = 27;
		14634: rom = 27;
		14635: rom = 27;
		14636: rom = 27;
		14637: rom = 27;
		14638: rom = 27;
		14639: rom = 27;
		14640: rom = 27;
		14641: rom = 27;
		14642: rom = 27;
		14643: rom = 27;
		14644: rom = 27;
		14645: rom = 27;
		14646: rom = 27;
		14647: rom = 27;
		14648: rom = 27;
		14649: rom = 27;
		14650: rom = 27;
		14651: rom = 27;
		14652: rom = 27;
		14653: rom = 27;
		14654: rom = 27;
		14655: rom = 27;
		14656: rom = 27;
		14657: rom = 27;
		14658: rom = 27;
		14659: rom = 27;
		14660: rom = 27;
		14661: rom = 27;
		14662: rom = 27;
		14663: rom = 27;
		14664: rom = 27;
		14665: rom = 27;
		14666: rom = 27;
		14667: rom = 27;
		14668: rom = 27;
		14669: rom = 27;
		14670: rom = 27;
		14671: rom = 27;
		14672: rom = 27;
		14673: rom = 27;
		14674: rom = 24;
		14675: rom = 14;
		14676: rom = 18;
		14677: rom = 18;
		14678: rom = 18;
		14679: rom = 18;
		14680: rom = 18;
		14681: rom = 18;
		14682: rom = 18;
		14683: rom = 18;
		14684: rom = 10;
		14685: rom = 11;
		14686: rom = 9;
		14687: rom = 24;
		14688: rom = 27;
		14689: rom = 16;
		14690: rom = 18;
		14691: rom = 18;
		14692: rom = 18;
		14693: rom = 18;
		14694: rom = 18;
		14695: rom = 18;
		14696: rom = 18;
		14697: rom = 18;
		14698: rom = 18;
		14699: rom = 18;
		14700: rom = 18;
		14701: rom = 18;
		14702: rom = 18;
		14703: rom = 4;
		14704: rom = 10;
		14705: rom = 18;
		14706: rom = 18;
		14707: rom = 15;
		14708: rom = 23;
		14709: rom = 27;
		14710: rom = 27;
		14711: rom = 27;
		14712: rom = 27;
		14713: rom = 27;
		14714: rom = 27;
		14720: rom = 27;
		14721: rom = 27;
		14722: rom = 27;
		14723: rom = 27;
		14724: rom = 27;
		14725: rom = 27;
		14726: rom = 27;
		14727: rom = 27;
		14728: rom = 27;
		14729: rom = 27;
		14730: rom = 22;
		14731: rom = 0;
		14732: rom = 0;
		14733: rom = 16;
		14734: rom = 26;
		14735: rom = 27;
		14736: rom = 27;
		14737: rom = 27;
		14738: rom = 27;
		14739: rom = 27;
		14740: rom = 27;
		14741: rom = 27;
		14742: rom = 27;
		14743: rom = 27;
		14744: rom = 27;
		14745: rom = 27;
		14746: rom = 27;
		14747: rom = 27;
		14748: rom = 27;
		14749: rom = 27;
		14750: rom = 27;
		14751: rom = 27;
		14752: rom = 27;
		14753: rom = 27;
		14754: rom = 27;
		14755: rom = 27;
		14756: rom = 27;
		14757: rom = 27;
		14758: rom = 27;
		14759: rom = 27;
		14760: rom = 27;
		14761: rom = 27;
		14762: rom = 27;
		14763: rom = 27;
		14764: rom = 27;
		14765: rom = 27;
		14766: rom = 27;
		14767: rom = 27;
		14768: rom = 27;
		14769: rom = 27;
		14770: rom = 27;
		14771: rom = 27;
		14772: rom = 27;
		14773: rom = 27;
		14774: rom = 27;
		14775: rom = 27;
		14776: rom = 27;
		14777: rom = 27;
		14778: rom = 27;
		14779: rom = 27;
		14780: rom = 27;
		14781: rom = 27;
		14782: rom = 27;
		14783: rom = 27;
		14784: rom = 27;
		14785: rom = 27;
		14786: rom = 27;
		14787: rom = 27;
		14788: rom = 27;
		14789: rom = 27;
		14790: rom = 27;
		14791: rom = 27;
		14792: rom = 27;
		14793: rom = 27;
		14794: rom = 27;
		14795: rom = 27;
		14796: rom = 27;
		14797: rom = 27;
		14798: rom = 27;
		14799: rom = 27;
		14800: rom = 27;
		14801: rom = 27;
		14802: rom = 27;
		14803: rom = 12;
		14804: rom = 18;
		14805: rom = 18;
		14806: rom = 18;
		14807: rom = 18;
		14808: rom = 18;
		14809: rom = 14;
		14810: rom = 16;
		14811: rom = 17;
		14812: rom = 11;
		14813: rom = 19;
		14814: rom = 16;
		14815: rom = 13;
		14816: rom = 23;
		14817: rom = 12;
		14818: rom = 18;
		14819: rom = 18;
		14820: rom = 18;
		14821: rom = 18;
		14822: rom = 18;
		14823: rom = 18;
		14824: rom = 18;
		14825: rom = 18;
		14826: rom = 18;
		14827: rom = 18;
		14828: rom = 18;
		14829: rom = 18;
		14830: rom = 18;
		14831: rom = 5;
		14832: rom = 7;
		14833: rom = 17;
		14834: rom = 18;
		14835: rom = 17;
		14836: rom = 19;
		14837: rom = 27;
		14838: rom = 27;
		14839: rom = 27;
		14840: rom = 27;
		14841: rom = 27;
		14842: rom = 27;
		14848: rom = 27;
		14849: rom = 27;
		14850: rom = 27;
		14851: rom = 27;
		14852: rom = 27;
		14853: rom = 27;
		14854: rom = 27;
		14855: rom = 27;
		14856: rom = 27;
		14857: rom = 27;
		14858: rom = 27;
		14859: rom = 27;
		14860: rom = 19;
		14861: rom = 0;
		14862: rom = 0;
		14863: rom = 22;
		14864: rom = 27;
		14865: rom = 27;
		14866: rom = 27;
		14867: rom = 27;
		14868: rom = 27;
		14869: rom = 27;
		14870: rom = 27;
		14871: rom = 27;
		14872: rom = 27;
		14873: rom = 27;
		14874: rom = 27;
		14875: rom = 27;
		14876: rom = 27;
		14877: rom = 27;
		14878: rom = 27;
		14879: rom = 27;
		14880: rom = 27;
		14881: rom = 27;
		14882: rom = 27;
		14883: rom = 27;
		14884: rom = 27;
		14885: rom = 27;
		14886: rom = 27;
		14887: rom = 27;
		14888: rom = 27;
		14889: rom = 27;
		14890: rom = 27;
		14891: rom = 27;
		14892: rom = 27;
		14893: rom = 27;
		14894: rom = 27;
		14895: rom = 27;
		14896: rom = 27;
		14897: rom = 27;
		14898: rom = 27;
		14899: rom = 27;
		14900: rom = 27;
		14901: rom = 27;
		14902: rom = 27;
		14903: rom = 27;
		14904: rom = 27;
		14905: rom = 27;
		14906: rom = 27;
		14907: rom = 27;
		14908: rom = 27;
		14909: rom = 27;
		14910: rom = 27;
		14911: rom = 27;
		14912: rom = 27;
		14913: rom = 27;
		14914: rom = 27;
		14915: rom = 27;
		14916: rom = 27;
		14917: rom = 27;
		14918: rom = 27;
		14919: rom = 27;
		14920: rom = 27;
		14921: rom = 27;
		14922: rom = 27;
		14923: rom = 27;
		14924: rom = 27;
		14925: rom = 27;
		14926: rom = 27;
		14927: rom = 27;
		14928: rom = 27;
		14929: rom = 27;
		14930: rom = 27;
		14931: rom = 15;
		14932: rom = 18;
		14933: rom = 18;
		14934: rom = 18;
		14935: rom = 18;
		14936: rom = 18;
		14937: rom = 18;
		14938: rom = 11;
		14939: rom = 15;
		14940: rom = 16;
		14941: rom = 11;
		14942: rom = 5;
		14943: rom = 15;
		14944: rom = 22;
		14945: rom = 11;
		14946: rom = 18;
		14947: rom = 18;
		14948: rom = 18;
		14949: rom = 18;
		14950: rom = 18;
		14951: rom = 18;
		14952: rom = 18;
		14953: rom = 18;
		14954: rom = 18;
		14955: rom = 18;
		14956: rom = 18;
		14957: rom = 18;
		14958: rom = 17;
		14959: rom = 12;
		14960: rom = 14;
		14961: rom = 18;
		14962: rom = 18;
		14963: rom = 18;
		14964: rom = 16;
		14965: rom = 27;
		14966: rom = 27;
		14967: rom = 27;
		14968: rom = 27;
		14969: rom = 27;
		14970: rom = 27;
		14976: rom = 27;
		14977: rom = 27;
		14978: rom = 27;
		14979: rom = 27;
		14980: rom = 17;
		14981: rom = 17;
		14982: rom = 17;
		14983: rom = 17;
		14984: rom = 17;
		14985: rom = 17;
		14986: rom = 17;
		14987: rom = 17;
		14988: rom = 17;
		14989: rom = 11;
		14990: rom = 0;
		14991: rom = 14;
		14992: rom = 27;
		14993: rom = 27;
		14994: rom = 27;
		14995: rom = 27;
		14996: rom = 27;
		14997: rom = 27;
		14998: rom = 27;
		14999: rom = 27;
		15000: rom = 27;
		15001: rom = 27;
		15002: rom = 27;
		15003: rom = 27;
		15004: rom = 27;
		15005: rom = 27;
		15006: rom = 27;
		15007: rom = 27;
		15008: rom = 27;
		15009: rom = 27;
		15010: rom = 27;
		15011: rom = 27;
		15012: rom = 27;
		15013: rom = 27;
		15014: rom = 27;
		15015: rom = 27;
		15016: rom = 27;
		15017: rom = 27;
		15018: rom = 27;
		15019: rom = 27;
		15020: rom = 27;
		15021: rom = 27;
		15022: rom = 27;
		15023: rom = 27;
		15024: rom = 27;
		15025: rom = 27;
		15026: rom = 27;
		15027: rom = 27;
		15028: rom = 27;
		15029: rom = 27;
		15030: rom = 27;
		15031: rom = 27;
		15032: rom = 27;
		15033: rom = 27;
		15034: rom = 27;
		15035: rom = 27;
		15036: rom = 27;
		15037: rom = 27;
		15038: rom = 27;
		15039: rom = 27;
		15040: rom = 27;
		15041: rom = 27;
		15042: rom = 27;
		15043: rom = 27;
		15044: rom = 27;
		15045: rom = 27;
		15046: rom = 27;
		15047: rom = 27;
		15048: rom = 27;
		15049: rom = 27;
		15050: rom = 27;
		15051: rom = 27;
		15052: rom = 27;
		15053: rom = 27;
		15054: rom = 27;
		15055: rom = 27;
		15056: rom = 27;
		15057: rom = 27;
		15058: rom = 27;
		15059: rom = 20;
		15060: rom = 17;
		15061: rom = 18;
		15062: rom = 18;
		15063: rom = 18;
		15064: rom = 18;
		15065: rom = 18;
		15066: rom = 18;
		15067: rom = 14;
		15068: rom = 9;
		15069: rom = 12;
		15070: rom = 17;
		15071: rom = 27;
		15072: rom = 25;
		15073: rom = 13;
		15074: rom = 18;
		15075: rom = 18;
		15076: rom = 18;
		15077: rom = 18;
		15078: rom = 18;
		15079: rom = 18;
		15080: rom = 18;
		15081: rom = 18;
		15082: rom = 18;
		15083: rom = 18;
		15084: rom = 18;
		15085: rom = 18;
		15086: rom = 16;
		15087: rom = 14;
		15088: rom = 18;
		15089: rom = 18;
		15090: rom = 18;
		15091: rom = 18;
		15092: rom = 11;
		15093: rom = 27;
		15094: rom = 27;
		15095: rom = 27;
		15096: rom = 27;
		15097: rom = 27;
		15098: rom = 27;
		15104: rom = 27;
		15105: rom = 27;
		15106: rom = 27;
		15107: rom = 27;
		15108: rom = 0;
		15109: rom = 0;
		15110: rom = 0;
		15111: rom = 0;
		15112: rom = 0;
		15113: rom = 0;
		15114: rom = 0;
		15115: rom = 0;
		15116: rom = 0;
		15117: rom = 0;
		15118: rom = 0;
		15119: rom = 14;
		15120: rom = 27;
		15121: rom = 27;
		15122: rom = 27;
		15123: rom = 27;
		15124: rom = 27;
		15125: rom = 27;
		15126: rom = 27;
		15127: rom = 27;
		15128: rom = 27;
		15129: rom = 27;
		15130: rom = 27;
		15131: rom = 27;
		15132: rom = 27;
		15133: rom = 27;
		15134: rom = 27;
		15135: rom = 27;
		15136: rom = 27;
		15137: rom = 27;
		15138: rom = 27;
		15139: rom = 27;
		15140: rom = 27;
		15141: rom = 27;
		15142: rom = 27;
		15143: rom = 27;
		15144: rom = 27;
		15145: rom = 27;
		15146: rom = 27;
		15147: rom = 27;
		15148: rom = 27;
		15149: rom = 27;
		15150: rom = 27;
		15151: rom = 27;
		15152: rom = 27;
		15153: rom = 27;
		15154: rom = 27;
		15155: rom = 27;
		15156: rom = 27;
		15157: rom = 27;
		15158: rom = 27;
		15159: rom = 27;
		15160: rom = 27;
		15161: rom = 27;
		15162: rom = 27;
		15163: rom = 27;
		15164: rom = 27;
		15165: rom = 27;
		15166: rom = 27;
		15167: rom = 27;
		15168: rom = 27;
		15169: rom = 27;
		15170: rom = 27;
		15171: rom = 27;
		15172: rom = 27;
		15173: rom = 27;
		15174: rom = 27;
		15175: rom = 27;
		15176: rom = 27;
		15177: rom = 27;
		15178: rom = 27;
		15179: rom = 27;
		15180: rom = 27;
		15181: rom = 27;
		15182: rom = 27;
		15183: rom = 27;
		15184: rom = 27;
		15185: rom = 27;
		15186: rom = 27;
		15187: rom = 25;
		15188: rom = 13;
		15189: rom = 18;
		15190: rom = 18;
		15191: rom = 16;
		15192: rom = 18;
		15193: rom = 18;
		15194: rom = 16;
		15195: rom = 18;
		15196: rom = 17;
		15197: rom = 16;
		15198: rom = 27;
		15199: rom = 27;
		15200: rom = 22;
		15201: rom = 15;
		15202: rom = 18;
		15203: rom = 18;
		15204: rom = 18;
		15205: rom = 18;
		15206: rom = 18;
		15207: rom = 18;
		15208: rom = 18;
		15209: rom = 18;
		15210: rom = 18;
		15211: rom = 18;
		15212: rom = 18;
		15213: rom = 18;
		15214: rom = 15;
		15215: rom = 15;
		15216: rom = 18;
		15217: rom = 18;
		15218: rom = 18;
		15219: rom = 18;
		15220: rom = 12;
		15221: rom = 25;
		15222: rom = 27;
		15223: rom = 27;
		15224: rom = 27;
		15225: rom = 27;
		15226: rom = 27;
		15232: rom = 27;
		15233: rom = 27;
		15234: rom = 27;
		15235: rom = 27;
		15236: rom = 26;
		15237: rom = 26;
		15238: rom = 26;
		15239: rom = 26;
		15240: rom = 26;
		15241: rom = 26;
		15242: rom = 26;
		15243: rom = 26;
		15244: rom = 26;
		15245: rom = 26;
		15246: rom = 26;
		15247: rom = 26;
		15248: rom = 27;
		15249: rom = 27;
		15250: rom = 27;
		15251: rom = 27;
		15252: rom = 27;
		15253: rom = 27;
		15254: rom = 27;
		15255: rom = 27;
		15256: rom = 27;
		15257: rom = 27;
		15258: rom = 27;
		15259: rom = 27;
		15260: rom = 27;
		15261: rom = 27;
		15262: rom = 27;
		15263: rom = 27;
		15264: rom = 27;
		15265: rom = 27;
		15266: rom = 27;
		15267: rom = 27;
		15268: rom = 27;
		15269: rom = 27;
		15270: rom = 27;
		15271: rom = 27;
		15272: rom = 27;
		15273: rom = 27;
		15274: rom = 27;
		15275: rom = 27;
		15276: rom = 27;
		15277: rom = 27;
		15278: rom = 27;
		15279: rom = 27;
		15280: rom = 27;
		15281: rom = 27;
		15282: rom = 27;
		15283: rom = 27;
		15284: rom = 27;
		15285: rom = 27;
		15286: rom = 27;
		15287: rom = 27;
		15288: rom = 27;
		15289: rom = 27;
		15290: rom = 27;
		15291: rom = 27;
		15292: rom = 27;
		15293: rom = 27;
		15294: rom = 27;
		15295: rom = 27;
		15296: rom = 27;
		15297: rom = 27;
		15298: rom = 27;
		15299: rom = 27;
		15300: rom = 27;
		15301: rom = 27;
		15302: rom = 27;
		15303: rom = 27;
		15304: rom = 27;
		15305: rom = 27;
		15306: rom = 27;
		15307: rom = 27;
		15308: rom = 27;
		15309: rom = 27;
		15310: rom = 27;
		15311: rom = 27;
		15312: rom = 27;
		15313: rom = 27;
		15314: rom = 27;
		15315: rom = 27;
		15316: rom = 12;
		15317: rom = 18;
		15318: rom = 18;
		15319: rom = 12;
		15320: rom = 18;
		15321: rom = 14;
		15322: rom = 13;
		15323: rom = 11;
		15324: rom = 13;
		15325: rom = 17;
		15326: rom = 27;
		15327: rom = 27;
		15328: rom = 19;
		15329: rom = 17;
		15330: rom = 18;
		15331: rom = 18;
		15332: rom = 18;
		15333: rom = 18;
		15334: rom = 18;
		15335: rom = 18;
		15336: rom = 18;
		15337: rom = 18;
		15338: rom = 18;
		15339: rom = 18;
		15340: rom = 18;
		15341: rom = 18;
		15342: rom = 13;
		15343: rom = 16;
		15344: rom = 18;
		15345: rom = 18;
		15346: rom = 18;
		15347: rom = 18;
		15348: rom = 15;
		15349: rom = 23;
		15350: rom = 27;
		15351: rom = 27;
		15352: rom = 27;
		15353: rom = 27;
		15354: rom = 27;
		15360: rom = 27;
		15361: rom = 27;
		15362: rom = 27;
		15363: rom = 27;
		15364: rom = 27;
		15365: rom = 27;
		15366: rom = 27;
		15367: rom = 27;
		15368: rom = 27;
		15369: rom = 27;
		15370: rom = 27;
		15371: rom = 27;
		15372: rom = 27;
		15373: rom = 27;
		15374: rom = 27;
		15375: rom = 27;
		15376: rom = 27;
		15377: rom = 27;
		15378: rom = 27;
		15379: rom = 27;
		15380: rom = 27;
		15381: rom = 27;
		15382: rom = 27;
		15383: rom = 27;
		15384: rom = 27;
		15385: rom = 27;
		15386: rom = 27;
		15387: rom = 27;
		15388: rom = 27;
		15389: rom = 27;
		15390: rom = 27;
		15391: rom = 27;
		15392: rom = 27;
		15393: rom = 27;
		15394: rom = 27;
		15395: rom = 27;
		15396: rom = 27;
		15397: rom = 27;
		15398: rom = 27;
		15399: rom = 27;
		15400: rom = 27;
		15401: rom = 27;
		15402: rom = 27;
		15403: rom = 27;
		15404: rom = 27;
		15405: rom = 27;
		15406: rom = 27;
		15407: rom = 27;
		15408: rom = 27;
		15409: rom = 27;
		15410: rom = 27;
		15411: rom = 27;
		15412: rom = 27;
		15413: rom = 27;
		15414: rom = 27;
		15415: rom = 27;
		15416: rom = 27;
		15417: rom = 27;
		15418: rom = 27;
		15419: rom = 27;
		15420: rom = 27;
		15421: rom = 27;
		15422: rom = 27;
		15423: rom = 27;
		15424: rom = 27;
		15425: rom = 27;
		15426: rom = 27;
		15427: rom = 27;
		15428: rom = 27;
		15429: rom = 27;
		15430: rom = 27;
		15431: rom = 27;
		15432: rom = 27;
		15433: rom = 27;
		15434: rom = 27;
		15435: rom = 27;
		15436: rom = 27;
		15437: rom = 27;
		15438: rom = 27;
		15439: rom = 27;
		15440: rom = 27;
		15441: rom = 27;
		15442: rom = 27;
		15443: rom = 27;
		15444: rom = 21;
		15445: rom = 15;
		15446: rom = 18;
		15447: rom = 15;
		15448: rom = 14;
		15449: rom = 17;
		15450: rom = 10;
		15451: rom = 16;
		15452: rom = 14;
		15453: rom = 11;
		15454: rom = 21;
		15455: rom = 27;
		15456: rom = 15;
		15457: rom = 18;
		15458: rom = 18;
		15459: rom = 18;
		15460: rom = 18;
		15461: rom = 18;
		15462: rom = 18;
		15463: rom = 18;
		15464: rom = 18;
		15465: rom = 18;
		15466: rom = 18;
		15467: rom = 18;
		15468: rom = 18;
		15469: rom = 18;
		15470: rom = 12;
		15471: rom = 18;
		15472: rom = 18;
		15473: rom = 18;
		15474: rom = 18;
		15475: rom = 18;
		15476: rom = 18;
		15477: rom = 17;
		15478: rom = 27;
		15479: rom = 27;
		15480: rom = 27;
		15481: rom = 27;
		15482: rom = 27;
		15488: rom = 27;
		15489: rom = 27;
		15490: rom = 27;
		15491: rom = 27;
		15492: rom = 27;
		15493: rom = 27;
		15494: rom = 27;
		15495: rom = 27;
		15496: rom = 27;
		15497: rom = 27;
		15498: rom = 27;
		15499: rom = 27;
		15500: rom = 27;
		15501: rom = 27;
		15502: rom = 27;
		15503: rom = 27;
		15504: rom = 27;
		15505: rom = 27;
		15506: rom = 27;
		15507: rom = 27;
		15508: rom = 27;
		15509: rom = 27;
		15510: rom = 27;
		15511: rom = 27;
		15512: rom = 27;
		15513: rom = 27;
		15514: rom = 27;
		15515: rom = 27;
		15516: rom = 27;
		15517: rom = 27;
		15518: rom = 27;
		15519: rom = 27;
		15520: rom = 27;
		15521: rom = 27;
		15522: rom = 27;
		15523: rom = 27;
		15524: rom = 27;
		15525: rom = 27;
		15526: rom = 27;
		15527: rom = 27;
		15528: rom = 27;
		15529: rom = 27;
		15530: rom = 27;
		15531: rom = 27;
		15532: rom = 27;
		15533: rom = 27;
		15534: rom = 27;
		15535: rom = 27;
		15536: rom = 27;
		15537: rom = 27;
		15538: rom = 27;
		15539: rom = 27;
		15540: rom = 27;
		15541: rom = 27;
		15542: rom = 27;
		15543: rom = 27;
		15544: rom = 27;
		15545: rom = 27;
		15546: rom = 27;
		15547: rom = 27;
		15548: rom = 27;
		15549: rom = 27;
		15550: rom = 27;
		15551: rom = 27;
		15552: rom = 27;
		15553: rom = 27;
		15554: rom = 27;
		15555: rom = 27;
		15556: rom = 27;
		15557: rom = 27;
		15558: rom = 27;
		15559: rom = 27;
		15560: rom = 27;
		15561: rom = 27;
		15562: rom = 27;
		15563: rom = 27;
		15564: rom = 27;
		15565: rom = 27;
		15566: rom = 27;
		15567: rom = 27;
		15568: rom = 27;
		15569: rom = 27;
		15570: rom = 27;
		15571: rom = 27;
		15572: rom = 27;
		15573: rom = 15;
		15574: rom = 16;
		15575: rom = 12;
		15576: rom = 7;
		15577: rom = 14;
		15578: rom = 16;
		15579: rom = 7;
		15580: rom = 13;
		15581: rom = 17;
		15582: rom = 19;
		15583: rom = 26;
		15584: rom = 11;
		15585: rom = 18;
		15586: rom = 18;
		15587: rom = 18;
		15588: rom = 18;
		15589: rom = 18;
		15590: rom = 18;
		15591: rom = 18;
		15592: rom = 18;
		15593: rom = 18;
		15594: rom = 18;
		15595: rom = 18;
		15596: rom = 18;
		15597: rom = 18;
		15598: rom = 11;
		15599: rom = 18;
		15600: rom = 18;
		15601: rom = 18;
		15602: rom = 18;
		15603: rom = 18;
		15604: rom = 18;
		15605: rom = 12;
		15606: rom = 27;
		15607: rom = 27;
		15608: rom = 27;
		15609: rom = 27;
		15610: rom = 27;
		15616: rom = 27;
		15617: rom = 27;
		15618: rom = 27;
		15619: rom = 27;
		15620: rom = 27;
		15621: rom = 27;
		15622: rom = 27;
		15623: rom = 27;
		15624: rom = 27;
		15625: rom = 27;
		15626: rom = 27;
		15627: rom = 27;
		15628: rom = 27;
		15629: rom = 27;
		15630: rom = 27;
		15631: rom = 27;
		15632: rom = 27;
		15633: rom = 27;
		15634: rom = 27;
		15635: rom = 27;
		15636: rom = 27;
		15637: rom = 27;
		15638: rom = 27;
		15639: rom = 27;
		15640: rom = 27;
		15641: rom = 27;
		15642: rom = 27;
		15643: rom = 27;
		15644: rom = 27;
		15645: rom = 27;
		15646: rom = 27;
		15647: rom = 27;
		15648: rom = 27;
		15649: rom = 27;
		15650: rom = 27;
		15651: rom = 27;
		15652: rom = 27;
		15653: rom = 27;
		15654: rom = 27;
		15655: rom = 27;
		15656: rom = 27;
		15657: rom = 27;
		15658: rom = 27;
		15659: rom = 27;
		15660: rom = 27;
		15661: rom = 27;
		15662: rom = 27;
		15663: rom = 27;
		15664: rom = 27;
		15665: rom = 27;
		15666: rom = 27;
		15667: rom = 27;
		15668: rom = 27;
		15669: rom = 27;
		15670: rom = 27;
		15671: rom = 27;
		15672: rom = 27;
		15673: rom = 27;
		15674: rom = 27;
		15675: rom = 27;
		15676: rom = 27;
		15677: rom = 27;
		15678: rom = 27;
		15679: rom = 27;
		15680: rom = 27;
		15681: rom = 27;
		15682: rom = 27;
		15683: rom = 27;
		15684: rom = 27;
		15685: rom = 27;
		15686: rom = 27;
		15687: rom = 27;
		15688: rom = 27;
		15689: rom = 27;
		15690: rom = 27;
		15691: rom = 27;
		15692: rom = 27;
		15693: rom = 27;
		15694: rom = 27;
		15695: rom = 27;
		15696: rom = 27;
		15697: rom = 27;
		15698: rom = 27;
		15699: rom = 27;
		15700: rom = 27;
		15701: rom = 27;
		15702: rom = 18;
		15703: rom = 7;
		15704: rom = 15;
		15705: rom = 13;
		15706: rom = 8;
		15707: rom = 21;
		15708: rom = 27;
		15709: rom = 27;
		15710: rom = 27;
		15711: rom = 23;
		15712: rom = 14;
		15713: rom = 18;
		15714: rom = 18;
		15715: rom = 18;
		15716: rom = 18;
		15717: rom = 18;
		15718: rom = 18;
		15719: rom = 18;
		15720: rom = 18;
		15721: rom = 18;
		15722: rom = 18;
		15723: rom = 18;
		15724: rom = 18;
		15725: rom = 18;
		15726: rom = 11;
		15727: rom = 18;
		15728: rom = 18;
		15729: rom = 18;
		15730: rom = 18;
		15731: rom = 18;
		15732: rom = 18;
		15733: rom = 16;
		15734: rom = 21;
		15735: rom = 27;
		15736: rom = 27;
		15737: rom = 27;
		15738: rom = 27;
		15744: rom = 27;
		15745: rom = 27;
		15746: rom = 27;
		15747: rom = 27;
		15748: rom = 27;
		15749: rom = 27;
		15750: rom = 27;
		15751: rom = 27;
		15752: rom = 27;
		15753: rom = 27;
		15754: rom = 27;
		15755: rom = 27;
		15756: rom = 27;
		15757: rom = 27;
		15758: rom = 27;
		15759: rom = 27;
		15760: rom = 27;
		15761: rom = 27;
		15762: rom = 27;
		15763: rom = 27;
		15764: rom = 27;
		15765: rom = 27;
		15766: rom = 27;
		15767: rom = 27;
		15768: rom = 27;
		15769: rom = 27;
		15770: rom = 27;
		15771: rom = 27;
		15772: rom = 27;
		15773: rom = 27;
		15774: rom = 27;
		15775: rom = 27;
		15776: rom = 27;
		15777: rom = 27;
		15778: rom = 27;
		15779: rom = 27;
		15780: rom = 27;
		15781: rom = 27;
		15782: rom = 27;
		15783: rom = 27;
		15784: rom = 27;
		15785: rom = 27;
		15786: rom = 27;
		15787: rom = 27;
		15788: rom = 27;
		15789: rom = 27;
		15790: rom = 27;
		15791: rom = 27;
		15792: rom = 27;
		15793: rom = 27;
		15794: rom = 27;
		15795: rom = 27;
		15796: rom = 27;
		15797: rom = 27;
		15798: rom = 27;
		15799: rom = 27;
		15800: rom = 27;
		15801: rom = 27;
		15802: rom = 27;
		15803: rom = 27;
		15804: rom = 27;
		15805: rom = 27;
		15806: rom = 27;
		15807: rom = 27;
		15808: rom = 27;
		15809: rom = 27;
		15810: rom = 27;
		15811: rom = 27;
		15812: rom = 27;
		15813: rom = 27;
		15814: rom = 27;
		15815: rom = 27;
		15816: rom = 27;
		15817: rom = 27;
		15818: rom = 27;
		15819: rom = 27;
		15820: rom = 27;
		15821: rom = 27;
		15822: rom = 27;
		15823: rom = 27;
		15824: rom = 27;
		15825: rom = 27;
		15826: rom = 27;
		15827: rom = 27;
		15828: rom = 27;
		15829: rom = 27;
		15830: rom = 27;
		15831: rom = 27;
		15832: rom = 22;
		15833: rom = 13;
		15834: rom = 5;
		15835: rom = 12;
		15836: rom = 27;
		15837: rom = 27;
		15838: rom = 27;
		15839: rom = 17;
		15840: rom = 17;
		15841: rom = 18;
		15842: rom = 18;
		15843: rom = 18;
		15844: rom = 18;
		15845: rom = 18;
		15846: rom = 18;
		15847: rom = 18;
		15848: rom = 18;
		15849: rom = 18;
		15850: rom = 18;
		15851: rom = 18;
		15852: rom = 18;
		15853: rom = 17;
		15854: rom = 12;
		15855: rom = 18;
		15856: rom = 18;
		15857: rom = 18;
		15858: rom = 18;
		15859: rom = 18;
		15860: rom = 18;
		15861: rom = 18;
		15862: rom = 13;
		15863: rom = 27;
		15864: rom = 27;
		15865: rom = 27;
		15866: rom = 27;
		15872: rom = 27;
		15873: rom = 27;
		15874: rom = 27;
		15875: rom = 27;
		15876: rom = 27;
		15877: rom = 27;
		15878: rom = 27;
		15879: rom = 27;
		15880: rom = 27;
		15881: rom = 27;
		15882: rom = 27;
		15883: rom = 27;
		15884: rom = 27;
		15885: rom = 27;
		15886: rom = 27;
		15887: rom = 27;
		15888: rom = 27;
		15889: rom = 27;
		15890: rom = 27;
		15891: rom = 27;
		15892: rom = 27;
		15893: rom = 27;
		15894: rom = 27;
		15895: rom = 27;
		15896: rom = 27;
		15897: rom = 27;
		15898: rom = 27;
		15899: rom = 27;
		15900: rom = 27;
		15901: rom = 27;
		15902: rom = 27;
		15903: rom = 27;
		15904: rom = 27;
		15905: rom = 27;
		15906: rom = 27;
		15907: rom = 27;
		15908: rom = 27;
		15909: rom = 27;
		15910: rom = 27;
		15911: rom = 27;
		15912: rom = 27;
		15913: rom = 27;
		15914: rom = 26;
		15915: rom = 23;
		15916: rom = 20;
		15917: rom = 16;
		15918: rom = 14;
		15919: rom = 13;
		15920: rom = 11;
		15921: rom = 14;
		15922: rom = 15;
		15923: rom = 19;
		15924: rom = 22;
		15925: rom = 26;
		15926: rom = 27;
		15927: rom = 27;
		15928: rom = 27;
		15929: rom = 27;
		15930: rom = 27;
		15931: rom = 27;
		15932: rom = 27;
		15933: rom = 27;
		15934: rom = 27;
		15935: rom = 27;
		15936: rom = 27;
		15937: rom = 27;
		15938: rom = 27;
		15939: rom = 27;
		15940: rom = 27;
		15941: rom = 27;
		15942: rom = 27;
		15943: rom = 27;
		15944: rom = 27;
		15945: rom = 27;
		15946: rom = 27;
		15947: rom = 27;
		15948: rom = 27;
		15949: rom = 27;
		15950: rom = 27;
		15951: rom = 27;
		15952: rom = 27;
		15953: rom = 27;
		15954: rom = 27;
		15955: rom = 27;
		15956: rom = 27;
		15957: rom = 27;
		15958: rom = 27;
		15959: rom = 27;
		15960: rom = 27;
		15961: rom = 27;
		15962: rom = 27;
		15963: rom = 27;
		15964: rom = 27;
		15965: rom = 27;
		15966: rom = 27;
		15967: rom = 12;
		15968: rom = 18;
		15969: rom = 18;
		15970: rom = 18;
		15971: rom = 18;
		15972: rom = 18;
		15973: rom = 18;
		15974: rom = 18;
		15975: rom = 18;
		15976: rom = 18;
		15977: rom = 18;
		15978: rom = 18;
		15979: rom = 18;
		15980: rom = 18;
		15981: rom = 15;
		15982: rom = 14;
		15983: rom = 18;
		15984: rom = 18;
		15985: rom = 18;
		15986: rom = 18;
		15987: rom = 18;
		15988: rom = 18;
		15989: rom = 18;
		15990: rom = 14;
		15991: rom = 24;
		15992: rom = 27;
		15993: rom = 27;
		15994: rom = 27;
		16000: rom = 27;
		16001: rom = 27;
		16002: rom = 27;
		16003: rom = 27;
		16004: rom = 27;
		16005: rom = 27;
		16006: rom = 27;
		16007: rom = 27;
		16008: rom = 27;
		16009: rom = 27;
		16010: rom = 27;
		16011: rom = 27;
		16012: rom = 27;
		16013: rom = 27;
		16014: rom = 27;
		16015: rom = 27;
		16016: rom = 27;
		16017: rom = 27;
		16018: rom = 27;
		16019: rom = 27;
		16020: rom = 27;
		16021: rom = 27;
		16022: rom = 27;
		16023: rom = 27;
		16024: rom = 27;
		16025: rom = 27;
		16026: rom = 27;
		16027: rom = 27;
		16028: rom = 27;
		16029: rom = 27;
		16030: rom = 27;
		16031: rom = 27;
		16032: rom = 27;
		16033: rom = 27;
		16034: rom = 27;
		16035: rom = 27;
		16036: rom = 27;
		16037: rom = 27;
		16038: rom = 27;
		16039: rom = 27;
		16040: rom = 24;
		16041: rom = 14;
		16042: rom = 9;
		16043: rom = 12;
		16044: rom = 15;
		16045: rom = 16;
		16046: rom = 17;
		16047: rom = 18;
		16048: rom = 18;
		16049: rom = 18;
		16050: rom = 17;
		16051: rom = 16;
		16052: rom = 14;
		16053: rom = 10;
		16054: rom = 13;
		16055: rom = 21;
		16056: rom = 26;
		16057: rom = 27;
		16058: rom = 27;
		16059: rom = 27;
		16060: rom = 27;
		16061: rom = 27;
		16062: rom = 27;
		16063: rom = 27;
		16064: rom = 27;
		16065: rom = 27;
		16066: rom = 27;
		16067: rom = 27;
		16068: rom = 27;
		16069: rom = 27;
		16070: rom = 27;
		16071: rom = 27;
		16072: rom = 27;
		16073: rom = 27;
		16074: rom = 27;
		16075: rom = 27;
		16076: rom = 27;
		16077: rom = 27;
		16078: rom = 27;
		16079: rom = 27;
		16080: rom = 27;
		16081: rom = 27;
		16082: rom = 27;
		16083: rom = 27;
		16084: rom = 27;
		16085: rom = 27;
		16086: rom = 27;
		16087: rom = 27;
		16088: rom = 27;
		16089: rom = 27;
		16090: rom = 27;
		16091: rom = 27;
		16092: rom = 27;
		16093: rom = 27;
		16094: rom = 22;
		16095: rom = 15;
		16096: rom = 18;
		16097: rom = 18;
		16098: rom = 18;
		16099: rom = 18;
		16100: rom = 18;
		16101: rom = 18;
		16102: rom = 18;
		16103: rom = 18;
		16104: rom = 18;
		16105: rom = 18;
		16106: rom = 18;
		16107: rom = 18;
		16108: rom = 18;
		16109: rom = 13;
		16110: rom = 17;
		16111: rom = 18;
		16112: rom = 18;
		16113: rom = 18;
		16114: rom = 18;
		16115: rom = 18;
		16116: rom = 18;
		16117: rom = 18;
		16118: rom = 18;
		16119: rom = 16;
		16120: rom = 27;
		16121: rom = 27;
		16122: rom = 27;
		16128: rom = 27;
		16129: rom = 27;
		16130: rom = 27;
		16131: rom = 27;
		16132: rom = 27;
		16133: rom = 27;
		16134: rom = 27;
		16135: rom = 27;
		16136: rom = 27;
		16137: rom = 27;
		16138: rom = 27;
		16139: rom = 27;
		16140: rom = 27;
		16141: rom = 27;
		16142: rom = 27;
		16143: rom = 27;
		16144: rom = 27;
		16145: rom = 27;
		16146: rom = 27;
		16147: rom = 27;
		16148: rom = 27;
		16149: rom = 27;
		16150: rom = 27;
		16151: rom = 27;
		16152: rom = 27;
		16153: rom = 27;
		16154: rom = 27;
		16155: rom = 27;
		16156: rom = 27;
		16157: rom = 27;
		16158: rom = 27;
		16159: rom = 27;
		16160: rom = 27;
		16161: rom = 27;
		16162: rom = 27;
		16163: rom = 27;
		16164: rom = 27;
		16165: rom = 27;
		16166: rom = 26;
		16167: rom = 16;
		16168: rom = 12;
		16169: rom = 16;
		16170: rom = 18;
		16171: rom = 18;
		16172: rom = 18;
		16173: rom = 18;
		16174: rom = 18;
		16175: rom = 18;
		16176: rom = 18;
		16177: rom = 18;
		16178: rom = 18;
		16179: rom = 18;
		16180: rom = 18;
		16181: rom = 18;
		16182: rom = 17;
		16183: rom = 14;
		16184: rom = 10;
		16185: rom = 17;
		16186: rom = 25;
		16187: rom = 27;
		16188: rom = 27;
		16189: rom = 27;
		16190: rom = 27;
		16191: rom = 27;
		16192: rom = 27;
		16193: rom = 27;
		16194: rom = 27;
		16195: rom = 27;
		16196: rom = 27;
		16197: rom = 27;
		16198: rom = 27;
		16199: rom = 27;
		16200: rom = 27;
		16201: rom = 27;
		16202: rom = 27;
		16203: rom = 27;
		16204: rom = 27;
		16205: rom = 27;
		16206: rom = 27;
		16207: rom = 27;
		16208: rom = 27;
		16209: rom = 27;
		16210: rom = 27;
		16211: rom = 27;
		16212: rom = 27;
		16213: rom = 27;
		16214: rom = 27;
		16215: rom = 27;
		16216: rom = 27;
		16217: rom = 27;
		16218: rom = 27;
		16219: rom = 27;
		16220: rom = 27;
		16221: rom = 27;
		16222: rom = 14;
		16223: rom = 17;
		16224: rom = 18;
		16225: rom = 18;
		16226: rom = 18;
		16227: rom = 18;
		16228: rom = 18;
		16229: rom = 18;
		16230: rom = 18;
		16231: rom = 18;
		16232: rom = 18;
		16233: rom = 18;
		16234: rom = 18;
		16235: rom = 18;
		16236: rom = 18;
		16237: rom = 9;
		16238: rom = 18;
		16239: rom = 18;
		16240: rom = 18;
		16241: rom = 18;
		16242: rom = 17;
		16243: rom = 18;
		16244: rom = 18;
		16245: rom = 18;
		16246: rom = 18;
		16247: rom = 12;
		16248: rom = 26;
		16249: rom = 27;
		16250: rom = 27;
		16256: rom = 27;
		16257: rom = 27;
		16258: rom = 27;
		16259: rom = 27;
		16260: rom = 27;
		16261: rom = 27;
		16262: rom = 27;
		16263: rom = 27;
		16264: rom = 27;
		16265: rom = 27;
		16266: rom = 27;
		16267: rom = 27;
		16268: rom = 27;
		16269: rom = 27;
		16270: rom = 27;
		16271: rom = 27;
		16272: rom = 27;
		16273: rom = 27;
		16274: rom = 27;
		16275: rom = 27;
		16276: rom = 27;
		16277: rom = 27;
		16278: rom = 27;
		16279: rom = 27;
		16280: rom = 27;
		16281: rom = 27;
		16282: rom = 27;
		16283: rom = 27;
		16284: rom = 27;
		16285: rom = 27;
		16286: rom = 27;
		16287: rom = 27;
		16288: rom = 27;
		16289: rom = 27;
		16290: rom = 27;
		16291: rom = 27;
		16292: rom = 27;
		16293: rom = 24;
		16294: rom = 11;
		16295: rom = 16;
		16296: rom = 18;
		16297: rom = 18;
		16298: rom = 18;
		16299: rom = 18;
		16300: rom = 18;
		16301: rom = 18;
		16302: rom = 18;
		16303: rom = 18;
		16304: rom = 18;
		16305: rom = 18;
		16306: rom = 18;
		16307: rom = 18;
		16308: rom = 18;
		16309: rom = 18;
		16310: rom = 18;
		16311: rom = 18;
		16312: rom = 18;
		16313: rom = 16;
		16314: rom = 11;
		16315: rom = 18;
		16316: rom = 26;
		16317: rom = 27;
		16318: rom = 27;
		16319: rom = 27;
		16320: rom = 27;
		16321: rom = 27;
		16322: rom = 27;
		16323: rom = 27;
		16324: rom = 27;
		16325: rom = 27;
		16326: rom = 27;
		16327: rom = 27;
		16328: rom = 27;
		16329: rom = 27;
		16330: rom = 27;
		16331: rom = 27;
		16332: rom = 27;
		16333: rom = 27;
		16334: rom = 27;
		16335: rom = 27;
		16336: rom = 27;
		16337: rom = 27;
		16338: rom = 27;
		16339: rom = 27;
		16340: rom = 27;
		16341: rom = 27;
		16342: rom = 27;
		16343: rom = 27;
		16344: rom = 27;
		16345: rom = 27;
		16346: rom = 27;
		16347: rom = 27;
		16348: rom = 27;
		16349: rom = 24;
		16350: rom = 13;
		16351: rom = 18;
		16352: rom = 18;
		16353: rom = 18;
		16354: rom = 18;
		16355: rom = 18;
		16356: rom = 18;
		16357: rom = 18;
		16358: rom = 18;
		16359: rom = 18;
		16360: rom = 18;
		16361: rom = 18;
		16362: rom = 18;
		16363: rom = 18;
		16364: rom = 17;
		16365: rom = 10;
		16366: rom = 15;
		16367: rom = 18;
		16368: rom = 18;
		16369: rom = 14;
		16370: rom = 16;
		16371: rom = 18;
		16372: rom = 18;
		16373: rom = 18;
		16374: rom = 18;
		16375: rom = 16;
		16376: rom = 22;
		16377: rom = 27;
		16378: rom = 27;
		16384: rom = 27;
		16385: rom = 27;
		16386: rom = 27;
		16387: rom = 27;
		16388: rom = 27;
		16389: rom = 27;
		16390: rom = 27;
		16391: rom = 27;
		16392: rom = 27;
		16393: rom = 27;
		16394: rom = 27;
		16395: rom = 27;
		16396: rom = 27;
		16397: rom = 27;
		16398: rom = 27;
		16399: rom = 27;
		16400: rom = 27;
		16401: rom = 27;
		16402: rom = 27;
		16403: rom = 27;
		16404: rom = 27;
		16405: rom = 27;
		16406: rom = 27;
		16407: rom = 27;
		16408: rom = 27;
		16409: rom = 27;
		16410: rom = 27;
		16411: rom = 27;
		16412: rom = 27;
		16413: rom = 27;
		16414: rom = 27;
		16415: rom = 27;
		16416: rom = 27;
		16417: rom = 27;
		16418: rom = 27;
		16419: rom = 27;
		16420: rom = 23;
		16421: rom = 11;
		16422: rom = 17;
		16423: rom = 18;
		16424: rom = 18;
		16425: rom = 18;
		16426: rom = 18;
		16427: rom = 18;
		16428: rom = 18;
		16429: rom = 18;
		16430: rom = 18;
		16431: rom = 18;
		16432: rom = 18;
		16433: rom = 18;
		16434: rom = 18;
		16435: rom = 18;
		16436: rom = 18;
		16437: rom = 18;
		16438: rom = 18;
		16439: rom = 18;
		16440: rom = 18;
		16441: rom = 18;
		16442: rom = 18;
		16443: rom = 16;
		16444: rom = 11;
		16445: rom = 21;
		16446: rom = 27;
		16447: rom = 27;
		16448: rom = 27;
		16449: rom = 27;
		16450: rom = 27;
		16451: rom = 27;
		16452: rom = 27;
		16453: rom = 27;
		16454: rom = 27;
		16455: rom = 27;
		16456: rom = 27;
		16457: rom = 27;
		16458: rom = 27;
		16459: rom = 27;
		16460: rom = 27;
		16461: rom = 27;
		16462: rom = 27;
		16463: rom = 27;
		16464: rom = 27;
		16465: rom = 27;
		16466: rom = 27;
		16467: rom = 27;
		16468: rom = 27;
		16469: rom = 27;
		16470: rom = 27;
		16471: rom = 27;
		16472: rom = 27;
		16473: rom = 27;
		16474: rom = 27;
		16475: rom = 27;
		16476: rom = 27;
		16477: rom = 14;
		16478: rom = 17;
		16479: rom = 18;
		16480: rom = 18;
		16481: rom = 18;
		16482: rom = 18;
		16483: rom = 18;
		16484: rom = 18;
		16485: rom = 18;
		16486: rom = 18;
		16487: rom = 18;
		16488: rom = 18;
		16489: rom = 18;
		16490: rom = 18;
		16491: rom = 18;
		16492: rom = 14;
		16493: rom = 23;
		16494: rom = 12;
		16495: rom = 18;
		16496: rom = 18;
		16497: rom = 12;
		16498: rom = 18;
		16499: rom = 18;
		16500: rom = 18;
		16501: rom = 18;
		16502: rom = 18;
		16503: rom = 17;
		16504: rom = 19;
		16505: rom = 27;
		16506: rom = 27;
		16512: rom = 27;
		16513: rom = 27;
		16514: rom = 27;
		16515: rom = 27;
		16516: rom = 27;
		16517: rom = 27;
		16518: rom = 27;
		16519: rom = 27;
		16520: rom = 27;
		16521: rom = 27;
		16522: rom = 27;
		16523: rom = 27;
		16524: rom = 27;
		16525: rom = 27;
		16526: rom = 27;
		16527: rom = 27;
		16528: rom = 27;
		16529: rom = 27;
		16530: rom = 27;
		16531: rom = 27;
		16532: rom = 27;
		16533: rom = 27;
		16534: rom = 27;
		16535: rom = 27;
		16536: rom = 27;
		16537: rom = 27;
		16538: rom = 27;
		16539: rom = 27;
		16540: rom = 27;
		16541: rom = 27;
		16542: rom = 27;
		16543: rom = 27;
		16544: rom = 27;
		16545: rom = 27;
		16546: rom = 27;
		16547: rom = 26;
		16548: rom = 12;
		16549: rom = 17;
		16550: rom = 18;
		16551: rom = 18;
		16552: rom = 18;
		16553: rom = 18;
		16554: rom = 18;
		16555: rom = 18;
		16556: rom = 18;
		16557: rom = 18;
		16558: rom = 18;
		16559: rom = 18;
		16560: rom = 18;
		16561: rom = 18;
		16562: rom = 18;
		16563: rom = 18;
		16564: rom = 18;
		16565: rom = 18;
		16566: rom = 18;
		16567: rom = 18;
		16568: rom = 18;
		16569: rom = 18;
		16570: rom = 18;
		16571: rom = 18;
		16572: rom = 17;
		16573: rom = 13;
		16574: rom = 15;
		16575: rom = 26;
		16576: rom = 27;
		16577: rom = 27;
		16578: rom = 27;
		16579: rom = 27;
		16580: rom = 27;
		16581: rom = 27;
		16582: rom = 27;
		16583: rom = 27;
		16584: rom = 27;
		16585: rom = 27;
		16586: rom = 27;
		16587: rom = 27;
		16588: rom = 27;
		16589: rom = 27;
		16590: rom = 27;
		16591: rom = 27;
		16592: rom = 27;
		16593: rom = 27;
		16594: rom = 27;
		16595: rom = 27;
		16596: rom = 27;
		16597: rom = 27;
		16598: rom = 27;
		16599: rom = 27;
		16600: rom = 27;
		16601: rom = 27;
		16602: rom = 27;
		16603: rom = 27;
		16604: rom = 22;
		16605: rom = 13;
		16606: rom = 18;
		16607: rom = 18;
		16608: rom = 18;
		16609: rom = 18;
		16610: rom = 18;
		16611: rom = 18;
		16612: rom = 18;
		16613: rom = 18;
		16614: rom = 18;
		16615: rom = 18;
		16616: rom = 18;
		16617: rom = 18;
		16618: rom = 18;
		16619: rom = 18;
		16620: rom = 12;
		16621: rom = 27;
		16622: rom = 12;
		16623: rom = 18;
		16624: rom = 18;
		16625: rom = 11;
		16626: rom = 18;
		16627: rom = 18;
		16628: rom = 18;
		16629: rom = 18;
		16630: rom = 18;
		16631: rom = 17;
		16632: rom = 20;
		16633: rom = 27;
		16634: rom = 27;
		16640: rom = 27;
		16641: rom = 27;
		16642: rom = 27;
		16643: rom = 27;
		16644: rom = 27;
		16645: rom = 27;
		16646: rom = 27;
		16647: rom = 27;
		16648: rom = 27;
		16649: rom = 27;
		16650: rom = 27;
		16651: rom = 27;
		16652: rom = 27;
		16653: rom = 27;
		16654: rom = 27;
		16655: rom = 27;
		16656: rom = 27;
		16657: rom = 27;
		16658: rom = 27;
		16659: rom = 27;
		16660: rom = 27;
		16661: rom = 27;
		16662: rom = 27;
		16663: rom = 27;
		16664: rom = 27;
		16665: rom = 27;
		16666: rom = 27;
		16667: rom = 27;
		16668: rom = 27;
		16669: rom = 27;
		16670: rom = 27;
		16671: rom = 27;
		16672: rom = 27;
		16673: rom = 27;
		16674: rom = 27;
		16675: rom = 14;
		16676: rom = 17;
		16677: rom = 18;
		16678: rom = 18;
		16679: rom = 18;
		16680: rom = 18;
		16681: rom = 18;
		16682: rom = 18;
		16683: rom = 18;
		16684: rom = 18;
		16685: rom = 18;
		16686: rom = 18;
		16687: rom = 18;
		16688: rom = 18;
		16689: rom = 18;
		16690: rom = 18;
		16691: rom = 18;
		16692: rom = 18;
		16693: rom = 18;
		16694: rom = 18;
		16695: rom = 18;
		16696: rom = 18;
		16697: rom = 18;
		16698: rom = 18;
		16699: rom = 18;
		16700: rom = 18;
		16701: rom = 18;
		16702: rom = 16;
		16703: rom = 11;
		16704: rom = 22;
		16705: rom = 27;
		16706: rom = 27;
		16707: rom = 27;
		16708: rom = 27;
		16709: rom = 27;
		16710: rom = 27;
		16711: rom = 27;
		16712: rom = 27;
		16713: rom = 27;
		16714: rom = 27;
		16715: rom = 27;
		16716: rom = 27;
		16717: rom = 27;
		16718: rom = 27;
		16719: rom = 27;
		16720: rom = 27;
		16721: rom = 27;
		16722: rom = 27;
		16723: rom = 27;
		16724: rom = 27;
		16725: rom = 27;
		16726: rom = 27;
		16727: rom = 27;
		16728: rom = 27;
		16729: rom = 27;
		16730: rom = 27;
		16731: rom = 26;
		16732: rom = 12;
		16733: rom = 17;
		16734: rom = 18;
		16735: rom = 18;
		16736: rom = 18;
		16737: rom = 18;
		16738: rom = 18;
		16739: rom = 18;
		16740: rom = 18;
		16741: rom = 18;
		16742: rom = 18;
		16743: rom = 18;
		16744: rom = 18;
		16745: rom = 18;
		16746: rom = 18;
		16747: rom = 16;
		16748: rom = 20;
		16749: rom = 27;
		16750: rom = 16;
		16751: rom = 18;
		16752: rom = 18;
		16753: rom = 12;
		16754: rom = 17;
		16755: rom = 18;
		16756: rom = 10;
		16757: rom = 10;
		16758: rom = 10;
		16759: rom = 8;
		16760: rom = 14;
		16761: rom = 22;
		16762: rom = 27;
		16768: rom = 27;
		16769: rom = 27;
		16770: rom = 27;
		16771: rom = 27;
		16772: rom = 27;
		16773: rom = 27;
		16774: rom = 27;
		16775: rom = 27;
		16776: rom = 27;
		16777: rom = 27;
		16778: rom = 27;
		16779: rom = 27;
		16780: rom = 27;
		16781: rom = 27;
		16782: rom = 27;
		16783: rom = 27;
		16784: rom = 27;
		16785: rom = 27;
		16786: rom = 27;
		16787: rom = 27;
		16788: rom = 27;
		16789: rom = 27;
		16790: rom = 27;
		16791: rom = 27;
		16792: rom = 27;
		16793: rom = 27;
		16794: rom = 27;
		16795: rom = 27;
		16796: rom = 27;
		16797: rom = 27;
		16798: rom = 27;
		16799: rom = 27;
		16800: rom = 27;
		16801: rom = 27;
		16802: rom = 22;
		16803: rom = 14;
		16804: rom = 18;
		16805: rom = 18;
		16806: rom = 18;
		16807: rom = 18;
		16808: rom = 18;
		16809: rom = 18;
		16810: rom = 18;
		16811: rom = 17;
		16812: rom = 16;
		16813: rom = 16;
		16814: rom = 17;
		16815: rom = 18;
		16816: rom = 18;
		16817: rom = 18;
		16818: rom = 18;
		16819: rom = 18;
		16820: rom = 18;
		16821: rom = 18;
		16822: rom = 18;
		16823: rom = 18;
		16824: rom = 18;
		16825: rom = 18;
		16826: rom = 18;
		16827: rom = 18;
		16828: rom = 18;
		16829: rom = 18;
		16830: rom = 18;
		16831: rom = 17;
		16832: rom = 12;
		16833: rom = 18;
		16834: rom = 27;
		16835: rom = 27;
		16836: rom = 27;
		16837: rom = 27;
		16838: rom = 27;
		16839: rom = 27;
		16840: rom = 27;
		16841: rom = 27;
		16842: rom = 27;
		16843: rom = 27;
		16844: rom = 27;
		16845: rom = 27;
		16846: rom = 27;
		16847: rom = 27;
		16848: rom = 27;
		16849: rom = 27;
		16850: rom = 27;
		16851: rom = 27;
		16852: rom = 27;
		16853: rom = 27;
		16854: rom = 27;
		16855: rom = 27;
		16856: rom = 27;
		16857: rom = 27;
		16858: rom = 27;
		16859: rom = 16;
		16860: rom = 16;
		16861: rom = 18;
		16862: rom = 18;
		16863: rom = 18;
		16864: rom = 18;
		16865: rom = 18;
		16866: rom = 18;
		16867: rom = 18;
		16868: rom = 18;
		16869: rom = 18;
		16870: rom = 18;
		16871: rom = 18;
		16872: rom = 18;
		16873: rom = 18;
		16874: rom = 18;
		16875: rom = 11;
		16876: rom = 26;
		16877: rom = 27;
		16878: rom = 16;
		16879: rom = 18;
		16880: rom = 18;
		16881: rom = 16;
		16882: rom = 12;
		16883: rom = 17;
		16884: rom = 10;
		16885: rom = 16;
		16886: rom = 15;
		16887: rom = 11;
		16888: rom = 19;
		16889: rom = 27;
		16890: rom = 27;
		16896: rom = 27;
		16897: rom = 27;
		16898: rom = 27;
		16899: rom = 27;
		16900: rom = 27;
		16901: rom = 27;
		16902: rom = 27;
		16903: rom = 27;
		16904: rom = 27;
		16905: rom = 27;
		16906: rom = 27;
		16907: rom = 27;
		16908: rom = 27;
		16909: rom = 27;
		16910: rom = 27;
		16911: rom = 27;
		16912: rom = 27;
		16913: rom = 27;
		16914: rom = 27;
		16915: rom = 27;
		16916: rom = 27;
		16917: rom = 27;
		16918: rom = 27;
		16919: rom = 27;
		16920: rom = 27;
		16921: rom = 27;
		16922: rom = 27;
		16923: rom = 27;
		16924: rom = 27;
		16925: rom = 27;
		16926: rom = 27;
		16927: rom = 27;
		16928: rom = 27;
		16929: rom = 27;
		16930: rom = 13;
		16931: rom = 17;
		16932: rom = 18;
		16933: rom = 18;
		16934: rom = 18;
		16935: rom = 18;
		16936: rom = 18;
		16937: rom = 16;
		16938: rom = 11;
		16939: rom = 16;
		16940: rom = 19;
		16941: rom = 19;
		16942: rom = 16;
		16943: rom = 13;
		16944: rom = 10;
		16945: rom = 14;
		16946: rom = 17;
		16947: rom = 18;
		16948: rom = 18;
		16949: rom = 18;
		16950: rom = 18;
		16951: rom = 18;
		16952: rom = 18;
		16953: rom = 18;
		16954: rom = 18;
		16955: rom = 18;
		16956: rom = 18;
		16957: rom = 18;
		16958: rom = 18;
		16959: rom = 18;
		16960: rom = 18;
		16961: rom = 15;
		16962: rom = 13;
		16963: rom = 25;
		16964: rom = 27;
		16965: rom = 27;
		16966: rom = 27;
		16967: rom = 27;
		16968: rom = 27;
		16969: rom = 27;
		16970: rom = 27;
		16971: rom = 27;
		16972: rom = 27;
		16973: rom = 27;
		16974: rom = 27;
		16975: rom = 27;
		16976: rom = 27;
		16977: rom = 27;
		16978: rom = 27;
		16979: rom = 27;
		16980: rom = 27;
		16981: rom = 27;
		16982: rom = 27;
		16983: rom = 27;
		16984: rom = 27;
		16985: rom = 27;
		16986: rom = 19;
		16987: rom = 14;
		16988: rom = 18;
		16989: rom = 18;
		16990: rom = 18;
		16991: rom = 18;
		16992: rom = 18;
		16993: rom = 18;
		16994: rom = 18;
		16995: rom = 18;
		16996: rom = 18;
		16997: rom = 18;
		16998: rom = 18;
		16999: rom = 18;
		17000: rom = 18;
		17001: rom = 18;
		17002: rom = 16;
		17003: rom = 18;
		17004: rom = 27;
		17005: rom = 27;
		17006: rom = 16;
		17007: rom = 18;
		17008: rom = 18;
		17009: rom = 18;
		17010: rom = 14;
		17011: rom = 9;
		17012: rom = 7;
		17013: rom = 9;
		17014: rom = 10;
		17015: rom = 23;
		17016: rom = 27;
		17017: rom = 27;
		17018: rom = 27;
		17024: rom = 27;
		17025: rom = 27;
		17026: rom = 27;
		17027: rom = 27;
		17028: rom = 27;
		17029: rom = 27;
		17030: rom = 27;
		17031: rom = 27;
		17032: rom = 27;
		17033: rom = 27;
		17034: rom = 27;
		17035: rom = 27;
		17036: rom = 27;
		17037: rom = 27;
		17038: rom = 27;
		17039: rom = 27;
		17040: rom = 27;
		17041: rom = 27;
		17042: rom = 27;
		17043: rom = 27;
		17044: rom = 27;
		17045: rom = 27;
		17046: rom = 27;
		17047: rom = 27;
		17048: rom = 27;
		17049: rom = 27;
		17050: rom = 27;
		17051: rom = 27;
		17052: rom = 27;
		17053: rom = 27;
		17054: rom = 27;
		17055: rom = 27;
		17056: rom = 27;
		17057: rom = 24;
		17058: rom = 13;
		17059: rom = 18;
		17060: rom = 18;
		17061: rom = 18;
		17062: rom = 18;
		17063: rom = 18;
		17064: rom = 16;
		17065: rom = 14;
		17066: rom = 26;
		17067: rom = 27;
		17068: rom = 27;
		17069: rom = 27;
		17070: rom = 27;
		17071: rom = 27;
		17072: rom = 27;
		17073: rom = 23;
		17074: rom = 16;
		17075: rom = 11;
		17076: rom = 16;
		17077: rom = 18;
		17078: rom = 18;
		17079: rom = 18;
		17080: rom = 18;
		17081: rom = 18;
		17082: rom = 18;
		17083: rom = 18;
		17084: rom = 18;
		17085: rom = 18;
		17086: rom = 18;
		17087: rom = 18;
		17088: rom = 18;
		17089: rom = 18;
		17090: rom = 17;
		17091: rom = 11;
		17092: rom = 19;
		17093: rom = 27;
		17094: rom = 27;
		17095: rom = 27;
		17096: rom = 27;
		17097: rom = 27;
		17098: rom = 27;
		17099: rom = 27;
		17100: rom = 27;
		17101: rom = 27;
		17102: rom = 27;
		17103: rom = 27;
		17104: rom = 27;
		17105: rom = 27;
		17106: rom = 27;
		17107: rom = 27;
		17108: rom = 27;
		17109: rom = 27;
		17110: rom = 27;
		17111: rom = 27;
		17112: rom = 27;
		17113: rom = 19;
		17114: rom = 13;
		17115: rom = 18;
		17116: rom = 18;
		17117: rom = 18;
		17118: rom = 18;
		17119: rom = 18;
		17120: rom = 18;
		17121: rom = 18;
		17122: rom = 18;
		17123: rom = 18;
		17124: rom = 18;
		17125: rom = 18;
		17126: rom = 18;
		17127: rom = 18;
		17128: rom = 18;
		17129: rom = 18;
		17130: rom = 11;
		17131: rom = 26;
		17132: rom = 27;
		17133: rom = 27;
		17134: rom = 17;
		17135: rom = 18;
		17136: rom = 15;
		17137: rom = 15;
		17138: rom = 18;
		17139: rom = 18;
		17140: rom = 18;
		17141: rom = 18;
		17142: rom = 18;
		17143: rom = 15;
		17144: rom = 27;
		17145: rom = 27;
		17146: rom = 27;
		17152: rom = 27;
		17153: rom = 27;
		17154: rom = 27;
		17155: rom = 27;
		17156: rom = 27;
		17157: rom = 27;
		17158: rom = 27;
		17159: rom = 27;
		17160: rom = 27;
		17161: rom = 27;
		17162: rom = 27;
		17163: rom = 27;
		17164: rom = 27;
		17165: rom = 27;
		17166: rom = 27;
		17167: rom = 27;
		17168: rom = 27;
		17169: rom = 27;
		17170: rom = 27;
		17171: rom = 27;
		17172: rom = 27;
		17173: rom = 27;
		17174: rom = 27;
		17175: rom = 27;
		17176: rom = 27;
		17177: rom = 27;
		17178: rom = 27;
		17179: rom = 27;
		17180: rom = 27;
		17181: rom = 27;
		17182: rom = 27;
		17183: rom = 27;
		17184: rom = 27;
		17185: rom = 18;
		17186: rom = 17;
		17187: rom = 18;
		17188: rom = 18;
		17189: rom = 18;
		17190: rom = 18;
		17191: rom = 17;
		17192: rom = 13;
		17193: rom = 27;
		17194: rom = 27;
		17195: rom = 27;
		17196: rom = 27;
		17197: rom = 27;
		17198: rom = 27;
		17199: rom = 27;
		17200: rom = 27;
		17201: rom = 27;
		17202: rom = 27;
		17203: rom = 25;
		17204: rom = 18;
		17205: rom = 11;
		17206: rom = 16;
		17207: rom = 18;
		17208: rom = 18;
		17209: rom = 18;
		17210: rom = 18;
		17211: rom = 18;
		17212: rom = 18;
		17213: rom = 18;
		17214: rom = 18;
		17215: rom = 18;
		17216: rom = 18;
		17217: rom = 18;
		17218: rom = 18;
		17219: rom = 18;
		17220: rom = 15;
		17221: rom = 12;
		17222: rom = 23;
		17223: rom = 27;
		17224: rom = 27;
		17225: rom = 27;
		17226: rom = 27;
		17227: rom = 27;
		17228: rom = 27;
		17229: rom = 27;
		17230: rom = 27;
		17231: rom = 27;
		17232: rom = 27;
		17233: rom = 27;
		17234: rom = 27;
		17235: rom = 27;
		17236: rom = 27;
		17237: rom = 27;
		17238: rom = 27;
		17239: rom = 27;
		17240: rom = 17;
		17241: rom = 13;
		17242: rom = 18;
		17243: rom = 18;
		17244: rom = 18;
		17245: rom = 18;
		17246: rom = 18;
		17247: rom = 18;
		17248: rom = 18;
		17249: rom = 18;
		17250: rom = 18;
		17251: rom = 18;
		17252: rom = 18;
		17253: rom = 18;
		17254: rom = 18;
		17255: rom = 18;
		17256: rom = 18;
		17257: rom = 15;
		17258: rom = 19;
		17259: rom = 27;
		17260: rom = 27;
		17261: rom = 27;
		17262: rom = 18;
		17263: rom = 18;
		17264: rom = 11;
		17265: rom = 18;
		17266: rom = 18;
		17267: rom = 18;
		17268: rom = 16;
		17269: rom = 15;
		17270: rom = 15;
		17271: rom = 11;
		17272: rom = 17;
		17273: rom = 27;
		17274: rom = 27;
		17280: rom = 27;
		17281: rom = 27;
		17282: rom = 27;
		17283: rom = 27;
		17284: rom = 27;
		17285: rom = 27;
		17286: rom = 27;
		17287: rom = 27;
		17288: rom = 27;
		17289: rom = 27;
		17290: rom = 27;
		17291: rom = 27;
		17292: rom = 27;
		17293: rom = 27;
		17294: rom = 27;
		17295: rom = 27;
		17296: rom = 27;
		17297: rom = 27;
		17298: rom = 27;
		17299: rom = 27;
		17300: rom = 27;
		17301: rom = 27;
		17302: rom = 27;
		17303: rom = 27;
		17304: rom = 27;
		17305: rom = 27;
		17306: rom = 27;
		17307: rom = 27;
		17308: rom = 27;
		17309: rom = 27;
		17310: rom = 27;
		17311: rom = 27;
		17312: rom = 27;
		17313: rom = 13;
		17314: rom = 18;
		17315: rom = 18;
		17316: rom = 18;
		17317: rom = 18;
		17318: rom = 18;
		17319: rom = 14;
		17320: rom = 23;
		17321: rom = 27;
		17322: rom = 27;
		17323: rom = 27;
		17324: rom = 27;
		17325: rom = 27;
		17326: rom = 27;
		17327: rom = 27;
		17328: rom = 27;
		17329: rom = 27;
		17330: rom = 27;
		17331: rom = 27;
		17332: rom = 27;
		17333: rom = 26;
		17334: rom = 17;
		17335: rom = 12;
		17336: rom = 17;
		17337: rom = 18;
		17338: rom = 18;
		17339: rom = 18;
		17340: rom = 18;
		17341: rom = 18;
		17342: rom = 18;
		17343: rom = 18;
		17344: rom = 18;
		17345: rom = 18;
		17346: rom = 18;
		17347: rom = 18;
		17348: rom = 18;
		17349: rom = 17;
		17350: rom = 13;
		17351: rom = 13;
		17352: rom = 23;
		17353: rom = 27;
		17354: rom = 27;
		17355: rom = 27;
		17356: rom = 27;
		17357: rom = 27;
		17358: rom = 27;
		17359: rom = 27;
		17360: rom = 27;
		17361: rom = 27;
		17362: rom = 27;
		17363: rom = 27;
		17364: rom = 27;
		17365: rom = 27;
		17366: rom = 23;
		17367: rom = 12;
		17368: rom = 15;
		17369: rom = 18;
		17370: rom = 18;
		17371: rom = 18;
		17372: rom = 18;
		17373: rom = 18;
		17374: rom = 18;
		17375: rom = 18;
		17376: rom = 18;
		17377: rom = 18;
		17378: rom = 18;
		17379: rom = 18;
		17380: rom = 18;
		17381: rom = 18;
		17382: rom = 18;
		17383: rom = 18;
		17384: rom = 17;
		17385: rom = 12;
		17386: rom = 21;
		17387: rom = 27;
		17388: rom = 27;
		17389: rom = 27;
		17390: rom = 20;
		17391: rom = 17;
		17392: rom = 11;
		17393: rom = 18;
		17394: rom = 18;
		17395: rom = 7;
		17396: rom = 13;
		17397: rom = 14;
		17398: rom = 10;
		17399: rom = 7;
		17400: rom = 23;
		17401: rom = 27;
		17402: rom = 27;
		17408: rom = 27;
		17409: rom = 27;
		17410: rom = 27;
		17411: rom = 27;
		17412: rom = 27;
		17413: rom = 27;
		17414: rom = 27;
		17415: rom = 27;
		17416: rom = 27;
		17417: rom = 27;
		17418: rom = 27;
		17419: rom = 27;
		17420: rom = 27;
		17421: rom = 27;
		17422: rom = 27;
		17423: rom = 27;
		17424: rom = 27;
		17425: rom = 27;
		17426: rom = 27;
		17427: rom = 27;
		17428: rom = 27;
		17429: rom = 27;
		17430: rom = 27;
		17431: rom = 27;
		17432: rom = 27;
		17433: rom = 27;
		17434: rom = 27;
		17435: rom = 27;
		17436: rom = 27;
		17437: rom = 27;
		17438: rom = 27;
		17439: rom = 27;
		17440: rom = 26;
		17441: rom = 12;
		17442: rom = 18;
		17443: rom = 18;
		17444: rom = 18;
		17445: rom = 18;
		17446: rom = 18;
		17447: rom = 12;
		17448: rom = 27;
		17449: rom = 27;
		17450: rom = 27;
		17451: rom = 27;
		17452: rom = 27;
		17453: rom = 27;
		17454: rom = 27;
		17455: rom = 27;
		17456: rom = 27;
		17457: rom = 27;
		17458: rom = 27;
		17459: rom = 27;
		17460: rom = 27;
		17461: rom = 27;
		17462: rom = 27;
		17463: rom = 24;
		17464: rom = 13;
		17465: rom = 15;
		17466: rom = 18;
		17467: rom = 18;
		17468: rom = 18;
		17469: rom = 18;
		17470: rom = 18;
		17471: rom = 18;
		17472: rom = 18;
		17473: rom = 18;
		17474: rom = 18;
		17475: rom = 18;
		17476: rom = 18;
		17477: rom = 18;
		17478: rom = 18;
		17479: rom = 17;
		17480: rom = 13;
		17481: rom = 12;
		17482: rom = 20;
		17483: rom = 26;
		17484: rom = 27;
		17485: rom = 27;
		17486: rom = 27;
		17487: rom = 27;
		17488: rom = 27;
		17489: rom = 27;
		17490: rom = 27;
		17491: rom = 27;
		17492: rom = 22;
		17493: rom = 14;
		17494: rom = 12;
		17495: rom = 17;
		17496: rom = 18;
		17497: rom = 18;
		17498: rom = 18;
		17499: rom = 18;
		17500: rom = 18;
		17501: rom = 18;
		17502: rom = 18;
		17503: rom = 18;
		17504: rom = 18;
		17505: rom = 18;
		17506: rom = 18;
		17507: rom = 18;
		17508: rom = 18;
		17509: rom = 18;
		17510: rom = 18;
		17511: rom = 18;
		17512: rom = 12;
		17513: rom = 24;
		17514: rom = 27;
		17515: rom = 27;
		17516: rom = 27;
		17517: rom = 27;
		17518: rom = 19;
		17519: rom = 16;
		17520: rom = 14;
		17521: rom = 15;
		17522: rom = 18;
		17523: rom = 13;
		17524: rom = 10;
		17525: rom = 9;
		17526: rom = 3;
		17527: rom = 23;
		17528: rom = 27;
		17529: rom = 27;
		17530: rom = 27;
		17536: rom = 27;
		17537: rom = 27;
		17538: rom = 27;
		17539: rom = 27;
		17540: rom = 27;
		17541: rom = 27;
		17542: rom = 27;
		17543: rom = 27;
		17544: rom = 27;
		17545: rom = 27;
		17546: rom = 27;
		17547: rom = 27;
		17548: rom = 27;
		17549: rom = 27;
		17550: rom = 27;
		17551: rom = 27;
		17552: rom = 27;
		17553: rom = 27;
		17554: rom = 27;
		17555: rom = 27;
		17556: rom = 27;
		17557: rom = 27;
		17558: rom = 27;
		17559: rom = 27;
		17560: rom = 27;
		17561: rom = 27;
		17562: rom = 27;
		17563: rom = 27;
		17564: rom = 27;
		17565: rom = 27;
		17566: rom = 27;
		17567: rom = 27;
		17568: rom = 24;
		17569: rom = 13;
		17570: rom = 18;
		17571: rom = 18;
		17572: rom = 18;
		17573: rom = 18;
		17574: rom = 18;
		17575: rom = 15;
		17576: rom = 27;
		17577: rom = 27;
		17578: rom = 27;
		17579: rom = 27;
		17580: rom = 27;
		17581: rom = 27;
		17582: rom = 27;
		17583: rom = 27;
		17584: rom = 27;
		17585: rom = 27;
		17586: rom = 27;
		17587: rom = 27;
		17588: rom = 27;
		17589: rom = 27;
		17590: rom = 27;
		17591: rom = 27;
		17592: rom = 27;
		17593: rom = 19;
		17594: rom = 11;
		17595: rom = 17;
		17596: rom = 18;
		17597: rom = 18;
		17598: rom = 18;
		17599: rom = 18;
		17600: rom = 18;
		17601: rom = 18;
		17602: rom = 18;
		17603: rom = 18;
		17604: rom = 18;
		17605: rom = 18;
		17606: rom = 18;
		17607: rom = 18;
		17608: rom = 18;
		17609: rom = 17;
		17610: rom = 15;
		17611: rom = 11;
		17612: rom = 13;
		17613: rom = 18;
		17614: rom = 21;
		17615: rom = 21;
		17616: rom = 20;
		17617: rom = 18;
		17618: rom = 14;
		17619: rom = 10;
		17620: rom = 14;
		17621: rom = 17;
		17622: rom = 18;
		17623: rom = 18;
		17624: rom = 18;
		17625: rom = 18;
		17626: rom = 18;
		17627: rom = 18;
		17628: rom = 18;
		17629: rom = 18;
		17630: rom = 18;
		17631: rom = 18;
		17632: rom = 18;
		17633: rom = 18;
		17634: rom = 18;
		17635: rom = 18;
		17636: rom = 18;
		17637: rom = 18;
		17638: rom = 18;
		17639: rom = 15;
		17640: rom = 18;
		17641: rom = 26;
		17642: rom = 27;
		17643: rom = 27;
		17644: rom = 27;
		17645: rom = 27;
		17646: rom = 21;
		17647: rom = 13;
		17648: rom = 18;
		17649: rom = 12;
		17650: rom = 10;
		17651: rom = 11;
		17652: rom = 9;
		17653: rom = 7;
		17654: rom = 22;
		17655: rom = 27;
		17656: rom = 27;
		17657: rom = 27;
		17658: rom = 27;
		17664: rom = 27;
		17665: rom = 27;
		17666: rom = 27;
		17667: rom = 27;
		17668: rom = 27;
		17669: rom = 27;
		17670: rom = 27;
		17671: rom = 27;
		17672: rom = 27;
		17673: rom = 27;
		17674: rom = 27;
		17675: rom = 27;
		17676: rom = 27;
		17677: rom = 27;
		17678: rom = 27;
		17679: rom = 27;
		17680: rom = 27;
		17681: rom = 27;
		17682: rom = 27;
		17683: rom = 27;
		17684: rom = 27;
		17685: rom = 27;
		17686: rom = 27;
		17687: rom = 27;
		17688: rom = 27;
		17689: rom = 27;
		17690: rom = 27;
		17691: rom = 27;
		17692: rom = 27;
		17693: rom = 27;
		17694: rom = 27;
		17695: rom = 27;
		17696: rom = 23;
		17697: rom = 14;
		17698: rom = 18;
		17699: rom = 18;
		17700: rom = 18;
		17701: rom = 18;
		17702: rom = 18;
		17703: rom = 16;
		17704: rom = 27;
		17705: rom = 27;
		17706: rom = 27;
		17707: rom = 27;
		17708: rom = 27;
		17709: rom = 27;
		17710: rom = 27;
		17711: rom = 27;
		17712: rom = 27;
		17713: rom = 27;
		17714: rom = 27;
		17715: rom = 27;
		17716: rom = 27;
		17717: rom = 27;
		17718: rom = 27;
		17719: rom = 27;
		17720: rom = 27;
		17721: rom = 27;
		17722: rom = 23;
		17723: rom = 11;
		17724: rom = 16;
		17725: rom = 18;
		17726: rom = 18;
		17727: rom = 18;
		17728: rom = 18;
		17729: rom = 18;
		17730: rom = 18;
		17731: rom = 18;
		17732: rom = 18;
		17733: rom = 18;
		17734: rom = 18;
		17735: rom = 18;
		17736: rom = 18;
		17737: rom = 18;
		17738: rom = 18;
		17739: rom = 18;
		17740: rom = 17;
		17741: rom = 16;
		17742: rom = 15;
		17743: rom = 14;
		17744: rom = 15;
		17745: rom = 16;
		17746: rom = 17;
		17747: rom = 18;
		17748: rom = 18;
		17749: rom = 18;
		17750: rom = 18;
		17751: rom = 18;
		17752: rom = 18;
		17753: rom = 18;
		17754: rom = 18;
		17755: rom = 18;
		17756: rom = 18;
		17757: rom = 18;
		17758: rom = 18;
		17759: rom = 18;
		17760: rom = 18;
		17761: rom = 18;
		17762: rom = 18;
		17763: rom = 18;
		17764: rom = 18;
		17765: rom = 18;
		17766: rom = 17;
		17767: rom = 14;
		17768: rom = 27;
		17769: rom = 27;
		17770: rom = 27;
		17771: rom = 27;
		17772: rom = 27;
		17773: rom = 27;
		17774: rom = 26;
		17775: rom = 16;
		17776: rom = 16;
		17777: rom = 13;
		17778: rom = 9;
		17779: rom = 8;
		17780: rom = 10;
		17781: rom = 5;
		17782: rom = 25;
		17783: rom = 27;
		17784: rom = 27;
		17785: rom = 27;
		17786: rom = 27;
		17792: rom = 27;
		17793: rom = 27;
		17794: rom = 27;
		17795: rom = 27;
		17796: rom = 27;
		17797: rom = 27;
		17798: rom = 27;
		17799: rom = 27;
		17800: rom = 27;
		17801: rom = 27;
		17802: rom = 27;
		17803: rom = 27;
		17804: rom = 27;
		17805: rom = 27;
		17806: rom = 27;
		17807: rom = 27;
		17808: rom = 27;
		17809: rom = 27;
		17810: rom = 27;
		17811: rom = 27;
		17812: rom = 27;
		17813: rom = 27;
		17814: rom = 27;
		17815: rom = 27;
		17816: rom = 27;
		17817: rom = 27;
		17818: rom = 27;
		17819: rom = 27;
		17820: rom = 27;
		17821: rom = 27;
		17822: rom = 27;
		17823: rom = 27;
		17824: rom = 23;
		17825: rom = 15;
		17826: rom = 18;
		17827: rom = 18;
		17828: rom = 18;
		17829: rom = 18;
		17830: rom = 18;
		17831: rom = 15;
		17832: rom = 27;
		17833: rom = 27;
		17834: rom = 27;
		17835: rom = 27;
		17836: rom = 27;
		17837: rom = 27;
		17838: rom = 27;
		17839: rom = 27;
		17840: rom = 27;
		17841: rom = 27;
		17842: rom = 27;
		17843: rom = 27;
		17844: rom = 27;
		17845: rom = 27;
		17846: rom = 27;
		17847: rom = 27;
		17848: rom = 27;
		17849: rom = 27;
		17850: rom = 27;
		17851: rom = 26;
		17852: rom = 15;
		17853: rom = 14;
		17854: rom = 18;
		17855: rom = 18;
		17856: rom = 18;
		17857: rom = 18;
		17858: rom = 18;
		17859: rom = 18;
		17860: rom = 18;
		17861: rom = 18;
		17862: rom = 18;
		17863: rom = 18;
		17864: rom = 18;
		17865: rom = 18;
		17866: rom = 18;
		17867: rom = 18;
		17868: rom = 18;
		17869: rom = 18;
		17870: rom = 18;
		17871: rom = 18;
		17872: rom = 18;
		17873: rom = 18;
		17874: rom = 18;
		17875: rom = 18;
		17876: rom = 18;
		17877: rom = 18;
		17878: rom = 18;
		17879: rom = 18;
		17880: rom = 18;
		17881: rom = 18;
		17882: rom = 18;
		17883: rom = 18;
		17884: rom = 18;
		17885: rom = 18;
		17886: rom = 18;
		17887: rom = 18;
		17888: rom = 18;
		17889: rom = 18;
		17890: rom = 18;
		17891: rom = 18;
		17892: rom = 18;
		17893: rom = 17;
		17894: rom = 11;
		17895: rom = 26;
		17896: rom = 27;
		17897: rom = 27;
		17898: rom = 27;
		17899: rom = 27;
		17900: rom = 27;
		17901: rom = 27;
		17902: rom = 27;
		17903: rom = 27;
		17904: rom = 19;
		17905: rom = 10;
		17906: rom = 20;
		17907: rom = 18;
		17908: rom = 11;
		17909: rom = 19;
		17910: rom = 27;
		17911: rom = 27;
		17912: rom = 27;
		17913: rom = 27;
		17914: rom = 27;
		17920: rom = 27;
		17921: rom = 27;
		17922: rom = 27;
		17923: rom = 27;
		17924: rom = 27;
		17925: rom = 27;
		17926: rom = 27;
		17927: rom = 27;
		17928: rom = 27;
		17929: rom = 27;
		17930: rom = 27;
		17931: rom = 27;
		17932: rom = 27;
		17933: rom = 27;
		17934: rom = 27;
		17935: rom = 27;
		17936: rom = 27;
		17937: rom = 27;
		17938: rom = 27;
		17939: rom = 27;
		17940: rom = 27;
		17941: rom = 27;
		17942: rom = 27;
		17943: rom = 27;
		17944: rom = 27;
		17945: rom = 27;
		17946: rom = 27;
		17947: rom = 27;
		17948: rom = 27;
		17949: rom = 27;
		17950: rom = 27;
		17951: rom = 27;
		17952: rom = 23;
		17953: rom = 15;
		17954: rom = 18;
		17955: rom = 18;
		17956: rom = 18;
		17957: rom = 18;
		17958: rom = 18;
		17959: rom = 12;
		17960: rom = 27;
		17961: rom = 27;
		17962: rom = 27;
		17963: rom = 27;
		17964: rom = 27;
		17965: rom = 27;
		17966: rom = 27;
		17967: rom = 27;
		17968: rom = 27;
		17969: rom = 27;
		17970: rom = 27;
		17971: rom = 27;
		17972: rom = 27;
		17973: rom = 27;
		17974: rom = 27;
		17975: rom = 27;
		17976: rom = 27;
		17977: rom = 27;
		17978: rom = 27;
		17979: rom = 27;
		17980: rom = 27;
		17981: rom = 19;
		17982: rom = 12;
		17983: rom = 17;
		17984: rom = 18;
		17985: rom = 18;
		17986: rom = 18;
		17987: rom = 18;
		17988: rom = 18;
		17989: rom = 18;
		17990: rom = 18;
		17991: rom = 18;
		17992: rom = 18;
		17993: rom = 18;
		17994: rom = 18;
		17995: rom = 18;
		17996: rom = 18;
		17997: rom = 18;
		17998: rom = 18;
		17999: rom = 18;
		18000: rom = 18;
		18001: rom = 18;
		18002: rom = 18;
		18003: rom = 18;
		18004: rom = 18;
		18005: rom = 18;
		18006: rom = 18;
		18007: rom = 18;
		18008: rom = 18;
		18009: rom = 18;
		18010: rom = 18;
		18011: rom = 18;
		18012: rom = 18;
		18013: rom = 18;
		18014: rom = 18;
		18015: rom = 18;
		18016: rom = 18;
		18017: rom = 18;
		18018: rom = 18;
		18019: rom = 18;
		18020: rom = 17;
		18021: rom = 11;
		18022: rom = 24;
		18023: rom = 27;
		18024: rom = 27;
		18025: rom = 27;
		18026: rom = 27;
		18027: rom = 27;
		18028: rom = 27;
		18029: rom = 27;
		18030: rom = 27;
		18031: rom = 27;
		18032: rom = 27;
		18033: rom = 23;
		18034: rom = 14;
		18035: rom = 18;
		18036: rom = 25;
		18037: rom = 25;
		18038: rom = 22;
		18039: rom = 27;
		18040: rom = 27;
		18041: rom = 27;
		18042: rom = 27;
		18048: rom = 27;
		18049: rom = 27;
		18050: rom = 27;
		18051: rom = 27;
		18052: rom = 27;
		18053: rom = 27;
		18054: rom = 27;
		18055: rom = 27;
		18056: rom = 27;
		18057: rom = 27;
		18058: rom = 27;
		18059: rom = 27;
		18060: rom = 27;
		18061: rom = 27;
		18062: rom = 27;
		18063: rom = 27;
		18064: rom = 27;
		18065: rom = 27;
		18066: rom = 27;
		18067: rom = 27;
		18068: rom = 27;
		18069: rom = 27;
		18070: rom = 27;
		18071: rom = 27;
		18072: rom = 27;
		18073: rom = 27;
		18074: rom = 27;
		18075: rom = 27;
		18076: rom = 27;
		18077: rom = 27;
		18078: rom = 27;
		18079: rom = 27;
		18080: rom = 23;
		18081: rom = 14;
		18082: rom = 18;
		18083: rom = 18;
		18084: rom = 18;
		18085: rom = 18;
		18086: rom = 18;
		18087: rom = 14;
		18088: rom = 23;
		18089: rom = 27;
		18090: rom = 27;
		18091: rom = 27;
		18092: rom = 27;
		18093: rom = 27;
		18094: rom = 27;
		18095: rom = 27;
		18096: rom = 27;
		18097: rom = 27;
		18098: rom = 27;
		18099: rom = 27;
		18100: rom = 27;
		18101: rom = 27;
		18102: rom = 27;
		18103: rom = 27;
		18104: rom = 27;
		18105: rom = 27;
		18106: rom = 27;
		18107: rom = 27;
		18108: rom = 27;
		18109: rom = 27;
		18110: rom = 23;
		18111: rom = 11;
		18112: rom = 17;
		18113: rom = 18;
		18114: rom = 18;
		18115: rom = 18;
		18116: rom = 18;
		18117: rom = 18;
		18118: rom = 18;
		18119: rom = 18;
		18120: rom = 18;
		18121: rom = 18;
		18122: rom = 18;
		18123: rom = 18;
		18124: rom = 18;
		18125: rom = 18;
		18126: rom = 18;
		18127: rom = 18;
		18128: rom = 18;
		18129: rom = 18;
		18130: rom = 18;
		18131: rom = 18;
		18132: rom = 18;
		18133: rom = 18;
		18134: rom = 18;
		18135: rom = 18;
		18136: rom = 18;
		18137: rom = 18;
		18138: rom = 18;
		18139: rom = 18;
		18140: rom = 18;
		18141: rom = 18;
		18142: rom = 18;
		18143: rom = 18;
		18144: rom = 18;
		18145: rom = 18;
		18146: rom = 18;
		18147: rom = 18;
		18148: rom = 12;
		18149: rom = 22;
		18150: rom = 27;
		18151: rom = 27;
		18152: rom = 27;
		18153: rom = 27;
		18154: rom = 27;
		18155: rom = 27;
		18156: rom = 27;
		18157: rom = 27;
		18158: rom = 27;
		18159: rom = 27;
		18160: rom = 27;
		18161: rom = 27;
		18162: rom = 27;
		18163: rom = 27;
		18164: rom = 21;
		18165: rom = 0;
		18166: rom = 19;
		18167: rom = 27;
		18168: rom = 27;
		18169: rom = 27;
		18170: rom = 27;
		18176: rom = 27;
		18177: rom = 27;
		18178: rom = 27;
		18179: rom = 27;
		18180: rom = 27;
		18181: rom = 27;
		18182: rom = 27;
		18183: rom = 27;
		18184: rom = 27;
		18185: rom = 27;
		18186: rom = 27;
		18187: rom = 27;
		18188: rom = 27;
		18189: rom = 27;
		18190: rom = 27;
		18191: rom = 27;
		18192: rom = 27;
		18193: rom = 27;
		18194: rom = 27;
		18195: rom = 27;
		18196: rom = 27;
		18197: rom = 27;
		18198: rom = 27;
		18199: rom = 27;
		18200: rom = 27;
		18201: rom = 27;
		18202: rom = 27;
		18203: rom = 27;
		18204: rom = 27;
		18205: rom = 27;
		18206: rom = 27;
		18207: rom = 27;
		18208: rom = 24;
		18209: rom = 13;
		18210: rom = 18;
		18211: rom = 18;
		18212: rom = 18;
		18213: rom = 18;
		18214: rom = 18;
		18215: rom = 17;
		18216: rom = 14;
		18217: rom = 27;
		18218: rom = 27;
		18219: rom = 27;
		18220: rom = 27;
		18221: rom = 27;
		18222: rom = 27;
		18223: rom = 27;
		18224: rom = 27;
		18225: rom = 27;
		18226: rom = 27;
		18227: rom = 27;
		18228: rom = 27;
		18229: rom = 27;
		18230: rom = 27;
		18231: rom = 27;
		18232: rom = 27;
		18233: rom = 27;
		18234: rom = 27;
		18235: rom = 27;
		18236: rom = 27;
		18237: rom = 27;
		18238: rom = 27;
		18239: rom = 25;
		18240: rom = 12;
		18241: rom = 16;
		18242: rom = 18;
		18243: rom = 18;
		18244: rom = 18;
		18245: rom = 18;
		18246: rom = 18;
		18247: rom = 18;
		18248: rom = 18;
		18249: rom = 18;
		18250: rom = 18;
		18251: rom = 18;
		18252: rom = 18;
		18253: rom = 18;
		18254: rom = 18;
		18255: rom = 18;
		18256: rom = 18;
		18257: rom = 18;
		18258: rom = 18;
		18259: rom = 18;
		18260: rom = 18;
		18261: rom = 18;
		18262: rom = 18;
		18263: rom = 18;
		18264: rom = 18;
		18265: rom = 18;
		18266: rom = 18;
		18267: rom = 18;
		18268: rom = 18;
		18269: rom = 18;
		18270: rom = 18;
		18271: rom = 18;
		18272: rom = 18;
		18273: rom = 18;
		18274: rom = 18;
		18275: rom = 12;
		18276: rom = 21;
		18277: rom = 27;
		18278: rom = 27;
		18279: rom = 27;
		18280: rom = 27;
		18281: rom = 27;
		18282: rom = 27;
		18283: rom = 27;
		18284: rom = 27;
		18285: rom = 27;
		18286: rom = 27;
		18287: rom = 27;
		18288: rom = 27;
		18289: rom = 27;
		18290: rom = 26;
		18291: rom = 15;
		18292: rom = 0;
		18293: rom = 0;
		18294: rom = 19;
		18295: rom = 27;
		18296: rom = 27;
		18297: rom = 27;
		18298: rom = 27;
		18304: rom = 27;
		18305: rom = 27;
		18306: rom = 27;
		18307: rom = 27;
		18308: rom = 27;
		18309: rom = 27;
		18310: rom = 27;
		18311: rom = 27;
		18312: rom = 27;
		18313: rom = 27;
		18314: rom = 27;
		18315: rom = 27;
		18316: rom = 27;
		18317: rom = 27;
		18318: rom = 27;
		18319: rom = 27;
		18320: rom = 27;
		18321: rom = 27;
		18322: rom = 27;
		18323: rom = 27;
		18324: rom = 27;
		18325: rom = 27;
		18326: rom = 27;
		18327: rom = 27;
		18328: rom = 27;
		18329: rom = 27;
		18330: rom = 27;
		18331: rom = 27;
		18332: rom = 27;
		18333: rom = 27;
		18334: rom = 27;
		18335: rom = 27;
		18336: rom = 26;
		18337: rom = 12;
		18338: rom = 18;
		18339: rom = 18;
		18340: rom = 18;
		18341: rom = 18;
		18342: rom = 18;
		18343: rom = 18;
		18344: rom = 14;
		18345: rom = 21;
		18346: rom = 27;
		18347: rom = 27;
		18348: rom = 27;
		18349: rom = 27;
		18350: rom = 27;
		18351: rom = 27;
		18352: rom = 27;
		18353: rom = 27;
		18354: rom = 27;
		18355: rom = 27;
		18356: rom = 27;
		18357: rom = 27;
		18358: rom = 27;
		18359: rom = 27;
		18360: rom = 27;
		18361: rom = 27;
		18362: rom = 27;
		18363: rom = 27;
		18364: rom = 27;
		18365: rom = 27;
		18366: rom = 27;
		18367: rom = 27;
		18368: rom = 26;
		18369: rom = 15;
		18370: rom = 15;
		18371: rom = 18;
		18372: rom = 18;
		18373: rom = 18;
		18374: rom = 18;
		18375: rom = 18;
		18376: rom = 18;
		18377: rom = 18;
		18378: rom = 18;
		18379: rom = 18;
		18380: rom = 18;
		18381: rom = 18;
		18382: rom = 18;
		18383: rom = 18;
		18384: rom = 18;
		18385: rom = 18;
		18386: rom = 18;
		18387: rom = 18;
		18388: rom = 18;
		18389: rom = 18;
		18390: rom = 18;
		18391: rom = 18;
		18392: rom = 18;
		18393: rom = 18;
		18394: rom = 18;
		18395: rom = 18;
		18396: rom = 18;
		18397: rom = 18;
		18398: rom = 18;
		18399: rom = 18;
		18400: rom = 18;
		18401: rom = 17;
		18402: rom = 11;
		18403: rom = 22;
		18404: rom = 27;
		18405: rom = 27;
		18406: rom = 27;
		18407: rom = 27;
		18408: rom = 27;
		18409: rom = 27;
		18410: rom = 27;
		18411: rom = 27;
		18412: rom = 27;
		18413: rom = 27;
		18414: rom = 27;
		18415: rom = 27;
		18416: rom = 27;
		18417: rom = 23;
		18418: rom = 8;
		18419: rom = 0;
		18420: rom = 0;
		18421: rom = 0;
		18422: rom = 19;
		18423: rom = 27;
		18424: rom = 27;
		18425: rom = 27;
		18426: rom = 27;
		18432: rom = 27;
		18433: rom = 27;
		18434: rom = 27;
		18435: rom = 27;
		18436: rom = 27;
		18437: rom = 27;
		18438: rom = 27;
		18439: rom = 27;
		18440: rom = 27;
		18441: rom = 27;
		18442: rom = 27;
		18443: rom = 27;
		18444: rom = 27;
		18445: rom = 27;
		18446: rom = 27;
		18447: rom = 27;
		18448: rom = 27;
		18449: rom = 27;
		18450: rom = 27;
		18451: rom = 27;
		18452: rom = 27;
		18453: rom = 27;
		18454: rom = 27;
		18455: rom = 27;
		18456: rom = 27;
		18457: rom = 27;
		18458: rom = 27;
		18459: rom = 27;
		18460: rom = 27;
		18461: rom = 27;
		18462: rom = 27;
		18463: rom = 27;
		18464: rom = 27;
		18465: rom = 11;
		18466: rom = 18;
		18467: rom = 18;
		18468: rom = 18;
		18469: rom = 18;
		18470: rom = 18;
		18471: rom = 18;
		18472: rom = 18;
		18473: rom = 12;
		18474: rom = 22;
		18475: rom = 27;
		18476: rom = 27;
		18477: rom = 27;
		18478: rom = 27;
		18479: rom = 27;
		18480: rom = 27;
		18481: rom = 27;
		18482: rom = 27;
		18483: rom = 27;
		18484: rom = 27;
		18485: rom = 27;
		18486: rom = 27;
		18487: rom = 27;
		18488: rom = 27;
		18489: rom = 27;
		18490: rom = 27;
		18491: rom = 27;
		18492: rom = 27;
		18493: rom = 27;
		18494: rom = 27;
		18495: rom = 27;
		18496: rom = 27;
		18497: rom = 27;
		18498: rom = 17;
		18499: rom = 13;
		18500: rom = 18;
		18501: rom = 18;
		18502: rom = 18;
		18503: rom = 18;
		18504: rom = 18;
		18505: rom = 18;
		18506: rom = 18;
		18507: rom = 18;
		18508: rom = 18;
		18509: rom = 18;
		18510: rom = 18;
		18511: rom = 18;
		18512: rom = 18;
		18513: rom = 18;
		18514: rom = 18;
		18515: rom = 18;
		18516: rom = 18;
		18517: rom = 18;
		18518: rom = 18;
		18519: rom = 18;
		18520: rom = 18;
		18521: rom = 18;
		18522: rom = 18;
		18523: rom = 18;
		18524: rom = 18;
		18525: rom = 18;
		18526: rom = 18;
		18527: rom = 18;
		18528: rom = 16;
		18529: rom = 11;
		18530: rom = 24;
		18531: rom = 27;
		18532: rom = 27;
		18533: rom = 27;
		18534: rom = 27;
		18535: rom = 27;
		18536: rom = 27;
		18537: rom = 27;
		18538: rom = 27;
		18539: rom = 22;
		18540: rom = 21;
		18541: rom = 20;
		18542: rom = 27;
		18543: rom = 27;
		18544: rom = 17;
		18545: rom = 0;
		18546: rom = 0;
		18547: rom = 0;
		18548: rom = 0;
		18549: rom = 0;
		18550: rom = 19;
		18551: rom = 27;
		18552: rom = 27;
		18553: rom = 27;
		18554: rom = 27;
		18560: rom = 27;
		18561: rom = 27;
		18562: rom = 27;
		18563: rom = 27;
		18564: rom = 27;
		18565: rom = 27;
		18566: rom = 27;
		18567: rom = 27;
		18568: rom = 27;
		18569: rom = 27;
		18570: rom = 27;
		18571: rom = 27;
		18572: rom = 27;
		18573: rom = 27;
		18574: rom = 27;
		18575: rom = 27;
		18576: rom = 27;
		18577: rom = 27;
		18578: rom = 27;
		18579: rom = 27;
		18580: rom = 27;
		18581: rom = 27;
		18582: rom = 27;
		18583: rom = 27;
		18584: rom = 27;
		18585: rom = 27;
		18586: rom = 27;
		18587: rom = 27;
		18588: rom = 27;
		18589: rom = 27;
		18590: rom = 27;
		18591: rom = 27;
		18592: rom = 27;
		18593: rom = 14;
		18594: rom = 18;
		18595: rom = 18;
		18596: rom = 18;
		18597: rom = 18;
		18598: rom = 18;
		18599: rom = 18;
		18600: rom = 18;
		18601: rom = 18;
		18602: rom = 13;
		18603: rom = 16;
		18604: rom = 26;
		18605: rom = 27;
		18606: rom = 27;
		18607: rom = 27;
		18608: rom = 27;
		18609: rom = 27;
		18610: rom = 27;
		18611: rom = 27;
		18612: rom = 27;
		18613: rom = 27;
		18614: rom = 27;
		18615: rom = 27;
		18616: rom = 27;
		18617: rom = 27;
		18618: rom = 27;
		18619: rom = 27;
		18620: rom = 27;
		18621: rom = 27;
		18622: rom = 27;
		18623: rom = 27;
		18624: rom = 27;
		18625: rom = 27;
		18626: rom = 27;
		18627: rom = 20;
		18628: rom = 11;
		18629: rom = 17;
		18630: rom = 18;
		18631: rom = 18;
		18632: rom = 18;
		18633: rom = 18;
		18634: rom = 18;
		18635: rom = 18;
		18636: rom = 18;
		18637: rom = 18;
		18638: rom = 18;
		18639: rom = 18;
		18640: rom = 18;
		18641: rom = 18;
		18642: rom = 18;
		18643: rom = 18;
		18644: rom = 18;
		18645: rom = 18;
		18646: rom = 18;
		18647: rom = 18;
		18648: rom = 18;
		18649: rom = 18;
		18650: rom = 18;
		18651: rom = 18;
		18652: rom = 18;
		18653: rom = 18;
		18654: rom = 18;
		18655: rom = 14;
		18656: rom = 14;
		18657: rom = 26;
		18658: rom = 27;
		18659: rom = 27;
		18660: rom = 27;
		18661: rom = 27;
		18662: rom = 25;
		18663: rom = 22;
		18664: rom = 19;
		18665: rom = 8;
		18666: rom = 0;
		18667: rom = 0;
		18668: rom = 0;
		18669: rom = 27;
		18670: rom = 27;
		18671: rom = 10;
		18672: rom = 0;
		18673: rom = 0;
		18674: rom = 0;
		18675: rom = 19;
		18676: rom = 12;
		18677: rom = 0;
		18678: rom = 19;
		18679: rom = 27;
		18680: rom = 27;
		18681: rom = 27;
		18682: rom = 27;
		18688: rom = 27;
		18689: rom = 27;
		18690: rom = 27;
		18691: rom = 27;
		18692: rom = 27;
		18693: rom = 27;
		18694: rom = 27;
		18695: rom = 27;
		18696: rom = 27;
		18697: rom = 27;
		18698: rom = 27;
		18699: rom = 27;
		18700: rom = 27;
		18701: rom = 27;
		18702: rom = 27;
		18703: rom = 27;
		18704: rom = 27;
		18705: rom = 27;
		18706: rom = 27;
		18707: rom = 27;
		18708: rom = 27;
		18709: rom = 27;
		18710: rom = 27;
		18711: rom = 27;
		18712: rom = 27;
		18713: rom = 27;
		18714: rom = 27;
		18715: rom = 27;
		18716: rom = 27;
		18717: rom = 27;
		18718: rom = 27;
		18719: rom = 27;
		18720: rom = 27;
		18721: rom = 18;
		18722: rom = 17;
		18723: rom = 18;
		18724: rom = 18;
		18725: rom = 18;
		18726: rom = 18;
		18727: rom = 18;
		18728: rom = 18;
		18729: rom = 18;
		18730: rom = 18;
		18731: rom = 16;
		18732: rom = 11;
		18733: rom = 16;
		18734: rom = 22;
		18735: rom = 27;
		18736: rom = 27;
		18737: rom = 27;
		18738: rom = 27;
		18739: rom = 27;
		18740: rom = 27;
		18741: rom = 27;
		18742: rom = 27;
		18743: rom = 27;
		18744: rom = 27;
		18745: rom = 27;
		18746: rom = 27;
		18747: rom = 27;
		18748: rom = 27;
		18749: rom = 27;
		18750: rom = 27;
		18751: rom = 27;
		18752: rom = 27;
		18753: rom = 27;
		18754: rom = 27;
		18755: rom = 27;
		18756: rom = 24;
		18757: rom = 11;
		18758: rom = 15;
		18759: rom = 18;
		18760: rom = 18;
		18761: rom = 18;
		18762: rom = 18;
		18763: rom = 18;
		18764: rom = 18;
		18765: rom = 18;
		18766: rom = 18;
		18767: rom = 18;
		18768: rom = 18;
		18769: rom = 18;
		18770: rom = 18;
		18771: rom = 18;
		18772: rom = 18;
		18773: rom = 18;
		18774: rom = 18;
		18775: rom = 18;
		18776: rom = 18;
		18777: rom = 18;
		18778: rom = 18;
		18779: rom = 18;
		18780: rom = 18;
		18781: rom = 16;
		18782: rom = 11;
		18783: rom = 20;
		18784: rom = 27;
		18785: rom = 27;
		18786: rom = 27;
		18787: rom = 27;
		18788: rom = 27;
		18789: rom = 21;
		18790: rom = 18;
		18791: rom = 0;
		18792: rom = 0;
		18793: rom = 0;
		18794: rom = 0;
		18795: rom = 0;
		18796: rom = 27;
		18797: rom = 27;
		18798: rom = 0;
		18799: rom = 0;
		18800: rom = 0;
		18801: rom = 27;
		18802: rom = 27;
		18803: rom = 27;
		18804: rom = 27;
		18805: rom = 0;
		18806: rom = 19;
		18807: rom = 27;
		18808: rom = 27;
		18809: rom = 27;
		18810: rom = 27;
		18816: rom = 27;
		18817: rom = 27;
		18818: rom = 27;
		18819: rom = 27;
		18820: rom = 27;
		18821: rom = 27;
		18822: rom = 27;
		18823: rom = 27;
		18824: rom = 27;
		18825: rom = 27;
		18826: rom = 27;
		18827: rom = 27;
		18828: rom = 27;
		18829: rom = 27;
		18830: rom = 27;
		18831: rom = 27;
		18832: rom = 27;
		18833: rom = 27;
		18834: rom = 27;
		18835: rom = 27;
		18836: rom = 27;
		18837: rom = 27;
		18838: rom = 27;
		18839: rom = 27;
		18840: rom = 27;
		18841: rom = 27;
		18842: rom = 27;
		18843: rom = 27;
		18844: rom = 27;
		18845: rom = 27;
		18846: rom = 27;
		18847: rom = 27;
		18848: rom = 27;
		18849: rom = 22;
		18850: rom = 15;
		18851: rom = 18;
		18852: rom = 18;
		18853: rom = 18;
		18854: rom = 18;
		18855: rom = 18;
		18856: rom = 18;
		18857: rom = 18;
		18858: rom = 18;
		18859: rom = 18;
		18860: rom = 18;
		18861: rom = 17;
		18862: rom = 14;
		18863: rom = 10;
		18864: rom = 15;
		18865: rom = 21;
		18866: rom = 26;
		18867: rom = 27;
		18868: rom = 27;
		18869: rom = 27;
		18870: rom = 27;
		18871: rom = 27;
		18872: rom = 27;
		18873: rom = 27;
		18874: rom = 27;
		18875: rom = 27;
		18876: rom = 27;
		18877: rom = 27;
		18878: rom = 27;
		18879: rom = 27;
		18880: rom = 27;
		18881: rom = 27;
		18882: rom = 27;
		18883: rom = 27;
		18884: rom = 27;
		18885: rom = 26;
		18886: rom = 18;
		18887: rom = 11;
		18888: rom = 17;
		18889: rom = 18;
		18890: rom = 18;
		18891: rom = 18;
		18892: rom = 18;
		18893: rom = 18;
		18894: rom = 18;
		18895: rom = 18;
		18896: rom = 18;
		18897: rom = 18;
		18898: rom = 18;
		18899: rom = 18;
		18900: rom = 18;
		18901: rom = 18;
		18902: rom = 18;
		18903: rom = 18;
		18904: rom = 18;
		18905: rom = 18;
		18906: rom = 18;
		18907: rom = 17;
		18908: rom = 12;
		18909: rom = 16;
		18910: rom = 26;
		18911: rom = 27;
		18912: rom = 27;
		18913: rom = 27;
		18914: rom = 27;
		18915: rom = 27;
		18916: rom = 27;
		18917: rom = 13;
		18918: rom = 0;
		18919: rom = 0;
		18920: rom = 0;
		18921: rom = 0;
		18922: rom = 27;
		18923: rom = 27;
		18924: rom = 27;
		18925: rom = 0;
		18926: rom = 0;
		18927: rom = 0;
		18928: rom = 27;
		18929: rom = 27;
		18930: rom = 2;
		18931: rom = 0;
		18932: rom = 27;
		18933: rom = 27;
		18934: rom = 27;
		18935: rom = 27;
		18936: rom = 27;
		18937: rom = 27;
		18938: rom = 27;
		18944: rom = 27;
		18945: rom = 27;
		18946: rom = 27;
		18947: rom = 27;
		18948: rom = 27;
		18949: rom = 27;
		18950: rom = 27;
		18951: rom = 27;
		18952: rom = 27;
		18953: rom = 27;
		18954: rom = 27;
		18955: rom = 27;
		18956: rom = 27;
		18957: rom = 27;
		18958: rom = 27;
		18959: rom = 27;
		18960: rom = 27;
		18961: rom = 27;
		18962: rom = 27;
		18963: rom = 27;
		18964: rom = 27;
		18965: rom = 27;
		18966: rom = 27;
		18967: rom = 27;
		18968: rom = 27;
		18969: rom = 27;
		18970: rom = 27;
		18971: rom = 27;
		18972: rom = 27;
		18973: rom = 27;
		18974: rom = 27;
		18975: rom = 27;
		18976: rom = 27;
		18977: rom = 26;
		18978: rom = 11;
		18979: rom = 18;
		18980: rom = 18;
		18981: rom = 18;
		18982: rom = 18;
		18983: rom = 18;
		18984: rom = 18;
		18985: rom = 18;
		18986: rom = 18;
		18987: rom = 18;
		18988: rom = 18;
		18989: rom = 18;
		18990: rom = 18;
		18991: rom = 18;
		18992: rom = 17;
		18993: rom = 14;
		18994: rom = 11;
		18995: rom = 15;
		18996: rom = 22;
		18997: rom = 27;
		18998: rom = 27;
		18999: rom = 27;
		19000: rom = 27;
		19001: rom = 27;
		19002: rom = 27;
		19003: rom = 27;
		19004: rom = 27;
		19005: rom = 27;
		19006: rom = 27;
		19007: rom = 27;
		19008: rom = 27;
		19009: rom = 27;
		19010: rom = 27;
		19011: rom = 27;
		19012: rom = 27;
		19013: rom = 27;
		19014: rom = 27;
		19015: rom = 24;
		19016: rom = 14;
		19017: rom = 12;
		19018: rom = 17;
		19019: rom = 18;
		19020: rom = 18;
		19021: rom = 18;
		19022: rom = 18;
		19023: rom = 18;
		19024: rom = 18;
		19025: rom = 18;
		19026: rom = 18;
		19027: rom = 18;
		19028: rom = 18;
		19029: rom = 18;
		19030: rom = 18;
		19031: rom = 18;
		19032: rom = 18;
		19033: rom = 17;
		19034: rom = 12;
		19035: rom = 14;
		19036: rom = 24;
		19037: rom = 27;
		19038: rom = 27;
		19039: rom = 27;
		19040: rom = 27;
		19041: rom = 27;
		19042: rom = 27;
		19043: rom = 26;
		19044: rom = 11;
		19045: rom = 0;
		19046: rom = 0;
		19047: rom = 4;
		19048: rom = 27;
		19049: rom = 27;
		19050: rom = 27;
		19051: rom = 3;
		19052: rom = 0;
		19053: rom = 0;
		19054: rom = 9;
		19055: rom = 23;
		19056: rom = 27;
		19057: rom = 20;
		19058: rom = 6;
		19059: rom = 0;
		19060: rom = 0;
		19061: rom = 10;
		19062: rom = 24;
		19063: rom = 27;
		19064: rom = 27;
		19065: rom = 27;
		19066: rom = 27;
		19072: rom = 27;
		19073: rom = 27;
		19074: rom = 27;
		19075: rom = 27;
		19076: rom = 27;
		19077: rom = 27;
		19078: rom = 27;
		19079: rom = 27;
		19080: rom = 27;
		19081: rom = 27;
		19082: rom = 27;
		19083: rom = 27;
		19084: rom = 27;
		19085: rom = 27;
		19086: rom = 27;
		19087: rom = 27;
		19088: rom = 27;
		19089: rom = 27;
		19090: rom = 27;
		19091: rom = 27;
		19092: rom = 27;
		19093: rom = 27;
		19094: rom = 27;
		19095: rom = 27;
		19096: rom = 27;
		19097: rom = 27;
		19098: rom = 27;
		19099: rom = 27;
		19100: rom = 27;
		19101: rom = 27;
		19102: rom = 27;
		19103: rom = 27;
		19104: rom = 27;
		19105: rom = 27;
		19106: rom = 16;
		19107: rom = 17;
		19108: rom = 18;
		19109: rom = 18;
		19110: rom = 18;
		19111: rom = 18;
		19112: rom = 18;
		19113: rom = 18;
		19114: rom = 18;
		19115: rom = 18;
		19116: rom = 18;
		19117: rom = 18;
		19118: rom = 18;
		19119: rom = 18;
		19120: rom = 18;
		19121: rom = 18;
		19122: rom = 18;
		19123: rom = 17;
		19124: rom = 14;
		19125: rom = 10;
		19126: rom = 18;
		19127: rom = 25;
		19128: rom = 27;
		19129: rom = 27;
		19130: rom = 27;
		19131: rom = 27;
		19132: rom = 27;
		19133: rom = 27;
		19134: rom = 27;
		19135: rom = 27;
		19136: rom = 27;
		19137: rom = 27;
		19138: rom = 27;
		19139: rom = 27;
		19140: rom = 27;
		19141: rom = 27;
		19142: rom = 27;
		19143: rom = 27;
		19144: rom = 27;
		19145: rom = 24;
		19146: rom = 16;
		19147: rom = 11;
		19148: rom = 15;
		19149: rom = 17;
		19150: rom = 18;
		19151: rom = 18;
		19152: rom = 18;
		19153: rom = 18;
		19154: rom = 18;
		19155: rom = 18;
		19156: rom = 18;
		19157: rom = 18;
		19158: rom = 18;
		19159: rom = 15;
		19160: rom = 11;
		19161: rom = 15;
		19162: rom = 24;
		19163: rom = 27;
		19164: rom = 27;
		19165: rom = 27;
		19166: rom = 27;
		19167: rom = 27;
		19168: rom = 27;
		19169: rom = 27;
		19170: rom = 27;
		19171: rom = 13;
		19172: rom = 0;
		19173: rom = 0;
		19174: rom = 11;
		19175: rom = 27;
		19176: rom = 27;
		19177: rom = 13;
		19178: rom = 0;
		19179: rom = 0;
		19180: rom = 0;
		19181: rom = 17;
		19182: rom = 26;
		19183: rom = 27;
		19184: rom = 27;
		19185: rom = 27;
		19186: rom = 25;
		19187: rom = 12;
		19188: rom = 0;
		19189: rom = 0;
		19190: rom = 13;
		19191: rom = 27;
		19192: rom = 27;
		19193: rom = 27;
		19194: rom = 27;
		19200: rom = 27;
		19201: rom = 27;
		19202: rom = 27;
		19203: rom = 27;
		19204: rom = 27;
		19205: rom = 27;
		19206: rom = 27;
		19207: rom = 27;
		19208: rom = 27;
		19209: rom = 27;
		19210: rom = 27;
		19211: rom = 27;
		19212: rom = 27;
		19213: rom = 27;
		19214: rom = 27;
		19215: rom = 27;
		19216: rom = 27;
		19217: rom = 27;
		19218: rom = 27;
		19219: rom = 26;
		19220: rom = 18;
		19221: rom = 10;
		19222: rom = 0;
		19223: rom = 0;
		19224: rom = 11;
		19225: rom = 19;
		19226: rom = 26;
		19227: rom = 27;
		19228: rom = 27;
		19229: rom = 27;
		19230: rom = 27;
		19231: rom = 27;
		19232: rom = 27;
		19233: rom = 27;
		19234: rom = 22;
		19235: rom = 14;
		19236: rom = 18;
		19237: rom = 18;
		19238: rom = 18;
		19239: rom = 18;
		19240: rom = 18;
		19241: rom = 18;
		19242: rom = 18;
		19243: rom = 18;
		19244: rom = 18;
		19245: rom = 18;
		19246: rom = 18;
		19247: rom = 18;
		19248: rom = 18;
		19249: rom = 18;
		19250: rom = 18;
		19251: rom = 18;
		19252: rom = 18;
		19253: rom = 18;
		19254: rom = 16;
		19255: rom = 10;
		19256: rom = 16;
		19257: rom = 25;
		19258: rom = 27;
		19259: rom = 27;
		19260: rom = 21;
		19261: rom = 27;
		19262: rom = 27;
		19263: rom = 27;
		19264: rom = 27;
		19265: rom = 27;
		19266: rom = 27;
		19267: rom = 27;
		19268: rom = 27;
		19269: rom = 27;
		19270: rom = 27;
		19271: rom = 27;
		19272: rom = 27;
		19273: rom = 27;
		19274: rom = 27;
		19275: rom = 26;
		19276: rom = 21;
		19277: rom = 14;
		19278: rom = 10;
		19279: rom = 12;
		19280: rom = 13;
		19281: rom = 14;
		19282: rom = 15;
		19283: rom = 14;
		19284: rom = 13;
		19285: rom = 11;
		19286: rom = 11;
		19287: rom = 19;
		19288: rom = 25;
		19289: rom = 27;
		19290: rom = 27;
		19291: rom = 27;
		19292: rom = 27;
		19293: rom = 27;
		19294: rom = 27;
		19295: rom = 27;
		19296: rom = 27;
		19297: rom = 27;
		19298: rom = 20;
		19299: rom = 0;
		19300: rom = 0;
		19301: rom = 12;
		19302: rom = 27;
		19303: rom = 27;
		19304: rom = 5;
		19305: rom = 0;
		19306: rom = 0;
		19307: rom = 7;
		19308: rom = 22;
		19309: rom = 27;
		19310: rom = 27;
		19311: rom = 27;
		19312: rom = 27;
		19313: rom = 27;
		19314: rom = 27;
		19315: rom = 27;
		19316: rom = 13;
		19317: rom = 0;
		19318: rom = 0;
		19319: rom = 19;
		19320: rom = 27;
		19321: rom = 27;
		19322: rom = 27;
		19328: rom = 27;
		19329: rom = 27;
		19330: rom = 27;
		19331: rom = 27;
		19332: rom = 27;
		19333: rom = 27;
		19334: rom = 27;
		19335: rom = 27;
		19336: rom = 27;
		19337: rom = 27;
		19338: rom = 27;
		19339: rom = 27;
		19340: rom = 27;
		19341: rom = 27;
		19342: rom = 27;
		19343: rom = 27;
		19344: rom = 27;
		19345: rom = 27;
		19346: rom = 22;
		19347: rom = 6;
		19348: rom = 0;
		19349: rom = 0;
		19350: rom = 0;
		19351: rom = 0;
		19352: rom = 0;
		19353: rom = 0;
		19354: rom = 7;
		19355: rom = 24;
		19356: rom = 27;
		19357: rom = 27;
		19358: rom = 27;
		19359: rom = 27;
		19360: rom = 27;
		19361: rom = 27;
		19362: rom = 27;
		19363: rom = 12;
		19364: rom = 18;
		19365: rom = 18;
		19366: rom = 18;
		19367: rom = 18;
		19368: rom = 18;
		19369: rom = 18;
		19370: rom = 18;
		19371: rom = 18;
		19372: rom = 18;
		19373: rom = 18;
		19374: rom = 18;
		19375: rom = 18;
		19376: rom = 18;
		19377: rom = 18;
		19378: rom = 18;
		19379: rom = 18;
		19380: rom = 18;
		19381: rom = 18;
		19382: rom = 18;
		19383: rom = 18;
		19384: rom = 16;
		19385: rom = 15;
		19386: rom = 27;
		19387: rom = 24;
		19388: rom = 10;
		19389: rom = 17;
		19390: rom = 27;
		19391: rom = 27;
		19392: rom = 27;
		19393: rom = 27;
		19394: rom = 27;
		19395: rom = 27;
		19396: rom = 27;
		19397: rom = 27;
		19398: rom = 27;
		19399: rom = 27;
		19400: rom = 27;
		19401: rom = 27;
		19402: rom = 27;
		19403: rom = 27;
		19404: rom = 27;
		19405: rom = 27;
		19406: rom = 27;
		19407: rom = 25;
		19408: rom = 24;
		19409: rom = 21;
		19410: rom = 21;
		19411: rom = 22;
		19412: rom = 24;
		19413: rom = 26;
		19414: rom = 27;
		19415: rom = 27;
		19416: rom = 27;
		19417: rom = 27;
		19418: rom = 27;
		19419: rom = 27;
		19420: rom = 27;
		19421: rom = 27;
		19422: rom = 27;
		19423: rom = 27;
		19424: rom = 27;
		19425: rom = 26;
		19426: rom = 4;
		19427: rom = 0;
		19428: rom = 8;
		19429: rom = 27;
		19430: rom = 27;
		19431: rom = 0;
		19432: rom = 0;
		19433: rom = 0;
		19434: rom = 15;
		19435: rom = 26;
		19436: rom = 27;
		19437: rom = 27;
		19438: rom = 27;
		19439: rom = 27;
		19440: rom = 27;
		19441: rom = 27;
		19442: rom = 27;
		19443: rom = 27;
		19444: rom = 27;
		19445: rom = 10;
		19446: rom = 0;
		19447: rom = 0;
		19448: rom = 25;
		19449: rom = 27;
		19450: rom = 27;
		19456: rom = 27;
		19457: rom = 27;
		19458: rom = 27;
		19459: rom = 27;
		19460: rom = 27;
		19461: rom = 27;
		19462: rom = 27;
		19463: rom = 27;
		19464: rom = 27;
		19465: rom = 27;
		19466: rom = 27;
		19467: rom = 27;
		19468: rom = 27;
		19469: rom = 27;
		19470: rom = 27;
		19471: rom = 27;
		19472: rom = 27;
		19473: rom = 21;
		19474: rom = 0;
		19475: rom = 0;
		19476: rom = 0;
		19477: rom = 0;
		19478: rom = 0;
		19479: rom = 0;
		19480: rom = 0;
		19481: rom = 0;
		19482: rom = 0;
		19483: rom = 0;
		19484: rom = 24;
		19485: rom = 27;
		19486: rom = 27;
		19487: rom = 27;
		19488: rom = 27;
		19489: rom = 27;
		19490: rom = 27;
		19491: rom = 20;
		19492: rom = 16;
		19493: rom = 18;
		19494: rom = 18;
		19495: rom = 18;
		19496: rom = 18;
		19497: rom = 18;
		19498: rom = 18;
		19499: rom = 18;
		19500: rom = 18;
		19501: rom = 18;
		19502: rom = 18;
		19503: rom = 18;
		19504: rom = 18;
		19505: rom = 18;
		19506: rom = 18;
		19507: rom = 18;
		19508: rom = 18;
		19509: rom = 18;
		19510: rom = 18;
		19511: rom = 18;
		19512: rom = 15;
		19513: rom = 22;
		19514: rom = 27;
		19515: rom = 14;
		19516: rom = 17;
		19517: rom = 13;
		19518: rom = 21;
		19519: rom = 27;
		19520: rom = 27;
		19521: rom = 27;
		19522: rom = 27;
		19523: rom = 27;
		19524: rom = 27;
		19525: rom = 27;
		19526: rom = 27;
		19527: rom = 27;
		19528: rom = 27;
		19529: rom = 27;
		19530: rom = 27;
		19531: rom = 27;
		19532: rom = 27;
		19533: rom = 27;
		19534: rom = 27;
		19535: rom = 27;
		19536: rom = 27;
		19537: rom = 27;
		19538: rom = 27;
		19539: rom = 27;
		19540: rom = 27;
		19541: rom = 27;
		19542: rom = 27;
		19543: rom = 27;
		19544: rom = 27;
		19545: rom = 27;
		19546: rom = 27;
		19547: rom = 27;
		19548: rom = 27;
		19549: rom = 27;
		19550: rom = 27;
		19551: rom = 27;
		19552: rom = 27;
		19553: rom = 18;
		19554: rom = 0;
		19555: rom = 0;
		19556: rom = 27;
		19557: rom = 27;
		19558: rom = 0;
		19559: rom = 0;
		19560: rom = 5;
		19561: rom = 21;
		19562: rom = 27;
		19563: rom = 27;
		19564: rom = 27;
		19565: rom = 27;
		19566: rom = 27;
		19567: rom = 27;
		19568: rom = 27;
		19569: rom = 27;
		19570: rom = 27;
		19571: rom = 27;
		19572: rom = 13;
		19573: rom = 27;
		19574: rom = 0;
		19575: rom = 0;
		19576: rom = 17;
		19577: rom = 27;
		19578: rom = 27;
		19584: rom = 27;
		19585: rom = 27;
		19586: rom = 27;
		19587: rom = 27;
		19588: rom = 27;
		19589: rom = 27;
		19590: rom = 27;
		19591: rom = 27;
		19592: rom = 27;
		19593: rom = 22;
		19594: rom = 13;
		19595: rom = 0;
		19596: rom = 0;
		19597: rom = 15;
		19598: rom = 24;
		19599: rom = 27;
		19600: rom = 23;
		19601: rom = 0;
		19602: rom = 0;
		19603: rom = 0;
		19604: rom = 10;
		19605: rom = 19;
		19606: rom = 22;
		19607: rom = 21;
		19608: rom = 15;
		19609: rom = 0;
		19610: rom = 0;
		19611: rom = 0;
		19612: rom = 10;
		19613: rom = 27;
		19614: rom = 27;
		19615: rom = 27;
		19616: rom = 27;
		19617: rom = 27;
		19618: rom = 27;
		19619: rom = 26;
		19620: rom = 11;
		19621: rom = 18;
		19622: rom = 18;
		19623: rom = 18;
		19624: rom = 18;
		19625: rom = 18;
		19626: rom = 18;
		19627: rom = 18;
		19628: rom = 18;
		19629: rom = 18;
		19630: rom = 18;
		19631: rom = 18;
		19632: rom = 18;
		19633: rom = 18;
		19634: rom = 18;
		19635: rom = 18;
		19636: rom = 18;
		19637: rom = 18;
		19638: rom = 18;
		19639: rom = 18;
		19640: rom = 12;
		19641: rom = 26;
		19642: rom = 23;
		19643: rom = 14;
		19644: rom = 18;
		19645: rom = 18;
		19646: rom = 11;
		19647: rom = 24;
		19648: rom = 27;
		19649: rom = 27;
		19650: rom = 27;
		19651: rom = 27;
		19652: rom = 27;
		19653: rom = 27;
		19654: rom = 27;
		19655: rom = 27;
		19656: rom = 27;
		19657: rom = 27;
		19658: rom = 27;
		19659: rom = 27;
		19660: rom = 27;
		19661: rom = 27;
		19662: rom = 27;
		19663: rom = 27;
		19664: rom = 27;
		19665: rom = 27;
		19666: rom = 27;
		19667: rom = 27;
		19668: rom = 27;
		19669: rom = 27;
		19670: rom = 27;
		19671: rom = 27;
		19672: rom = 27;
		19673: rom = 27;
		19674: rom = 27;
		19675: rom = 27;
		19676: rom = 27;
		19677: rom = 27;
		19678: rom = 27;
		19679: rom = 27;
		19680: rom = 27;
		19681: rom = 6;
		19682: rom = 0;
		19683: rom = 27;
		19684: rom = 27;
		19685: rom = 0;
		19686: rom = 0;
		19687: rom = 13;
		19688: rom = 25;
		19689: rom = 27;
		19690: rom = 27;
		19691: rom = 27;
		19692: rom = 27;
		19693: rom = 27;
		19694: rom = 27;
		19695: rom = 27;
		19696: rom = 27;
		19697: rom = 27;
		19698: rom = 27;
		19699: rom = 27;
		19700: rom = 13;
		19701: rom = 8;
		19702: rom = 27;
		19703: rom = 0;
		19704: rom = 0;
		19705: rom = 26;
		19706: rom = 27;
		19712: rom = 27;
		19713: rom = 27;
		19714: rom = 27;
		19715: rom = 27;
		19716: rom = 27;
		19717: rom = 27;
		19718: rom = 27;
		19719: rom = 27;
		19720: rom = 18;
		19721: rom = 0;
		19722: rom = 0;
		19723: rom = 0;
		19724: rom = 0;
		19725: rom = 0;
		19726: rom = 0;
		19727: rom = 18;
		19728: rom = 8;
		19729: rom = 0;
		19730: rom = 0;
		19731: rom = 19;
		19732: rom = 27;
		19733: rom = 27;
		19734: rom = 27;
		19735: rom = 27;
		19736: rom = 27;
		19737: rom = 23;
		19738: rom = 0;
		19739: rom = 0;
		19740: rom = 0;
		19741: rom = 20;
		19742: rom = 27;
		19743: rom = 27;
		19744: rom = 27;
		19745: rom = 27;
		19746: rom = 27;
		19747: rom = 27;
		19748: rom = 18;
		19749: rom = 16;
		19750: rom = 18;
		19751: rom = 18;
		19752: rom = 18;
		19753: rom = 18;
		19754: rom = 18;
		19755: rom = 18;
		19756: rom = 18;
		19757: rom = 18;
		19758: rom = 18;
		19759: rom = 18;
		19760: rom = 18;
		19761: rom = 18;
		19762: rom = 18;
		19763: rom = 18;
		19764: rom = 18;
		19765: rom = 18;
		19766: rom = 18;
		19767: rom = 18;
		19768: rom = 13;
		19769: rom = 27;
		19770: rom = 12;
		19771: rom = 17;
		19772: rom = 18;
		19773: rom = 18;
		19774: rom = 17;
		19775: rom = 12;
		19776: rom = 26;
		19777: rom = 27;
		19778: rom = 27;
		19779: rom = 27;
		19780: rom = 27;
		19781: rom = 27;
		19782: rom = 27;
		19783: rom = 27;
		19784: rom = 27;
		19785: rom = 27;
		19786: rom = 27;
		19787: rom = 27;
		19788: rom = 27;
		19789: rom = 27;
		19790: rom = 27;
		19791: rom = 27;
		19792: rom = 27;
		19793: rom = 27;
		19794: rom = 27;
		19795: rom = 27;
		19796: rom = 27;
		19797: rom = 27;
		19798: rom = 27;
		19799: rom = 27;
		19800: rom = 27;
		19801: rom = 27;
		19802: rom = 27;
		19803: rom = 27;
		19804: rom = 27;
		19805: rom = 27;
		19806: rom = 27;
		19807: rom = 27;
		19808: rom = 23;
		19809: rom = 0;
		19810: rom = 0;
		19811: rom = 27;
		19812: rom = 0;
		19813: rom = 0;
		19814: rom = 20;
		19815: rom = 27;
		19816: rom = 27;
		19817: rom = 27;
		19818: rom = 27;
		19819: rom = 27;
		19820: rom = 27;
		19821: rom = 27;
		19822: rom = 27;
		19823: rom = 27;
		19824: rom = 27;
		19825: rom = 27;
		19826: rom = 27;
		19827: rom = 27;
		19828: rom = 13;
		19829: rom = 0;
		19830: rom = 27;
		19831: rom = 0;
		19832: rom = 0;
		19833: rom = 22;
		19834: rom = 27;
		19840: rom = 27;
		19841: rom = 27;
		19842: rom = 27;
		19843: rom = 27;
		19844: rom = 27;
		19845: rom = 27;
		19846: rom = 27;
		19847: rom = 22;
		19848: rom = 0;
		19849: rom = 0;
		19850: rom = 0;
		19851: rom = 0;
		19852: rom = 0;
		19853: rom = 0;
		19854: rom = 0;
		19855: rom = 0;
		19856: rom = 0;
		19857: rom = 0;
		19858: rom = 21;
		19859: rom = 27;
		19860: rom = 27;
		19861: rom = 27;
		19862: rom = 27;
		19863: rom = 27;
		19864: rom = 27;
		19865: rom = 27;
		19866: rom = 22;
		19867: rom = 0;
		19868: rom = 0;
		19869: rom = 10;
		19870: rom = 27;
		19871: rom = 27;
		19872: rom = 27;
		19873: rom = 27;
		19874: rom = 27;
		19875: rom = 27;
		19876: rom = 25;
		19877: rom = 11;
		19878: rom = 18;
		19879: rom = 18;
		19880: rom = 18;
		19881: rom = 18;
		19882: rom = 18;
		19883: rom = 18;
		19884: rom = 18;
		19885: rom = 18;
		19886: rom = 18;
		19887: rom = 18;
		19888: rom = 18;
		19889: rom = 18;
		19890: rom = 18;
		19891: rom = 18;
		19892: rom = 18;
		19893: rom = 18;
		19894: rom = 18;
		19895: rom = 18;
		19896: rom = 16;
		19897: rom = 21;
		19898: rom = 15;
		19899: rom = 18;
		19900: rom = 18;
		19901: rom = 18;
		19902: rom = 18;
		19903: rom = 17;
		19904: rom = 13;
		19905: rom = 27;
		19906: rom = 27;
		19907: rom = 27;
		19908: rom = 27;
		19909: rom = 27;
		19910: rom = 27;
		19911: rom = 27;
		19912: rom = 27;
		19913: rom = 27;
		19914: rom = 27;
		19915: rom = 27;
		19916: rom = 27;
		19917: rom = 27;
		19918: rom = 27;
		19919: rom = 27;
		19920: rom = 27;
		19921: rom = 27;
		19922: rom = 27;
		19923: rom = 27;
		19924: rom = 27;
		19925: rom = 27;
		19926: rom = 27;
		19927: rom = 27;
		19928: rom = 27;
		19929: rom = 27;
		19930: rom = 27;
		19931: rom = 27;
		19932: rom = 27;
		19933: rom = 27;
		19934: rom = 27;
		19935: rom = 27;
		19936: rom = 18;
		19937: rom = 0;
		19938: rom = 0;
		19939: rom = 27;
		19940: rom = 12;
		19941: rom = 25;
		19942: rom = 27;
		19943: rom = 27;
		19944: rom = 27;
		19945: rom = 27;
		19946: rom = 27;
		19947: rom = 0;
		19948: rom = 0;
		19949: rom = 0;
		19950: rom = 0;
		19951: rom = 27;
		19952: rom = 27;
		19953: rom = 27;
		19954: rom = 27;
		19955: rom = 27;
		19956: rom = 13;
		19957: rom = 0;
		19958: rom = 27;
		19959: rom = 8;
		19960: rom = 0;
		19961: rom = 17;
		19962: rom = 27;
		19968: rom = 27;
		19969: rom = 27;
		19970: rom = 27;
		19971: rom = 27;
		19972: rom = 27;
		19973: rom = 27;
		19974: rom = 27;
		19975: rom = 10;
		19976: rom = 0;
		19977: rom = 0;
		19978: rom = 14;
		19979: rom = 22;
		19980: rom = 21;
		19981: rom = 12;
		19982: rom = 0;
		19983: rom = 0;
		19984: rom = 0;
		19985: rom = 14;
		19986: rom = 27;
		19987: rom = 27;
		19988: rom = 27;
		19989: rom = 27;
		19990: rom = 27;
		19991: rom = 27;
		19992: rom = 27;
		19993: rom = 27;
		19994: rom = 27;
		19995: rom = 14;
		19996: rom = 0;
		19997: rom = 0;
		19998: rom = 25;
		19999: rom = 27;
		20000: rom = 27;
		20001: rom = 27;
		20002: rom = 27;
		20003: rom = 27;
		20004: rom = 27;
		20005: rom = 16;
		20006: rom = 17;
		20007: rom = 18;
		20008: rom = 18;
		20009: rom = 18;
		20010: rom = 18;
		20011: rom = 18;
		20012: rom = 18;
		20013: rom = 18;
		20014: rom = 18;
		20015: rom = 18;
		20016: rom = 18;
		20017: rom = 18;
		20018: rom = 18;
		20019: rom = 18;
		20020: rom = 18;
		20021: rom = 18;
		20022: rom = 18;
		20023: rom = 16;
		20024: rom = 19;
		20025: rom = 12;
		20026: rom = 18;
		20027: rom = 18;
		20028: rom = 18;
		20029: rom = 18;
		20030: rom = 18;
		20031: rom = 18;
		20032: rom = 15;
		20033: rom = 17;
		20034: rom = 27;
		20035: rom = 27;
		20036: rom = 27;
		20037: rom = 27;
		20038: rom = 27;
		20039: rom = 27;
		20040: rom = 27;
		20041: rom = 27;
		20042: rom = 27;
		20043: rom = 27;
		20044: rom = 27;
		20045: rom = 27;
		20046: rom = 27;
		20047: rom = 27;
		20048: rom = 27;
		20049: rom = 27;
		20050: rom = 27;
		20051: rom = 27;
		20052: rom = 27;
		20053: rom = 27;
		20054: rom = 27;
		20055: rom = 27;
		20056: rom = 27;
		20057: rom = 27;
		20058: rom = 27;
		20059: rom = 27;
		20060: rom = 27;
		20061: rom = 27;
		20062: rom = 23;
		20063: rom = 27;
		20064: rom = 13;
		20065: rom = 0;
		20066: rom = 14;
		20067: rom = 27;
		20068: rom = 27;
		20069: rom = 27;
		20070: rom = 27;
		20071: rom = 27;
		20072: rom = 27;
		20073: rom = 27;
		20074: rom = 27;
		20075: rom = 27;
		20076: rom = 0;
		20077: rom = 0;
		20078: rom = 27;
		20079: rom = 27;
		20080: rom = 27;
		20081: rom = 27;
		20082: rom = 27;
		20083: rom = 27;
		20084: rom = 13;
		20085: rom = 0;
		20086: rom = 27;
		20087: rom = 16;
		20088: rom = 0;
		20089: rom = 11;
		20090: rom = 27;
		20096: rom = 27;
		20097: rom = 27;
		20098: rom = 27;
		20099: rom = 27;
		20100: rom = 27;
		20101: rom = 27;
		20102: rom = 24;
		20103: rom = 0;
		20104: rom = 0;
		20105: rom = 15;
		20106: rom = 27;
		20107: rom = 27;
		20108: rom = 27;
		20109: rom = 27;
		20110: rom = 17;
		20111: rom = 0;
		20112: rom = 0;
		20113: rom = 0;
		20114: rom = 21;
		20115: rom = 27;
		20116: rom = 27;
		20117: rom = 27;
		20118: rom = 27;
		20119: rom = 27;
		20120: rom = 27;
		20121: rom = 27;
		20122: rom = 27;
		20123: rom = 22;
		20124: rom = 0;
		20125: rom = 0;
		20126: rom = 23;
		20127: rom = 27;
		20128: rom = 27;
		20129: rom = 27;
		20130: rom = 27;
		20131: rom = 27;
		20132: rom = 27;
		20133: rom = 24;
		20134: rom = 13;
		20135: rom = 18;
		20136: rom = 18;
		20137: rom = 18;
		20138: rom = 18;
		20139: rom = 18;
		20140: rom = 18;
		20141: rom = 18;
		20142: rom = 18;
		20143: rom = 18;
		20144: rom = 18;
		20145: rom = 18;
		20146: rom = 18;
		20147: rom = 18;
		20148: rom = 18;
		20149: rom = 18;
		20150: rom = 18;
		20151: rom = 15;
		20152: rom = 10;
		20153: rom = 16;
		20154: rom = 18;
		20155: rom = 18;
		20156: rom = 18;
		20157: rom = 18;
		20158: rom = 18;
		20159: rom = 18;
		20160: rom = 23;
		20161: rom = 20;
		20162: rom = 21;
		20163: rom = 27;
		20164: rom = 27;
		20165: rom = 27;
		20166: rom = 27;
		20167: rom = 27;
		20168: rom = 27;
		20169: rom = 27;
		20170: rom = 27;
		20171: rom = 27;
		20172: rom = 27;
		20173: rom = 27;
		20174: rom = 27;
		20175: rom = 27;
		20176: rom = 27;
		20177: rom = 27;
		20178: rom = 27;
		20179: rom = 27;
		20180: rom = 27;
		20181: rom = 27;
		20182: rom = 27;
		20183: rom = 27;
		20184: rom = 27;
		20185: rom = 27;
		20186: rom = 27;
		20187: rom = 27;
		20188: rom = 27;
		20189: rom = 17;
		20190: rom = 0;
		20191: rom = 27;
		20192: rom = 0;
		20193: rom = 0;
		20194: rom = 19;
		20195: rom = 27;
		20196: rom = 27;
		20197: rom = 27;
		20198: rom = 27;
		20199: rom = 27;
		20200: rom = 27;
		20201: rom = 27;
		20202: rom = 27;
		20203: rom = 27;
		20204: rom = 0;
		20205: rom = 0;
		20206: rom = 27;
		20207: rom = 27;
		20208: rom = 27;
		20209: rom = 27;
		20210: rom = 27;
		20211: rom = 27;
		20212: rom = 13;
		20213: rom = 0;
		20214: rom = 27;
		20215: rom = 20;
		20216: rom = 0;
		20217: rom = 0;
		20218: rom = 27;
		20224: rom = 27;
		20225: rom = 27;
		20226: rom = 27;
		20227: rom = 27;
		20228: rom = 27;
		20229: rom = 27;
		20230: rom = 21;
		20231: rom = 0;
		20232: rom = 0;
		20233: rom = 25;
		20234: rom = 27;
		20235: rom = 27;
		20236: rom = 27;
		20237: rom = 27;
		20238: rom = 27;
		20239: rom = 17;
		20240: rom = 0;
		20241: rom = 0;
		20242: rom = 0;
		20243: rom = 22;
		20244: rom = 27;
		20245: rom = 27;
		20246: rom = 27;
		20247: rom = 27;
		20248: rom = 27;
		20249: rom = 27;
		20250: rom = 27;
		20251: rom = 25;
		20252: rom = 0;
		20253: rom = 0;
		20254: rom = 21;
		20255: rom = 27;
		20256: rom = 27;
		20257: rom = 27;
		20258: rom = 27;
		20259: rom = 27;
		20260: rom = 27;
		20261: rom = 27;
		20262: rom = 15;
		20263: rom = 17;
		20264: rom = 18;
		20265: rom = 18;
		20266: rom = 18;
		20267: rom = 18;
		20268: rom = 18;
		20269: rom = 18;
		20270: rom = 18;
		20271: rom = 18;
		20272: rom = 18;
		20273: rom = 18;
		20274: rom = 18;
		20275: rom = 18;
		20276: rom = 18;
		20277: rom = 18;
		20278: rom = 18;
		20279: rom = 14;
		20280: rom = 9;
		20281: rom = 18;
		20282: rom = 18;
		20283: rom = 18;
		20284: rom = 18;
		20285: rom = 18;
		20286: rom = 18;
		20287: rom = 23;
		20288: rom = 25;
		20289: rom = 24;
		20290: rom = 13;
		20291: rom = 23;
		20292: rom = 27;
		20293: rom = 27;
		20294: rom = 27;
		20295: rom = 27;
		20296: rom = 27;
		20297: rom = 27;
		20298: rom = 27;
		20299: rom = 27;
		20300: rom = 27;
		20301: rom = 27;
		20302: rom = 27;
		20303: rom = 27;
		20304: rom = 27;
		20305: rom = 27;
		20306: rom = 27;
		20307: rom = 27;
		20308: rom = 27;
		20309: rom = 27;
		20310: rom = 27;
		20311: rom = 27;
		20312: rom = 27;
		20313: rom = 27;
		20314: rom = 27;
		20315: rom = 24;
		20316: rom = 10;
		20317: rom = 0;
		20318: rom = 0;
		20319: rom = 27;
		20320: rom = 0;
		20321: rom = 0;
		20322: rom = 20;
		20323: rom = 27;
		20324: rom = 27;
		20325: rom = 27;
		20326: rom = 27;
		20327: rom = 27;
		20328: rom = 27;
		20329: rom = 27;
		20330: rom = 27;
		20331: rom = 27;
		20332: rom = 0;
		20333: rom = 0;
		20334: rom = 27;
		20335: rom = 27;
		20336: rom = 27;
		20337: rom = 27;
		20338: rom = 27;
		20339: rom = 27;
		20340: rom = 13;
		20341: rom = 0;
		20342: rom = 27;
		20343: rom = 21;
		20344: rom = 0;
		20345: rom = 0;
		20346: rom = 26;
		20352: rom = 27;
		20353: rom = 27;
		20354: rom = 27;
		20355: rom = 27;
		20356: rom = 27;
		20357: rom = 27;
		20358: rom = 20;
		20359: rom = 0;
		20360: rom = 0;
		20361: rom = 27;
		20362: rom = 27;
		20363: rom = 27;
		20364: rom = 27;
		20365: rom = 27;
		20366: rom = 27;
		20367: rom = 27;
		20368: rom = 16;
		20369: rom = 0;
		20370: rom = 0;
		20371: rom = 0;
		20372: rom = 24;
		20373: rom = 27;
		20374: rom = 27;
		20375: rom = 27;
		20376: rom = 27;
		20377: rom = 27;
		20378: rom = 27;
		20379: rom = 27;
		20380: rom = 0;
		20381: rom = 0;
		20382: rom = 20;
		20383: rom = 27;
		20384: rom = 27;
		20385: rom = 27;
		20386: rom = 27;
		20387: rom = 27;
		20388: rom = 27;
		20389: rom = 27;
		20390: rom = 25;
		20391: rom = 12;
		20392: rom = 18;
		20393: rom = 18;
		20394: rom = 18;
		20395: rom = 18;
		20396: rom = 18;
		20397: rom = 18;
		20398: rom = 18;
		20399: rom = 18;
		20400: rom = 18;
		20401: rom = 18;
		20402: rom = 18;
		20403: rom = 18;
		20404: rom = 18;
		20405: rom = 18;
		20406: rom = 18;
		20407: rom = 14;
		20408: rom = 15;
		20409: rom = 18;
		20410: rom = 18;
		20411: rom = 18;
		20412: rom = 18;
		20413: rom = 18;
		20414: rom = 24;
		20415: rom = 25;
		20416: rom = 24;
		20417: rom = 19;
		20418: rom = 18;
		20419: rom = 11;
		20420: rom = 25;
		20421: rom = 27;
		20422: rom = 27;
		20423: rom = 27;
		20424: rom = 27;
		20425: rom = 27;
		20426: rom = 27;
		20427: rom = 27;
		20428: rom = 27;
		20429: rom = 27;
		20430: rom = 27;
		20431: rom = 27;
		20432: rom = 27;
		20433: rom = 27;
		20434: rom = 27;
		20435: rom = 27;
		20436: rom = 27;
		20437: rom = 27;
		20438: rom = 27;
		20439: rom = 27;
		20440: rom = 27;
		20441: rom = 27;
		20442: rom = 20;
		20443: rom = 2;
		20444: rom = 0;
		20445: rom = 0;
		20446: rom = 27;
		20447: rom = 27;
		20448: rom = 0;
		20449: rom = 0;
		20450: rom = 20;
		20451: rom = 27;
		20452: rom = 27;
		20453: rom = 27;
		20454: rom = 27;
		20455: rom = 27;
		20456: rom = 27;
		20457: rom = 27;
		20458: rom = 27;
		20459: rom = 27;
		20460: rom = 0;
		20461: rom = 0;
		20462: rom = 27;
		20463: rom = 27;
		20464: rom = 27;
		20465: rom = 27;
		20466: rom = 27;
		20467: rom = 27;
		20468: rom = 13;
		20469: rom = 0;
		20470: rom = 27;
		20471: rom = 21;
		20472: rom = 0;
		20473: rom = 0;
		20474: rom = 26;
		20480: rom = 27;
		20481: rom = 27;
		20482: rom = 27;
		20483: rom = 27;
		20484: rom = 27;
		20485: rom = 27;
		20486: rom = 20;
		20487: rom = 0;
		20488: rom = 0;
		20489: rom = 27;
		20490: rom = 27;
		20491: rom = 27;
		20492: rom = 27;
		20493: rom = 27;
		20494: rom = 27;
		20495: rom = 27;
		20496: rom = 27;
		20497: rom = 13;
		20498: rom = 0;
		20499: rom = 0;
		20500: rom = 6;
		20501: rom = 25;
		20502: rom = 27;
		20503: rom = 27;
		20504: rom = 27;
		20505: rom = 27;
		20506: rom = 27;
		20507: rom = 27;
		20508: rom = 0;
		20509: rom = 0;
		20510: rom = 20;
		20511: rom = 27;
		20512: rom = 27;
		20513: rom = 27;
		20514: rom = 27;
		20515: rom = 27;
		20516: rom = 27;
		20517: rom = 27;
		20518: rom = 27;
		20519: rom = 18;
		20520: rom = 16;
		20521: rom = 18;
		20522: rom = 18;
		20523: rom = 18;
		20524: rom = 18;
		20525: rom = 18;
		20526: rom = 18;
		20527: rom = 18;
		20528: rom = 18;
		20529: rom = 18;
		20530: rom = 18;
		20531: rom = 18;
		20532: rom = 18;
		20533: rom = 18;
		20534: rom = 18;
		20535: rom = 17;
		20536: rom = 18;
		20537: rom = 18;
		20538: rom = 18;
		20539: rom = 18;
		20540: rom = 18;
		20541: rom = 24;
		20542: rom = 25;
		20543: rom = 24;
		20544: rom = 19;
		20545: rom = 18;
		20546: rom = 18;
		20547: rom = 18;
		20548: rom = 11;
		20549: rom = 26;
		20550: rom = 27;
		20551: rom = 27;
		20552: rom = 27;
		20553: rom = 27;
		20554: rom = 27;
		20555: rom = 27;
		20556: rom = 27;
		20557: rom = 27;
		20558: rom = 27;
		20559: rom = 27;
		20560: rom = 27;
		20561: rom = 27;
		20562: rom = 27;
		20563: rom = 27;
		20564: rom = 27;
		20565: rom = 27;
		20566: rom = 27;
		20567: rom = 27;
		20568: rom = 27;
		20569: rom = 27;
		20570: rom = 25;
		20571: rom = 14;
		20572: rom = 0;
		20573: rom = 0;
		20574: rom = 0;
		20575: rom = 27;
		20576: rom = 27;
		20577: rom = 27;
		20578: rom = 27;
		20579: rom = 27;
		20580: rom = 27;
		20581: rom = 27;
		20582: rom = 27;
		20583: rom = 27;
		20584: rom = 27;
		20585: rom = 27;
		20586: rom = 27;
		20587: rom = 27;
		20588: rom = 0;
		20589: rom = 0;
		20590: rom = 27;
		20591: rom = 27;
		20592: rom = 27;
		20593: rom = 27;
		20594: rom = 27;
		20595: rom = 27;
		20596: rom = 13;
		20597: rom = 0;
		20598: rom = 27;
		20599: rom = 20;
		20600: rom = 0;
		20601: rom = 0;
		20602: rom = 27;
		20608: rom = 27;
		20609: rom = 27;
		20610: rom = 27;
		20611: rom = 27;
		20612: rom = 27;
		20613: rom = 27;
		20614: rom = 20;
		20615: rom = 0;
		20616: rom = 0;
		20617: rom = 27;
		20618: rom = 27;
		20619: rom = 27;
		20620: rom = 27;
		20621: rom = 27;
		20622: rom = 27;
		20623: rom = 27;
		20624: rom = 27;
		20625: rom = 26;
		20626: rom = 11;
		20627: rom = 0;
		20628: rom = 0;
		20629: rom = 8;
		20630: rom = 25;
		20631: rom = 27;
		20632: rom = 27;
		20633: rom = 27;
		20634: rom = 27;
		20635: rom = 25;
		20636: rom = 0;
		20637: rom = 0;
		20638: rom = 22;
		20639: rom = 27;
		20640: rom = 27;
		20641: rom = 27;
		20642: rom = 27;
		20643: rom = 27;
		20644: rom = 27;
		20645: rom = 27;
		20646: rom = 27;
		20647: rom = 26;
		20648: rom = 12;
		20649: rom = 18;
		20650: rom = 18;
		20651: rom = 18;
		20652: rom = 18;
		20653: rom = 18;
		20654: rom = 18;
		20655: rom = 18;
		20656: rom = 18;
		20657: rom = 18;
		20658: rom = 18;
		20659: rom = 18;
		20660: rom = 18;
		20661: rom = 18;
		20662: rom = 18;
		20663: rom = 18;
		20664: rom = 18;
		20665: rom = 18;
		20666: rom = 18;
		20667: rom = 18;
		20668: rom = 24;
		20669: rom = 25;
		20670: rom = 23;
		20671: rom = 19;
		20672: rom = 18;
		20673: rom = 18;
		20674: rom = 18;
		20675: rom = 18;
		20676: rom = 17;
		20677: rom = 13;
		20678: rom = 26;
		20679: rom = 27;
		20680: rom = 27;
		20681: rom = 27;
		20682: rom = 27;
		20683: rom = 27;
		20684: rom = 27;
		20685: rom = 27;
		20686: rom = 27;
		20687: rom = 27;
		20688: rom = 27;
		20689: rom = 27;
		20690: rom = 27;
		20691: rom = 27;
		20692: rom = 27;
		20693: rom = 27;
		20694: rom = 27;
		20695: rom = 27;
		20696: rom = 27;
		20697: rom = 27;
		20698: rom = 27;
		20699: rom = 27;
		20700: rom = 21;
		20701: rom = 6;
		20702: rom = 0;
		20703: rom = 0;
		20704: rom = 5;
		20705: rom = 27;
		20706: rom = 27;
		20707: rom = 27;
		20708: rom = 27;
		20709: rom = 27;
		20710: rom = 27;
		20711: rom = 27;
		20712: rom = 27;
		20713: rom = 27;
		20714: rom = 27;
		20715: rom = 27;
		20716: rom = 0;
		20717: rom = 0;
		20718: rom = 27;
		20719: rom = 27;
		20720: rom = 27;
		20721: rom = 27;
		20722: rom = 27;
		20723: rom = 27;
		20724: rom = 13;
		20725: rom = 0;
		20726: rom = 27;
		20727: rom = 18;
		20728: rom = 0;
		20729: rom = 8;
		20730: rom = 27;
		20736: rom = 27;
		20737: rom = 27;
		20738: rom = 27;
		20739: rom = 27;
		20740: rom = 27;
		20741: rom = 27;
		20742: rom = 22;
		20743: rom = 0;
		20744: rom = 0;
		20745: rom = 26;
		20746: rom = 27;
		20747: rom = 27;
		20748: rom = 27;
		20749: rom = 27;
		20750: rom = 27;
		20751: rom = 27;
		20752: rom = 27;
		20753: rom = 27;
		20754: rom = 26;
		20755: rom = 9;
		20756: rom = 0;
		20757: rom = 0;
		20758: rom = 11;
		20759: rom = 26;
		20760: rom = 27;
		20761: rom = 27;
		20762: rom = 27;
		20763: rom = 22;
		20764: rom = 0;
		20765: rom = 0;
		20766: rom = 25;
		20767: rom = 27;
		20768: rom = 27;
		20769: rom = 27;
		20770: rom = 27;
		20771: rom = 27;
		20772: rom = 27;
		20773: rom = 27;
		20774: rom = 27;
		20775: rom = 27;
		20776: rom = 18;
		20777: rom = 16;
		20778: rom = 18;
		20779: rom = 18;
		20780: rom = 18;
		20781: rom = 18;
		20782: rom = 18;
		20783: rom = 18;
		20784: rom = 18;
		20785: rom = 18;
		20786: rom = 18;
		20787: rom = 18;
		20788: rom = 18;
		20789: rom = 18;
		20790: rom = 18;
		20791: rom = 18;
		20792: rom = 18;
		20793: rom = 18;
		20794: rom = 18;
		20795: rom = 24;
		20796: rom = 25;
		20797: rom = 23;
		20798: rom = 19;
		20799: rom = 18;
		20800: rom = 18;
		20801: rom = 18;
		20802: rom = 18;
		20803: rom = 18;
		20804: rom = 18;
		20805: rom = 17;
		20806: rom = 13;
		20807: rom = 26;
		20808: rom = 27;
		20809: rom = 27;
		20810: rom = 27;
		20811: rom = 27;
		20812: rom = 27;
		20813: rom = 27;
		20814: rom = 27;
		20815: rom = 27;
		20816: rom = 27;
		20817: rom = 27;
		20818: rom = 27;
		20819: rom = 27;
		20820: rom = 27;
		20821: rom = 27;
		20822: rom = 27;
		20823: rom = 27;
		20824: rom = 27;
		20825: rom = 27;
		20826: rom = 27;
		20827: rom = 27;
		20828: rom = 27;
		20829: rom = 26;
		20830: rom = 14;
		20831: rom = 0;
		20832: rom = 0;
		20833: rom = 0;
		20834: rom = 12;
		20835: rom = 25;
		20836: rom = 27;
		20837: rom = 27;
		20838: rom = 27;
		20839: rom = 27;
		20840: rom = 27;
		20841: rom = 27;
		20842: rom = 27;
		20843: rom = 27;
		20844: rom = 0;
		20845: rom = 0;
		20846: rom = 27;
		20847: rom = 27;
		20848: rom = 27;
		20849: rom = 27;
		20850: rom = 27;
		20851: rom = 27;
		20852: rom = 13;
		20853: rom = 0;
		20854: rom = 27;
		20855: rom = 13;
		20856: rom = 0;
		20857: rom = 14;
		20858: rom = 27;
		20864: rom = 27;
		20865: rom = 27;
		20866: rom = 27;
		20867: rom = 27;
		20868: rom = 27;
		20869: rom = 27;
		20870: rom = 25;
		20871: rom = 0;
		20872: rom = 0;
		20873: rom = 22;
		20874: rom = 27;
		20875: rom = 27;
		20876: rom = 27;
		20877: rom = 27;
		20878: rom = 27;
		20879: rom = 27;
		20880: rom = 27;
		20881: rom = 27;
		20882: rom = 27;
		20883: rom = 25;
		20884: rom = 7;
		20885: rom = 0;
		20886: rom = 0;
		20887: rom = 13;
		20888: rom = 27;
		20889: rom = 27;
		20890: rom = 27;
		20891: rom = 17;
		20892: rom = 0;
		20893: rom = 7;
		20894: rom = 27;
		20895: rom = 27;
		20896: rom = 27;
		20897: rom = 27;
		20898: rom = 27;
		20899: rom = 27;
		20900: rom = 27;
		20901: rom = 27;
		20902: rom = 27;
		20903: rom = 27;
		20904: rom = 26;
		20905: rom = 11;
		20906: rom = 18;
		20907: rom = 18;
		20908: rom = 18;
		20909: rom = 18;
		20910: rom = 18;
		20911: rom = 18;
		20912: rom = 18;
		20913: rom = 18;
		20914: rom = 18;
		20915: rom = 18;
		20916: rom = 18;
		20917: rom = 18;
		20918: rom = 18;
		20919: rom = 18;
		20920: rom = 18;
		20921: rom = 18;
		20922: rom = 23;
		20923: rom = 25;
		20924: rom = 24;
		20925: rom = 19;
		20926: rom = 18;
		20927: rom = 18;
		20928: rom = 18;
		20929: rom = 18;
		20930: rom = 18;
		20931: rom = 18;
		20932: rom = 18;
		20933: rom = 18;
		20934: rom = 17;
		20935: rom = 13;
		20936: rom = 26;
		20937: rom = 27;
		20938: rom = 27;
		20939: rom = 27;
		20940: rom = 27;
		20941: rom = 27;
		20942: rom = 27;
		20943: rom = 27;
		20944: rom = 27;
		20945: rom = 27;
		20946: rom = 27;
		20947: rom = 27;
		20948: rom = 27;
		20949: rom = 27;
		20950: rom = 27;
		20951: rom = 27;
		20952: rom = 27;
		20953: rom = 27;
		20954: rom = 27;
		20955: rom = 27;
		20956: rom = 27;
		20957: rom = 27;
		20958: rom = 27;
		20959: rom = 21;
		20960: rom = 7;
		20961: rom = 0;
		20962: rom = 0;
		20963: rom = 2;
		20964: rom = 20;
		20965: rom = 27;
		20966: rom = 27;
		20967: rom = 27;
		20968: rom = 27;
		20969: rom = 27;
		20970: rom = 27;
		20971: rom = 0;
		20972: rom = 0;
		20973: rom = 0;
		20974: rom = 0;
		20975: rom = 27;
		20976: rom = 27;
		20977: rom = 27;
		20978: rom = 27;
		20979: rom = 27;
		20980: rom = 13;
		20981: rom = 0;
		20982: rom = 27;
		20983: rom = 0;
		20984: rom = 0;
		20985: rom = 19;
		20986: rom = 27;
		20992: rom = 27;
		20993: rom = 27;
		20994: rom = 27;
		20995: rom = 27;
		20996: rom = 27;
		20997: rom = 27;
		20998: rom = 27;
		20999: rom = 0;
		21000: rom = 0;
		21001: rom = 15;
		21002: rom = 27;
		21003: rom = 27;
		21004: rom = 27;
		21005: rom = 27;
		21006: rom = 27;
		21007: rom = 27;
		21008: rom = 27;
		21009: rom = 27;
		21010: rom = 27;
		21011: rom = 27;
		21012: rom = 24;
		21013: rom = 0;
		21014: rom = 0;
		21015: rom = 0;
		21016: rom = 15;
		21017: rom = 27;
		21018: rom = 25;
		21019: rom = 0;
		21020: rom = 0;
		21021: rom = 17;
		21022: rom = 27;
		21023: rom = 27;
		21024: rom = 27;
		21025: rom = 27;
		21026: rom = 27;
		21027: rom = 27;
		21028: rom = 27;
		21029: rom = 27;
		21030: rom = 27;
		21031: rom = 27;
		21032: rom = 27;
		21033: rom = 20;
		21034: rom = 15;
		21035: rom = 18;
		21036: rom = 18;
		21037: rom = 18;
		21038: rom = 18;
		21039: rom = 18;
		21040: rom = 18;
		21041: rom = 18;
		21042: rom = 18;
		21043: rom = 18;
		21044: rom = 18;
		21045: rom = 18;
		21046: rom = 18;
		21047: rom = 18;
		21048: rom = 18;
		21049: rom = 22;
		21050: rom = 25;
		21051: rom = 24;
		21052: rom = 19;
		21053: rom = 18;
		21054: rom = 18;
		21055: rom = 18;
		21056: rom = 18;
		21057: rom = 18;
		21058: rom = 18;
		21059: rom = 18;
		21060: rom = 18;
		21061: rom = 18;
		21062: rom = 18;
		21063: rom = 17;
		21064: rom = 13;
		21065: rom = 26;
		21066: rom = 27;
		21067: rom = 27;
		21068: rom = 27;
		21069: rom = 27;
		21070: rom = 27;
		21071: rom = 27;
		21072: rom = 27;
		21073: rom = 27;
		21074: rom = 27;
		21075: rom = 27;
		21076: rom = 27;
		21077: rom = 27;
		21078: rom = 27;
		21079: rom = 27;
		21080: rom = 27;
		21081: rom = 27;
		21082: rom = 27;
		21083: rom = 27;
		21084: rom = 27;
		21085: rom = 27;
		21086: rom = 27;
		21087: rom = 27;
		21088: rom = 25;
		21089: rom = 14;
		21090: rom = 0;
		21091: rom = 0;
		21092: rom = 0;
		21093: rom = 12;
		21094: rom = 24;
		21095: rom = 27;
		21096: rom = 27;
		21097: rom = 27;
		21098: rom = 27;
		21099: rom = 27;
		21100: rom = 27;
		21101: rom = 27;
		21102: rom = 27;
		21103: rom = 27;
		21104: rom = 27;
		21105: rom = 27;
		21106: rom = 27;
		21107: rom = 27;
		21108: rom = 13;
		21109: rom = 0;
		21110: rom = 27;
		21111: rom = 0;
		21112: rom = 0;
		21113: rom = 24;
		21114: rom = 27;
		21120: rom = 27;
		21121: rom = 27;
		21122: rom = 27;
		21123: rom = 27;
		21124: rom = 27;
		21125: rom = 27;
		21126: rom = 27;
		21127: rom = 18;
		21128: rom = 0;
		21129: rom = 0;
		21130: rom = 26;
		21131: rom = 27;
		21132: rom = 27;
		21133: rom = 27;
		21134: rom = 27;
		21135: rom = 27;
		21136: rom = 27;
		21137: rom = 27;
		21138: rom = 27;
		21139: rom = 27;
		21140: rom = 27;
		21141: rom = 23;
		21142: rom = 0;
		21143: rom = 0;
		21144: rom = 0;
		21145: rom = 17;
		21146: rom = 15;
		21147: rom = 0;
		21148: rom = 0;
		21149: rom = 25;
		21150: rom = 27;
		21151: rom = 27;
		21152: rom = 27;
		21153: rom = 27;
		21154: rom = 27;
		21155: rom = 27;
		21156: rom = 27;
		21157: rom = 27;
		21158: rom = 27;
		21159: rom = 27;
		21160: rom = 27;
		21161: rom = 27;
		21162: rom = 13;
		21163: rom = 17;
		21164: rom = 18;
		21165: rom = 18;
		21166: rom = 18;
		21167: rom = 18;
		21168: rom = 18;
		21169: rom = 18;
		21170: rom = 18;
		21171: rom = 18;
		21172: rom = 18;
		21173: rom = 18;
		21174: rom = 18;
		21175: rom = 18;
		21176: rom = 19;
		21177: rom = 25;
		21178: rom = 25;
		21179: rom = 19;
		21180: rom = 18;
		21181: rom = 18;
		21182: rom = 18;
		21183: rom = 18;
		21184: rom = 18;
		21185: rom = 18;
		21186: rom = 18;
		21187: rom = 18;
		21188: rom = 18;
		21189: rom = 18;
		21190: rom = 18;
		21191: rom = 18;
		21192: rom = 17;
		21193: rom = 12;
		21194: rom = 25;
		21195: rom = 27;
		21196: rom = 27;
		21197: rom = 27;
		21198: rom = 27;
		21199: rom = 27;
		21200: rom = 27;
		21201: rom = 27;
		21202: rom = 27;
		21203: rom = 27;
		21204: rom = 27;
		21205: rom = 27;
		21206: rom = 27;
		21207: rom = 27;
		21208: rom = 27;
		21209: rom = 27;
		21210: rom = 27;
		21211: rom = 27;
		21212: rom = 27;
		21213: rom = 27;
		21214: rom = 27;
		21215: rom = 27;
		21216: rom = 27;
		21217: rom = 27;
		21218: rom = 27;
		21219: rom = 27;
		21220: rom = 0;
		21221: rom = 0;
		21222: rom = 2;
		21223: rom = 19;
		21224: rom = 27;
		21225: rom = 27;
		21226: rom = 27;
		21227: rom = 27;
		21228: rom = 27;
		21229: rom = 27;
		21230: rom = 27;
		21231: rom = 27;
		21232: rom = 27;
		21233: rom = 27;
		21234: rom = 27;
		21235: rom = 27;
		21236: rom = 13;
		21237: rom = 0;
		21238: rom = 27;
		21239: rom = 0;
		21240: rom = 9;
		21241: rom = 27;
		21242: rom = 27;
		21248: rom = 27;
		21249: rom = 27;
		21250: rom = 27;
		21251: rom = 27;
		21252: rom = 27;
		21253: rom = 27;
		21254: rom = 27;
		21255: rom = 27;
		21256: rom = 27;
		21257: rom = 27;
		21258: rom = 27;
		21259: rom = 27;
		21260: rom = 27;
		21261: rom = 27;
		21262: rom = 27;
		21263: rom = 27;
		21264: rom = 27;
		21265: rom = 27;
		21266: rom = 27;
		21267: rom = 27;
		21268: rom = 27;
		21269: rom = 27;
		21270: rom = 21;
		21271: rom = 0;
		21272: rom = 0;
		21273: rom = 0;
		21274: rom = 0;
		21275: rom = 0;
		21276: rom = 17;
		21277: rom = 27;
		21278: rom = 27;
		21279: rom = 27;
		21280: rom = 27;
		21281: rom = 27;
		21282: rom = 27;
		21283: rom = 27;
		21284: rom = 27;
		21285: rom = 27;
		21286: rom = 27;
		21287: rom = 27;
		21288: rom = 27;
		21289: rom = 27;
		21290: rom = 24;
		21291: rom = 12;
		21292: rom = 18;
		21293: rom = 18;
		21294: rom = 18;
		21295: rom = 18;
		21296: rom = 18;
		21297: rom = 18;
		21298: rom = 18;
		21299: rom = 18;
		21300: rom = 18;
		21301: rom = 18;
		21302: rom = 18;
		21303: rom = 18;
		21304: rom = 23;
		21305: rom = 25;
		21306: rom = 21;
		21307: rom = 18;
		21308: rom = 18;
		21309: rom = 18;
		21310: rom = 18;
		21311: rom = 18;
		21312: rom = 18;
		21313: rom = 18;
		21314: rom = 18;
		21315: rom = 18;
		21316: rom = 18;
		21317: rom = 18;
		21318: rom = 18;
		21319: rom = 18;
		21320: rom = 18;
		21321: rom = 17;
		21322: rom = 12;
		21323: rom = 25;
		21324: rom = 27;
		21325: rom = 27;
		21326: rom = 27;
		21327: rom = 27;
		21328: rom = 27;
		21329: rom = 27;
		21330: rom = 27;
		21331: rom = 27;
		21332: rom = 27;
		21333: rom = 27;
		21334: rom = 27;
		21335: rom = 27;
		21336: rom = 27;
		21337: rom = 27;
		21338: rom = 27;
		21339: rom = 27;
		21340: rom = 27;
		21341: rom = 27;
		21342: rom = 27;
		21343: rom = 27;
		21344: rom = 27;
		21345: rom = 20;
		21346: rom = 0;
		21347: rom = 27;
		21348: rom = 27;
		21349: rom = 0;
		21350: rom = 0;
		21351: rom = 0;
		21352: rom = 11;
		21353: rom = 24;
		21354: rom = 27;
		21355: rom = 27;
		21356: rom = 27;
		21357: rom = 27;
		21358: rom = 27;
		21359: rom = 27;
		21360: rom = 27;
		21361: rom = 27;
		21362: rom = 27;
		21363: rom = 27;
		21364: rom = 13;
		21365: rom = 0;
		21366: rom = 27;
		21367: rom = 0;
		21368: rom = 20;
		21369: rom = 27;
		21370: rom = 27;
		21376: rom = 27;
		21377: rom = 27;
		21378: rom = 27;
		21379: rom = 27;
		21380: rom = 27;
		21381: rom = 27;
		21382: rom = 27;
		21383: rom = 27;
		21384: rom = 27;
		21385: rom = 27;
		21386: rom = 27;
		21387: rom = 27;
		21388: rom = 27;
		21389: rom = 27;
		21390: rom = 27;
		21391: rom = 27;
		21392: rom = 27;
		21393: rom = 27;
		21394: rom = 27;
		21395: rom = 27;
		21396: rom = 27;
		21397: rom = 27;
		21398: rom = 27;
		21399: rom = 19;
		21400: rom = 0;
		21401: rom = 0;
		21402: rom = 0;
		21403: rom = 8;
		21404: rom = 26;
		21405: rom = 27;
		21406: rom = 27;
		21407: rom = 27;
		21408: rom = 27;
		21409: rom = 27;
		21410: rom = 27;
		21411: rom = 27;
		21412: rom = 27;
		21413: rom = 27;
		21414: rom = 27;
		21415: rom = 27;
		21416: rom = 27;
		21417: rom = 27;
		21418: rom = 27;
		21419: rom = 19;
		21420: rom = 15;
		21421: rom = 18;
		21422: rom = 18;
		21423: rom = 18;
		21424: rom = 18;
		21425: rom = 18;
		21426: rom = 18;
		21427: rom = 18;
		21428: rom = 18;
		21429: rom = 18;
		21430: rom = 18;
		21431: rom = 18;
		21432: rom = 23;
		21433: rom = 25;
		21434: rom = 19;
		21435: rom = 18;
		21436: rom = 18;
		21437: rom = 18;
		21438: rom = 18;
		21439: rom = 18;
		21440: rom = 18;
		21441: rom = 18;
		21442: rom = 18;
		21443: rom = 18;
		21444: rom = 18;
		21445: rom = 18;
		21446: rom = 18;
		21447: rom = 18;
		21448: rom = 18;
		21449: rom = 18;
		21450: rom = 18;
		21451: rom = 11;
		21452: rom = 24;
		21453: rom = 27;
		21454: rom = 27;
		21455: rom = 27;
		21456: rom = 27;
		21457: rom = 27;
		21458: rom = 27;
		21459: rom = 27;
		21460: rom = 27;
		21461: rom = 27;
		21462: rom = 27;
		21463: rom = 27;
		21464: rom = 27;
		21465: rom = 27;
		21466: rom = 27;
		21467: rom = 27;
		21468: rom = 27;
		21469: rom = 27;
		21470: rom = 27;
		21471: rom = 27;
		21472: rom = 27;
		21473: rom = 27;
		21474: rom = 9;
		21475: rom = 0;
		21476: rom = 27;
		21477: rom = 27;
		21478: rom = 8;
		21479: rom = 0;
		21480: rom = 0;
		21481: rom = 1;
		21482: rom = 18;
		21483: rom = 27;
		21484: rom = 27;
		21485: rom = 27;
		21486: rom = 27;
		21487: rom = 27;
		21488: rom = 27;
		21489: rom = 27;
		21490: rom = 27;
		21491: rom = 27;
		21492: rom = 13;
		21493: rom = 0;
		21494: rom = 27;
		21495: rom = 8;
		21496: rom = 27;
		21497: rom = 27;
		21498: rom = 27;
		21504: rom = 27;
		21505: rom = 27;
		21506: rom = 27;
		21507: rom = 27;
		21508: rom = 27;
		21509: rom = 27;
		21510: rom = 27;
		21511: rom = 27;
		21512: rom = 27;
		21513: rom = 27;
		21514: rom = 27;
		21515: rom = 27;
		21516: rom = 27;
		21517: rom = 27;
		21518: rom = 27;
		21519: rom = 27;
		21520: rom = 27;
		21521: rom = 27;
		21522: rom = 27;
		21523: rom = 27;
		21524: rom = 27;
		21525: rom = 27;
		21526: rom = 26;
		21527: rom = 15;
		21528: rom = 0;
		21529: rom = 0;
		21530: rom = 0;
		21531: rom = 0;
		21532: rom = 23;
		21533: rom = 27;
		21534: rom = 27;
		21535: rom = 27;
		21536: rom = 27;
		21537: rom = 27;
		21538: rom = 27;
		21539: rom = 27;
		21540: rom = 27;
		21541: rom = 27;
		21542: rom = 27;
		21543: rom = 27;
		21544: rom = 27;
		21545: rom = 27;
		21546: rom = 27;
		21547: rom = 27;
		21548: rom = 14;
		21549: rom = 16;
		21550: rom = 18;
		21551: rom = 18;
		21552: rom = 18;
		21553: rom = 18;
		21554: rom = 18;
		21555: rom = 18;
		21556: rom = 18;
		21557: rom = 18;
		21558: rom = 18;
		21559: rom = 18;
		21560: rom = 21;
		21561: rom = 25;
		21562: rom = 21;
		21563: rom = 18;
		21564: rom = 18;
		21565: rom = 18;
		21566: rom = 18;
		21567: rom = 18;
		21568: rom = 18;
		21569: rom = 18;
		21570: rom = 18;
		21571: rom = 18;
		21572: rom = 18;
		21573: rom = 18;
		21574: rom = 18;
		21575: rom = 18;
		21576: rom = 18;
		21577: rom = 18;
		21578: rom = 18;
		21579: rom = 18;
		21580: rom = 11;
		21581: rom = 23;
		21582: rom = 27;
		21583: rom = 27;
		21584: rom = 27;
		21585: rom = 27;
		21586: rom = 27;
		21587: rom = 27;
		21588: rom = 27;
		21589: rom = 27;
		21590: rom = 27;
		21591: rom = 27;
		21592: rom = 27;
		21593: rom = 27;
		21594: rom = 27;
		21595: rom = 27;
		21596: rom = 27;
		21597: rom = 27;
		21598: rom = 27;
		21599: rom = 27;
		21600: rom = 27;
		21601: rom = 27;
		21602: rom = 23;
		21603: rom = 0;
		21604: rom = 0;
		21605: rom = 27;
		21606: rom = 27;
		21607: rom = 27;
		21608: rom = 0;
		21609: rom = 0;
		21610: rom = 0;
		21611: rom = 9;
		21612: rom = 23;
		21613: rom = 27;
		21614: rom = 27;
		21615: rom = 27;
		21616: rom = 27;
		21617: rom = 27;
		21618: rom = 27;
		21619: rom = 26;
		21620: rom = 13;
		21621: rom = 0;
		21622: rom = 27;
		21623: rom = 22;
		21624: rom = 27;
		21625: rom = 27;
		21626: rom = 27;
		21632: rom = 27;
		21633: rom = 27;
		21634: rom = 27;
		21635: rom = 27;
		21636: rom = 27;
		21637: rom = 27;
		21638: rom = 27;
		21639: rom = 27;
		21640: rom = 27;
		21641: rom = 27;
		21642: rom = 27;
		21643: rom = 27;
		21644: rom = 27;
		21645: rom = 27;
		21646: rom = 27;
		21647: rom = 27;
		21648: rom = 27;
		21649: rom = 27;
		21650: rom = 27;
		21651: rom = 27;
		21652: rom = 24;
		21653: rom = 17;
		21654: rom = 0;
		21655: rom = 0;
		21656: rom = 0;
		21657: rom = 3;
		21658: rom = 0;
		21659: rom = 0;
		21660: rom = 0;
		21661: rom = 24;
		21662: rom = 27;
		21663: rom = 27;
		21664: rom = 27;
		21665: rom = 27;
		21666: rom = 27;
		21667: rom = 27;
		21668: rom = 27;
		21669: rom = 27;
		21670: rom = 27;
		21671: rom = 27;
		21672: rom = 27;
		21673: rom = 27;
		21674: rom = 27;
		21675: rom = 27;
		21676: rom = 26;
		21677: rom = 12;
		21678: rom = 17;
		21679: rom = 18;
		21680: rom = 18;
		21681: rom = 18;
		21682: rom = 18;
		21683: rom = 18;
		21684: rom = 18;
		21685: rom = 18;
		21686: rom = 18;
		21687: rom = 18;
		21688: rom = 19;
		21689: rom = 25;
		21690: rom = 24;
		21691: rom = 18;
		21692: rom = 18;
		21693: rom = 18;
		21694: rom = 18;
		21695: rom = 18;
		21696: rom = 18;
		21697: rom = 18;
		21698: rom = 18;
		21699: rom = 18;
		21700: rom = 18;
		21701: rom = 18;
		21702: rom = 18;
		21703: rom = 18;
		21704: rom = 18;
		21705: rom = 18;
		21706: rom = 18;
		21707: rom = 18;
		21708: rom = 18;
		21709: rom = 12;
		21710: rom = 22;
		21711: rom = 27;
		21712: rom = 27;
		21713: rom = 27;
		21714: rom = 27;
		21715: rom = 27;
		21716: rom = 27;
		21717: rom = 27;
		21718: rom = 27;
		21719: rom = 27;
		21720: rom = 27;
		21721: rom = 27;
		21722: rom = 27;
		21723: rom = 27;
		21724: rom = 27;
		21725: rom = 27;
		21726: rom = 27;
		21727: rom = 27;
		21728: rom = 27;
		21729: rom = 27;
		21730: rom = 27;
		21731: rom = 18;
		21732: rom = 0;
		21733: rom = 0;
		21734: rom = 8;
		21735: rom = 27;
		21736: rom = 27;
		21737: rom = 9;
		21738: rom = 0;
		21739: rom = 0;
		21740: rom = 0;
		21741: rom = 17;
		21742: rom = 26;
		21743: rom = 27;
		21744: rom = 27;
		21745: rom = 27;
		21746: rom = 23;
		21747: rom = 27;
		21748: rom = 13;
		21749: rom = 0;
		21750: rom = 27;
		21751: rom = 27;
		21752: rom = 27;
		21753: rom = 27;
		21754: rom = 27;
		21760: rom = 27;
		21761: rom = 27;
		21762: rom = 27;
		21763: rom = 27;
		21764: rom = 27;
		21765: rom = 27;
		21766: rom = 27;
		21767: rom = 27;
		21768: rom = 27;
		21769: rom = 27;
		21770: rom = 27;
		21771: rom = 27;
		21772: rom = 27;
		21773: rom = 27;
		21774: rom = 27;
		21775: rom = 27;
		21776: rom = 27;
		21777: rom = 23;
		21778: rom = 13;
		21779: rom = 0;
		21780: rom = 0;
		21781: rom = 0;
		21782: rom = 0;
		21783: rom = 0;
		21784: rom = 14;
		21785: rom = 26;
		21786: rom = 12;
		21787: rom = 0;
		21788: rom = 0;
		21789: rom = 0;
		21790: rom = 27;
		21791: rom = 27;
		21792: rom = 27;
		21793: rom = 27;
		21794: rom = 27;
		21795: rom = 27;
		21796: rom = 27;
		21797: rom = 27;
		21798: rom = 27;
		21799: rom = 27;
		21800: rom = 27;
		21801: rom = 27;
		21802: rom = 27;
		21803: rom = 27;
		21804: rom = 27;
		21805: rom = 25;
		21806: rom = 11;
		21807: rom = 17;
		21808: rom = 18;
		21809: rom = 18;
		21810: rom = 18;
		21811: rom = 18;
		21812: rom = 18;
		21813: rom = 15;
		21814: rom = 18;
		21815: rom = 18;
		21816: rom = 18;
		21817: rom = 24;
		21818: rom = 25;
		21819: rom = 19;
		21820: rom = 18;
		21821: rom = 18;
		21822: rom = 18;
		21823: rom = 18;
		21824: rom = 18;
		21825: rom = 18;
		21826: rom = 18;
		21827: rom = 18;
		21828: rom = 18;
		21829: rom = 18;
		21830: rom = 18;
		21831: rom = 18;
		21832: rom = 18;
		21833: rom = 18;
		21834: rom = 18;
		21835: rom = 18;
		21836: rom = 18;
		21837: rom = 18;
		21838: rom = 13;
		21839: rom = 22;
		21840: rom = 27;
		21841: rom = 27;
		21842: rom = 27;
		21843: rom = 27;
		21844: rom = 27;
		21845: rom = 27;
		21846: rom = 27;
		21847: rom = 27;
		21848: rom = 27;
		21849: rom = 27;
		21850: rom = 27;
		21851: rom = 27;
		21852: rom = 27;
		21853: rom = 27;
		21854: rom = 27;
		21855: rom = 27;
		21856: rom = 27;
		21857: rom = 27;
		21858: rom = 27;
		21859: rom = 27;
		21860: rom = 15;
		21861: rom = 0;
		21862: rom = 0;
		21863: rom = 1;
		21864: rom = 27;
		21865: rom = 27;
		21866: rom = 27;
		21867: rom = 1;
		21868: rom = 0;
		21869: rom = 0;
		21870: rom = 27;
		21871: rom = 27;
		21872: rom = 24;
		21873: rom = 15;
		21874: rom = 0;
		21875: rom = 27;
		21876: rom = 13;
		21877: rom = 0;
		21878: rom = 27;
		21879: rom = 27;
		21880: rom = 27;
		21881: rom = 27;
		21882: rom = 27;
		21888: rom = 27;
		21889: rom = 27;
		21890: rom = 27;
		21891: rom = 27;
		21892: rom = 27;
		21893: rom = 27;
		21894: rom = 27;
		21895: rom = 27;
		21896: rom = 27;
		21897: rom = 27;
		21898: rom = 27;
		21899: rom = 27;
		21900: rom = 27;
		21901: rom = 27;
		21902: rom = 27;
		21903: rom = 27;
		21904: rom = 27;
		21905: rom = 21;
		21906: rom = 0;
		21907: rom = 0;
		21908: rom = 0;
		21909: rom = 0;
		21910: rom = 0;
		21911: rom = 21;
		21912: rom = 27;
		21913: rom = 27;
		21914: rom = 26;
		21915: rom = 10;
		21916: rom = 0;
		21917: rom = 0;
		21918: rom = 27;
		21919: rom = 27;
		21920: rom = 27;
		21921: rom = 27;
		21922: rom = 27;
		21923: rom = 27;
		21924: rom = 27;
		21925: rom = 27;
		21926: rom = 27;
		21927: rom = 27;
		21928: rom = 27;
		21929: rom = 27;
		21930: rom = 27;
		21931: rom = 27;
		21932: rom = 27;
		21933: rom = 27;
		21934: rom = 25;
		21935: rom = 11;
		21936: rom = 17;
		21937: rom = 18;
		21938: rom = 18;
		21939: rom = 18;
		21940: rom = 18;
		21941: rom = 7;
		21942: rom = 16;
		21943: rom = 18;
		21944: rom = 18;
		21945: rom = 21;
		21946: rom = 25;
		21947: rom = 22;
		21948: rom = 18;
		21949: rom = 18;
		21950: rom = 18;
		21951: rom = 18;
		21952: rom = 18;
		21953: rom = 18;
		21954: rom = 18;
		21955: rom = 18;
		21956: rom = 18;
		21957: rom = 18;
		21958: rom = 18;
		21959: rom = 18;
		21960: rom = 18;
		21961: rom = 18;
		21962: rom = 18;
		21963: rom = 18;
		21964: rom = 18;
		21965: rom = 18;
		21966: rom = 14;
		21967: rom = 14;
		21968: rom = 27;
		21969: rom = 27;
		21970: rom = 27;
		21971: rom = 27;
		21972: rom = 27;
		21973: rom = 27;
		21974: rom = 27;
		21975: rom = 27;
		21976: rom = 27;
		21977: rom = 27;
		21978: rom = 27;
		21979: rom = 27;
		21980: rom = 27;
		21981: rom = 27;
		21982: rom = 27;
		21983: rom = 27;
		21984: rom = 27;
		21985: rom = 27;
		21986: rom = 27;
		21987: rom = 27;
		21988: rom = 27;
		21989: rom = 16;
		21990: rom = 0;
		21991: rom = 0;
		21992: rom = 0;
		21993: rom = 0;
		21994: rom = 27;
		21995: rom = 27;
		21996: rom = 27;
		21997: rom = 27;
		21998: rom = 27;
		21999: rom = 10;
		22000: rom = 0;
		22001: rom = 0;
		22002: rom = 0;
		22003: rom = 27;
		22004: rom = 13;
		22005: rom = 0;
		22006: rom = 27;
		22007: rom = 27;
		22008: rom = 27;
		22009: rom = 27;
		22010: rom = 27;
		22016: rom = 27;
		22017: rom = 27;
		22018: rom = 27;
		22019: rom = 27;
		22020: rom = 27;
		22021: rom = 27;
		22022: rom = 27;
		22023: rom = 27;
		22024: rom = 27;
		22025: rom = 27;
		22026: rom = 27;
		22027: rom = 27;
		22028: rom = 27;
		22029: rom = 27;
		22030: rom = 27;
		22031: rom = 27;
		22032: rom = 27;
		22033: rom = 21;
		22034: rom = 0;
		22035: rom = 0;
		22036: rom = 9;
		22037: rom = 19;
		22038: rom = 26;
		22039: rom = 27;
		22040: rom = 27;
		22041: rom = 27;
		22042: rom = 27;
		22043: rom = 25;
		22044: rom = 0;
		22045: rom = 0;
		22046: rom = 27;
		22047: rom = 27;
		22048: rom = 27;
		22049: rom = 27;
		22050: rom = 27;
		22051: rom = 27;
		22052: rom = 27;
		22053: rom = 27;
		22054: rom = 27;
		22055: rom = 27;
		22056: rom = 27;
		22057: rom = 27;
		22058: rom = 27;
		22059: rom = 27;
		22060: rom = 27;
		22061: rom = 27;
		22062: rom = 27;
		22063: rom = 25;
		22064: rom = 11;
		22065: rom = 17;
		22066: rom = 18;
		22067: rom = 18;
		22068: rom = 18;
		22069: rom = 6;
		22070: rom = 14;
		22071: rom = 18;
		22072: rom = 18;
		22073: rom = 18;
		22074: rom = 25;
		22075: rom = 25;
		22076: rom = 19;
		22077: rom = 18;
		22078: rom = 18;
		22079: rom = 18;
		22080: rom = 18;
		22081: rom = 18;
		22082: rom = 18;
		22083: rom = 18;
		22084: rom = 18;
		22085: rom = 18;
		22086: rom = 18;
		22087: rom = 18;
		22088: rom = 18;
		22089: rom = 18;
		22090: rom = 18;
		22091: rom = 18;
		22092: rom = 14;
		22093: rom = 12;
		22094: rom = 22;
		22095: rom = 27;
		22096: rom = 27;
		22097: rom = 27;
		22098: rom = 27;
		22099: rom = 27;
		22100: rom = 27;
		22101: rom = 27;
		22102: rom = 27;
		22103: rom = 27;
		22104: rom = 27;
		22105: rom = 27;
		22106: rom = 27;
		22107: rom = 27;
		22108: rom = 27;
		22109: rom = 27;
		22110: rom = 27;
		22111: rom = 27;
		22112: rom = 27;
		22113: rom = 27;
		22114: rom = 27;
		22115: rom = 27;
		22116: rom = 27;
		22117: rom = 27;
		22118: rom = 21;
		22119: rom = 6;
		22120: rom = 0;
		22121: rom = 0;
		22122: rom = 0;
		22123: rom = 0;
		22124: rom = 0;
		22125: rom = 0;
		22126: rom = 0;
		22127: rom = 0;
		22128: rom = 0;
		22129: rom = 0;
		22130: rom = 27;
		22131: rom = 27;
		22132: rom = 13;
		22133: rom = 0;
		22134: rom = 19;
		22135: rom = 27;
		22136: rom = 27;
		22137: rom = 27;
		22138: rom = 27;
		22144: rom = 27;
		22145: rom = 27;
		22146: rom = 27;
		22147: rom = 27;
		22148: rom = 27;
		22149: rom = 27;
		22150: rom = 27;
		22151: rom = 27;
		22152: rom = 27;
		22153: rom = 27;
		22154: rom = 27;
		22155: rom = 27;
		22156: rom = 27;
		22157: rom = 27;
		22158: rom = 27;
		22159: rom = 27;
		22160: rom = 27;
		22161: rom = 24;
		22162: rom = 21;
		22163: rom = 24;
		22164: rom = 27;
		22165: rom = 27;
		22166: rom = 27;
		22167: rom = 27;
		22168: rom = 27;
		22169: rom = 27;
		22170: rom = 27;
		22171: rom = 27;
		22172: rom = 24;
		22173: rom = 0;
		22174: rom = 27;
		22175: rom = 27;
		22176: rom = 27;
		22177: rom = 27;
		22178: rom = 27;
		22179: rom = 27;
		22180: rom = 27;
		22181: rom = 27;
		22182: rom = 27;
		22183: rom = 27;
		22184: rom = 27;
		22185: rom = 27;
		22186: rom = 27;
		22187: rom = 27;
		22188: rom = 27;
		22189: rom = 27;
		22190: rom = 27;
		22191: rom = 27;
		22192: rom = 25;
		22193: rom = 12;
		22194: rom = 15;
		22195: rom = 18;
		22196: rom = 18;
		22197: rom = 14;
		22198: rom = 11;
		22199: rom = 18;
		22200: rom = 18;
		22201: rom = 18;
		22202: rom = 22;
		22203: rom = 25;
		22204: rom = 22;
		22205: rom = 18;
		22206: rom = 18;
		22207: rom = 18;
		22208: rom = 18;
		22209: rom = 18;
		22210: rom = 18;
		22211: rom = 18;
		22212: rom = 18;
		22213: rom = 18;
		22214: rom = 18;
		22215: rom = 18;
		22216: rom = 18;
		22217: rom = 17;
		22218: rom = 12;
		22219: rom = 14;
		22220: rom = 22;
		22221: rom = 27;
		22222: rom = 27;
		22223: rom = 27;
		22224: rom = 27;
		22225: rom = 27;
		22226: rom = 27;
		22227: rom = 27;
		22228: rom = 27;
		22229: rom = 27;
		22230: rom = 27;
		22231: rom = 27;
		22232: rom = 27;
		22233: rom = 27;
		22234: rom = 27;
		22235: rom = 27;
		22236: rom = 27;
		22237: rom = 27;
		22238: rom = 27;
		22239: rom = 27;
		22240: rom = 27;
		22241: rom = 27;
		22242: rom = 27;
		22243: rom = 27;
		22244: rom = 27;
		22245: rom = 27;
		22246: rom = 27;
		22247: rom = 26;
		22248: rom = 19;
		22249: rom = 8;
		22250: rom = 0;
		22251: rom = 0;
		22252: rom = 0;
		22253: rom = 0;
		22254: rom = 0;
		22255: rom = 0;
		22256: rom = 27;
		22257: rom = 27;
		22258: rom = 27;
		22259: rom = 18;
		22260: rom = 11;
		22261: rom = 0;
		22262: rom = 19;
		22263: rom = 27;
		22264: rom = 27;
		22265: rom = 27;
		22266: rom = 27;
		22272: rom = 27;
		22273: rom = 27;
		22274: rom = 27;
		22275: rom = 27;
		22276: rom = 27;
		22277: rom = 27;
		22278: rom = 27;
		22279: rom = 27;
		22280: rom = 27;
		22281: rom = 27;
		22282: rom = 27;
		22283: rom = 27;
		22284: rom = 27;
		22285: rom = 27;
		22286: rom = 27;
		22287: rom = 27;
		22288: rom = 27;
		22289: rom = 27;
		22290: rom = 27;
		22291: rom = 27;
		22292: rom = 27;
		22293: rom = 27;
		22294: rom = 27;
		22295: rom = 27;
		22296: rom = 27;
		22297: rom = 27;
		22298: rom = 27;
		22299: rom = 27;
		22300: rom = 27;
		22301: rom = 23;
		22302: rom = 27;
		22303: rom = 27;
		22304: rom = 27;
		22305: rom = 27;
		22306: rom = 27;
		22307: rom = 27;
		22308: rom = 27;
		22309: rom = 27;
		22310: rom = 27;
		22311: rom = 27;
		22312: rom = 27;
		22313: rom = 27;
		22314: rom = 27;
		22315: rom = 27;
		22316: rom = 27;
		22317: rom = 27;
		22318: rom = 27;
		22319: rom = 27;
		22320: rom = 27;
		22321: rom = 26;
		22322: rom = 15;
		22323: rom = 13;
		22324: rom = 17;
		22325: rom = 15;
		22326: rom = 15;
		22327: rom = 17;
		22328: rom = 18;
		22329: rom = 18;
		22330: rom = 18;
		22331: rom = 25;
		22332: rom = 25;
		22333: rom = 19;
		22334: rom = 18;
		22335: rom = 18;
		22336: rom = 18;
		22337: rom = 18;
		22338: rom = 18;
		22339: rom = 18;
		22340: rom = 18;
		22341: rom = 18;
		22342: rom = 17;
		22343: rom = 14;
		22344: rom = 11;
		22345: rom = 18;
		22346: rom = 24;
		22347: rom = 27;
		22348: rom = 27;
		22349: rom = 27;
		22350: rom = 27;
		22351: rom = 27;
		22352: rom = 27;
		22353: rom = 27;
		22354: rom = 27;
		22355: rom = 27;
		22356: rom = 27;
		22357: rom = 27;
		22358: rom = 27;
		22359: rom = 27;
		22360: rom = 27;
		22361: rom = 27;
		22362: rom = 27;
		22363: rom = 27;
		22364: rom = 27;
		22365: rom = 27;
		22366: rom = 27;
		22367: rom = 27;
		22368: rom = 27;
		22369: rom = 27;
		22370: rom = 27;
		22371: rom = 27;
		22372: rom = 27;
		22373: rom = 27;
		22374: rom = 27;
		22375: rom = 27;
		22376: rom = 27;
		22377: rom = 27;
		22378: rom = 24;
		22379: rom = 22;
		22380: rom = 20;
		22381: rom = 20;
		22382: rom = 22;
		22383: rom = 27;
		22384: rom = 27;
		22385: rom = 1;
		22386: rom = 0;
		22387: rom = 0;
		22388: rom = 0;
		22389: rom = 0;
		22390: rom = 19;
		22391: rom = 27;
		22392: rom = 27;
		22393: rom = 27;
		22394: rom = 27;
		22400: rom = 27;
		22401: rom = 27;
		22402: rom = 27;
		22403: rom = 27;
		22404: rom = 27;
		22405: rom = 27;
		22406: rom = 27;
		22407: rom = 27;
		22408: rom = 27;
		22409: rom = 27;
		22410: rom = 27;
		22411: rom = 27;
		22412: rom = 27;
		22413: rom = 27;
		22414: rom = 27;
		22415: rom = 27;
		22416: rom = 27;
		22417: rom = 27;
		22418: rom = 27;
		22419: rom = 27;
		22420: rom = 27;
		22421: rom = 27;
		22422: rom = 27;
		22423: rom = 27;
		22424: rom = 27;
		22425: rom = 27;
		22426: rom = 27;
		22427: rom = 27;
		22428: rom = 27;
		22429: rom = 27;
		22430: rom = 27;
		22431: rom = 27;
		22432: rom = 27;
		22433: rom = 27;
		22434: rom = 27;
		22435: rom = 27;
		22436: rom = 27;
		22437: rom = 27;
		22438: rom = 27;
		22439: rom = 27;
		22440: rom = 27;
		22441: rom = 27;
		22442: rom = 27;
		22443: rom = 27;
		22444: rom = 27;
		22445: rom = 27;
		22446: rom = 27;
		22447: rom = 27;
		22448: rom = 27;
		22449: rom = 27;
		22450: rom = 27;
		22451: rom = 22;
		22452: rom = 11;
		22453: rom = 7;
		22454: rom = 23;
		22455: rom = 11;
		22456: rom = 16;
		22457: rom = 17;
		22458: rom = 18;
		22459: rom = 22;
		22460: rom = 25;
		22461: rom = 23;
		22462: rom = 18;
		22463: rom = 18;
		22464: rom = 18;
		22465: rom = 18;
		22466: rom = 17;
		22467: rom = 15;
		22468: rom = 12;
		22469: rom = 12;
		22470: rom = 18;
		22471: rom = 23;
		22472: rom = 27;
		22473: rom = 27;
		22474: rom = 27;
		22475: rom = 27;
		22476: rom = 27;
		22477: rom = 0;
		22478: rom = 27;
		22479: rom = 27;
		22480: rom = 27;
		22481: rom = 27;
		22482: rom = 27;
		22483: rom = 27;
		22484: rom = 27;
		22485: rom = 27;
		22486: rom = 27;
		22487: rom = 27;
		22488: rom = 27;
		22489: rom = 27;
		22490: rom = 27;
		22491: rom = 27;
		22492: rom = 27;
		22493: rom = 27;
		22494: rom = 27;
		22495: rom = 27;
		22496: rom = 27;
		22497: rom = 27;
		22498: rom = 27;
		22499: rom = 27;
		22500: rom = 27;
		22501: rom = 27;
		22502: rom = 27;
		22503: rom = 27;
		22504: rom = 27;
		22505: rom = 27;
		22506: rom = 27;
		22507: rom = 27;
		22508: rom = 27;
		22509: rom = 27;
		22510: rom = 27;
		22511: rom = 27;
		22512: rom = 27;
		22513: rom = 24;
		22514: rom = 10;
		22515: rom = 0;
		22516: rom = 0;
		22517: rom = 0;
		22518: rom = 19;
		22519: rom = 27;
		22520: rom = 27;
		22521: rom = 27;
		22522: rom = 27;
		22528: rom = 27;
		22529: rom = 27;
		22530: rom = 27;
		22531: rom = 27;
		22532: rom = 27;
		22533: rom = 27;
		22534: rom = 27;
		22535: rom = 27;
		22536: rom = 27;
		22537: rom = 27;
		22538: rom = 27;
		22539: rom = 27;
		22540: rom = 27;
		22541: rom = 27;
		22542: rom = 27;
		22543: rom = 27;
		22544: rom = 27;
		22545: rom = 27;
		22546: rom = 27;
		22547: rom = 27;
		22548: rom = 27;
		22549: rom = 27;
		22550: rom = 27;
		22551: rom = 27;
		22552: rom = 27;
		22553: rom = 27;
		22554: rom = 27;
		22555: rom = 27;
		22556: rom = 27;
		22557: rom = 27;
		22558: rom = 27;
		22559: rom = 27;
		22560: rom = 27;
		22561: rom = 27;
		22562: rom = 27;
		22563: rom = 27;
		22564: rom = 27;
		22565: rom = 27;
		22566: rom = 27;
		22567: rom = 27;
		22568: rom = 27;
		22569: rom = 27;
		22570: rom = 27;
		22571: rom = 27;
		22572: rom = 27;
		22573: rom = 27;
		22574: rom = 27;
		22575: rom = 27;
		22576: rom = 27;
		22577: rom = 27;
		22578: rom = 27;
		22579: rom = 27;
		22580: rom = 26;
		22581: rom = 20;
		22582: rom = 26;
		22583: rom = 23;
		22584: rom = 19;
		22585: rom = 15;
		22586: rom = 11;
		22587: rom = 10;
		22588: rom = 16;
		22589: rom = 17;
		22590: rom = 12;
		22591: rom = 10;
		22592: rom = 11;
		22593: rom = 14;
		22594: rom = 18;
		22595: rom = 22;
		22596: rom = 25;
		22597: rom = 27;
		22598: rom = 27;
		22599: rom = 27;
		22600: rom = 27;
		22601: rom = 27;
		22602: rom = 27;
		22603: rom = 27;
		22604: rom = 27;
		22605: rom = 0;
		22606: rom = 0;
		22607: rom = 0;
		22608: rom = 0;
		22609: rom = 0;
		22610: rom = 27;
		22611: rom = 27;
		22612: rom = 27;
		22613: rom = 27;
		22614: rom = 27;
		22615: rom = 27;
		22616: rom = 27;
		22617: rom = 27;
		22618: rom = 27;
		22619: rom = 27;
		22620: rom = 27;
		22621: rom = 27;
		22622: rom = 27;
		22623: rom = 27;
		22624: rom = 27;
		22625: rom = 27;
		22626: rom = 27;
		22627: rom = 27;
		22628: rom = 27;
		22629: rom = 27;
		22630: rom = 27;
		22631: rom = 27;
		22632: rom = 27;
		22633: rom = 27;
		22634: rom = 27;
		22635: rom = 27;
		22636: rom = 27;
		22637: rom = 27;
		22638: rom = 27;
		22639: rom = 27;
		22640: rom = 27;
		22641: rom = 27;
		22642: rom = 27;
		22643: rom = 18;
		22644: rom = 0;
		22645: rom = 0;
		22646: rom = 19;
		22647: rom = 27;
		22648: rom = 27;
		22649: rom = 27;
		22650: rom = 27;
		22656: rom = 27;
		22657: rom = 27;
		22658: rom = 27;
		22659: rom = 27;
		22660: rom = 27;
		22661: rom = 27;
		22662: rom = 27;
		22663: rom = 27;
		22664: rom = 27;
		22665: rom = 27;
		22666: rom = 27;
		22667: rom = 27;
		22668: rom = 27;
		22669: rom = 27;
		22670: rom = 27;
		22671: rom = 27;
		22672: rom = 27;
		22673: rom = 27;
		22674: rom = 27;
		22675: rom = 27;
		22676: rom = 27;
		22677: rom = 27;
		22678: rom = 27;
		22679: rom = 27;
		22680: rom = 27;
		22681: rom = 27;
		22682: rom = 27;
		22683: rom = 27;
		22684: rom = 27;
		22685: rom = 27;
		22686: rom = 27;
		22687: rom = 27;
		22688: rom = 27;
		22689: rom = 27;
		22690: rom = 27;
		22691: rom = 27;
		22692: rom = 27;
		22693: rom = 27;
		22694: rom = 27;
		22695: rom = 27;
		22696: rom = 27;
		22697: rom = 27;
		22698: rom = 27;
		22699: rom = 27;
		22700: rom = 27;
		22701: rom = 27;
		22702: rom = 27;
		22703: rom = 27;
		22704: rom = 27;
		22705: rom = 27;
		22706: rom = 27;
		22707: rom = 27;
		22708: rom = 27;
		22709: rom = 27;
		22710: rom = 27;
		22711: rom = 27;
		22712: rom = 27;
		22713: rom = 27;
		22714: rom = 27;
		22715: rom = 27;
		22716: rom = 26;
		22717: rom = 26;
		22718: rom = 26;
		22719: rom = 27;
		22720: rom = 27;
		22721: rom = 27;
		22722: rom = 27;
		22723: rom = 27;
		22724: rom = 27;
		22725: rom = 27;
		22726: rom = 27;
		22727: rom = 27;
		22728: rom = 27;
		22729: rom = 27;
		22730: rom = 27;
		22731: rom = 27;
		22732: rom = 27;
		22733: rom = 0;
		22734: rom = 27;
		22735: rom = 27;
		22736: rom = 27;
		22737: rom = 27;
		22738: rom = 27;
		22739: rom = 27;
		22740: rom = 27;
		22741: rom = 27;
		22742: rom = 27;
		22743: rom = 27;
		22744: rom = 27;
		22745: rom = 27;
		22746: rom = 27;
		22747: rom = 27;
		22748: rom = 27;
		22749: rom = 27;
		22750: rom = 27;
		22751: rom = 27;
		22752: rom = 27;
		22753: rom = 27;
		22754: rom = 27;
		22755: rom = 27;
		22756: rom = 27;
		22757: rom = 27;
		22758: rom = 27;
		22759: rom = 27;
		22760: rom = 27;
		22761: rom = 27;
		22762: rom = 27;
		22763: rom = 27;
		22764: rom = 27;
		22765: rom = 27;
		22766: rom = 27;
		22767: rom = 27;
		22768: rom = 27;
		22769: rom = 27;
		22770: rom = 27;
		22771: rom = 27;
		22772: rom = 24;
		22773: rom = 10;
		22774: rom = 19;
		22775: rom = 27;
		22776: rom = 27;
		22777: rom = 27;
		22778: rom = 27;
		22784: rom = 27;
		22785: rom = 27;
		22786: rom = 27;
		22787: rom = 27;
		22788: rom = 27;
		22789: rom = 27;
		22790: rom = 27;
		22791: rom = 27;
		22792: rom = 27;
		22793: rom = 27;
		22794: rom = 27;
		22795: rom = 27;
		22796: rom = 27;
		22797: rom = 27;
		22798: rom = 27;
		22799: rom = 27;
		22800: rom = 27;
		22801: rom = 27;
		22802: rom = 27;
		22803: rom = 27;
		22804: rom = 27;
		22805: rom = 27;
		22806: rom = 27;
		22807: rom = 27;
		22808: rom = 27;
		22809: rom = 27;
		22810: rom = 27;
		22811: rom = 27;
		22812: rom = 27;
		22813: rom = 27;
		22814: rom = 27;
		22815: rom = 27;
		22816: rom = 27;
		22817: rom = 27;
		22818: rom = 27;
		22819: rom = 27;
		22820: rom = 27;
		22821: rom = 27;
		22822: rom = 27;
		22823: rom = 27;
		22824: rom = 27;
		22825: rom = 27;
		22826: rom = 27;
		22827: rom = 27;
		22828: rom = 27;
		22829: rom = 27;
		22830: rom = 27;
		22831: rom = 27;
		22832: rom = 27;
		22833: rom = 27;
		22834: rom = 27;
		22835: rom = 27;
		22836: rom = 27;
		22837: rom = 27;
		22838: rom = 27;
		22839: rom = 27;
		22840: rom = 27;
		22841: rom = 27;
		22842: rom = 27;
		22843: rom = 27;
		22844: rom = 27;
		22845: rom = 27;
		22846: rom = 27;
		22847: rom = 27;
		22848: rom = 27;
		22849: rom = 27;
		22850: rom = 27;
		22851: rom = 27;
		22852: rom = 27;
		22853: rom = 27;
		22854: rom = 27;
		22855: rom = 27;
		22856: rom = 27;
		22857: rom = 27;
		22858: rom = 27;
		22859: rom = 27;
		22860: rom = 27;
		22861: rom = 27;
		22862: rom = 27;
		22863: rom = 27;
		22864: rom = 27;
		22865: rom = 27;
		22866: rom = 27;
		22867: rom = 27;
		22868: rom = 27;
		22869: rom = 27;
		22870: rom = 27;
		22871: rom = 27;
		22872: rom = 27;
		22873: rom = 27;
		22874: rom = 27;
		22875: rom = 27;
		22876: rom = 27;
		22877: rom = 27;
		22878: rom = 27;
		22879: rom = 27;
		22880: rom = 27;
		22881: rom = 27;
		22882: rom = 27;
		22883: rom = 27;
		22884: rom = 27;
		22885: rom = 27;
		22886: rom = 27;
		22887: rom = 27;
		22888: rom = 27;
		22889: rom = 27;
		22890: rom = 27;
		22891: rom = 27;
		22892: rom = 27;
		22893: rom = 27;
		22894: rom = 27;
		22895: rom = 27;
		22896: rom = 27;
		22897: rom = 27;
		22898: rom = 27;
		22899: rom = 27;
		22900: rom = 27;
		22901: rom = 27;
		22902: rom = 27;
		22903: rom = 27;
		22904: rom = 0;
		22905: rom = 0;
		22906: rom = 27;
		22912: rom = 31;
		22913: rom = 31;
		22914: rom = 31;
		22915: rom = 31;
		22916: rom = 31;
		22917: rom = 31;
		22918: rom = 31;
		22919: rom = 31;
		22920: rom = 31;
		22921: rom = 31;
		22922: rom = 31;
		22923: rom = 31;
		22924: rom = 31;
		22925: rom = 31;
		22926: rom = 31;
		22927: rom = 31;
		22928: rom = 31;
		22929: rom = 31;
		22930: rom = 31;
		22931: rom = 31;
		22932: rom = 31;
		22933: rom = 31;
		22934: rom = 31;
		22935: rom = 31;
		22936: rom = 31;
		22937: rom = 31;
		22938: rom = 31;
		22939: rom = 31;
		22940: rom = 31;
		22941: rom = 31;
		22942: rom = 31;
		22943: rom = 31;
		22944: rom = 31;
		22945: rom = 31;
		22946: rom = 31;
		22947: rom = 31;
		22948: rom = 31;
		22949: rom = 31;
		22950: rom = 31;
		22951: rom = 31;
		22952: rom = 31;
		22953: rom = 31;
		22954: rom = 31;
		22955: rom = 31;
		22956: rom = 31;
		22957: rom = 31;
		22958: rom = 31;
		22959: rom = 31;
		22960: rom = 31;
		22961: rom = 31;
		22962: rom = 31;
		22963: rom = 31;
		22964: rom = 31;
		22965: rom = 31;
		22966: rom = 31;
		22967: rom = 31;
		22968: rom = 31;
		22969: rom = 31;
		22970: rom = 31;
		22971: rom = 31;
		22972: rom = 31;
		22973: rom = 31;
		22974: rom = 31;
		22975: rom = 31;
		22976: rom = 31;
		22977: rom = 31;
		22978: rom = 31;
		22979: rom = 31;
		22980: rom = 31;
		22981: rom = 31;
		22982: rom = 31;
		22983: rom = 31;
		22984: rom = 31;
		22985: rom = 31;
		22986: rom = 31;
		22987: rom = 31;
		22988: rom = 31;
		22989: rom = 0;
		22990: rom = 0;
		22991: rom = 0;
		22992: rom = 0;
		22993: rom = 0;
		22994: rom = 31;
		22995: rom = 31;
		22996: rom = 0;
		22997: rom = 31;
		22998: rom = 0;
		22999: rom = 31;
		23000: rom = 0;
		23001: rom = 31;
		23002: rom = 0;
		23003: rom = 31;
		23004: rom = 0;
		23005: rom = 31;
		23006: rom = 31;
		23007: rom = 0;
		23008: rom = 31;
		23009: rom = 0;
		23010: rom = 31;
		23011: rom = 0;
		23012: rom = 31;
		23013: rom = 0;
		23014: rom = 31;
		23015: rom = 31;
		23016: rom = 0;
		23017: rom = 0;
		23018: rom = 0;
		23019: rom = 0;
		23020: rom = 0;
		23021: rom = 0;
		23022: rom = 0;
		23023: rom = 31;
		23024: rom = 31;
		23025: rom = 31;
		23026: rom = 0;
		23027: rom = 31;
		23028: rom = 0;
		23029: rom = 31;
		23030: rom = 31;
		23031: rom = 0;
		23032: rom = 31;
		23033: rom = 0;
		23034: rom = 31;
		23040: rom = 31;
		23041: rom = 31;
		23042: rom = 31;
		23043: rom = 31;
		23044: rom = 31;
		23045: rom = 31;
		23046: rom = 31;
		23047: rom = 31;
		23048: rom = 31;
		23049: rom = 31;
		23050: rom = 31;
		23051: rom = 31;
		23052: rom = 31;
		23053: rom = 31;
		23054: rom = 31;
		23055: rom = 31;
		23056: rom = 31;
		23057: rom = 31;
		23058: rom = 31;
		23059: rom = 31;
		23060: rom = 31;
		23061: rom = 31;
		23062: rom = 31;
		23063: rom = 31;
		23064: rom = 31;
		23065: rom = 31;
		23066: rom = 31;
		23067: rom = 31;
		23068: rom = 31;
		23069: rom = 31;
		23070: rom = 31;
		23071: rom = 31;
		23072: rom = 31;
		23073: rom = 31;
		23074: rom = 31;
		23075: rom = 31;
		23076: rom = 31;
		23077: rom = 31;
		23078: rom = 31;
		23079: rom = 31;
		23080: rom = 31;
		23081: rom = 31;
		23082: rom = 31;
		23083: rom = 31;
		23084: rom = 31;
		23085: rom = 31;
		23086: rom = 31;
		23087: rom = 31;
		23088: rom = 31;
		23089: rom = 31;
		23090: rom = 31;
		23091: rom = 31;
		23092: rom = 31;
		23093: rom = 31;
		23094: rom = 31;
		23095: rom = 31;
		23096: rom = 31;
		23097: rom = 31;
		23098: rom = 31;
		23099: rom = 31;
		23100: rom = 31;
		23101: rom = 31;
		23102: rom = 31;
		23103: rom = 31;
		23104: rom = 31;
		23105: rom = 31;
		23106: rom = 31;
		23107: rom = 31;
		23108: rom = 31;
		23109: rom = 31;
		23110: rom = 31;
		23111: rom = 31;
		23112: rom = 31;
		23113: rom = 31;
		23114: rom = 31;
		23115: rom = 31;
		23116: rom = 31;
		23117: rom = 0;
		23118: rom = 31;
		23119: rom = 0;
		23120: rom = 31;
		23121: rom = 0;
		23122: rom = 31;
		23123: rom = 31;
		23124: rom = 31;
		23125: rom = 0;
		23126: rom = 31;
		23127: rom = 0;
		23128: rom = 31;
		23129: rom = 0;
		23130: rom = 31;
		23131: rom = 0;
		23132: rom = 31;
		23133: rom = 31;
		23134: rom = 31;
		23135: rom = 0;
		23136: rom = 31;
		23137: rom = 0;
		23138: rom = 31;
		23139: rom = 0;
		23140: rom = 31;
		23141: rom = 0;
		23142: rom = 31;
		23143: rom = 31;
		23144: rom = 31;
		23145: rom = 31;
		23146: rom = 31;
		23147: rom = 31;
		23148: rom = 31;
		23149: rom = 31;
		23150: rom = 31;
		23151: rom = 31;
		23152: rom = 31;
		23153: rom = 31;
		23154: rom = 31;
		23155: rom = 0;
		23156: rom = 31;
		23157: rom = 31;
		23158: rom = 0;
		23159: rom = 31;
		23160: rom = 31;
		23161: rom = 0;
		23162: rom = 31;
		23168: rom = 31;
		23169: rom = 31;
		23170: rom = 31;
		23171: rom = 31;
		23172: rom = 31;
		23173: rom = 31;
		23174: rom = 31;
		23175: rom = 31;
		23176: rom = 31;
		23177: rom = 31;
		23178: rom = 31;
		23179: rom = 31;
		23180: rom = 31;
		23181: rom = 31;
		23182: rom = 31;
		23183: rom = 31;
		23184: rom = 31;
		23185: rom = 31;
		23186: rom = 31;
		23187: rom = 31;
		23188: rom = 31;
		23189: rom = 31;
		23190: rom = 31;
		23191: rom = 31;
		23192: rom = 31;
		23193: rom = 31;
		23194: rom = 31;
		23195: rom = 31;
		23196: rom = 31;
		23197: rom = 31;
		23198: rom = 31;
		23199: rom = 31;
		23200: rom = 31;
		23201: rom = 31;
		23202: rom = 31;
		23203: rom = 31;
		23204: rom = 31;
		23205: rom = 31;
		23206: rom = 31;
		23207: rom = 31;
		23208: rom = 31;
		23209: rom = 31;
		23210: rom = 31;
		23211: rom = 31;
		23212: rom = 31;
		23213: rom = 31;
		23214: rom = 31;
		23215: rom = 31;
		23216: rom = 31;
		23217: rom = 31;
		23218: rom = 31;
		23219: rom = 31;
		23220: rom = 31;
		23221: rom = 31;
		23222: rom = 31;
		23223: rom = 31;
		23224: rom = 31;
		23225: rom = 31;
		23226: rom = 31;
		23227: rom = 31;
		23228: rom = 31;
		23229: rom = 31;
		23230: rom = 31;
		23231: rom = 31;
		23232: rom = 31;
		23233: rom = 31;
		23234: rom = 31;
		23235: rom = 31;
		23236: rom = 31;
		23237: rom = 31;
		23238: rom = 31;
		23239: rom = 31;
		23240: rom = 31;
		23241: rom = 31;
		23242: rom = 31;
		23243: rom = 31;
		23244: rom = 31;
		23245: rom = 31;
		23246: rom = 31;
		23247: rom = 31;
		23248: rom = 31;
		23249: rom = 31;
		23250: rom = 31;
		23251: rom = 31;
		23252: rom = 0;
		23253: rom = 31;
		23254: rom = 0;
		23255: rom = 31;
		23256: rom = 0;
		23257: rom = 31;
		23258: rom = 0;
		23259: rom = 31;
		23260: rom = 0;
		23261: rom = 31;
		23262: rom = 31;
		23263: rom = 0;
		23264: rom = 31;
		23265: rom = 0;
		23266: rom = 31;
		23267: rom = 0;
		23268: rom = 31;
		23269: rom = 0;
		23270: rom = 31;
		23271: rom = 31;
		23272: rom = 0;
		23273: rom = 0;
		23274: rom = 0;
		23275: rom = 0;
		23276: rom = 0;
		23277: rom = 0;
		23278: rom = 0;
		23279: rom = 31;
		23280: rom = 31;
		23281: rom = 31;
		23282: rom = 0;
		23283: rom = 31;
		23284: rom = 0;
		23285: rom = 31;
		23286: rom = 31;
		23287: rom = 0;
		23288: rom = 31;
		23289: rom = 0;
		23290: rom = 31;
		23296: rom = 31;
		23297: rom = 31;
		23298: rom = 31;
		23299: rom = 31;
		23300: rom = 31;
		23301: rom = 31;
		23302: rom = 31;
		23303: rom = 31;
		23304: rom = 31;
		23305: rom = 31;
		23306: rom = 31;
		23307: rom = 31;
		23308: rom = 31;
		23309: rom = 31;
		23310: rom = 31;
		23311: rom = 31;
		23312: rom = 31;
		23313: rom = 31;
		23314: rom = 31;
		23315: rom = 31;
		23316: rom = 31;
		23317: rom = 31;
		23318: rom = 31;
		23319: rom = 31;
		23320: rom = 31;
		23321: rom = 31;
		23322: rom = 31;
		23323: rom = 31;
		23324: rom = 31;
		23325: rom = 31;
		23326: rom = 31;
		23327: rom = 31;
		23328: rom = 31;
		23329: rom = 31;
		23330: rom = 31;
		23331: rom = 31;
		23332: rom = 31;
		23333: rom = 31;
		23334: rom = 31;
		23335: rom = 31;
		23336: rom = 31;
		23337: rom = 31;
		23338: rom = 31;
		23339: rom = 31;
		23340: rom = 31;
		23341: rom = 31;
		23342: rom = 31;
		23343: rom = 31;
		23344: rom = 31;
		23345: rom = 31;
		23346: rom = 31;
		23347: rom = 31;
		23348: rom = 31;
		23349: rom = 31;
		23350: rom = 31;
		23351: rom = 31;
		23352: rom = 31;
		23353: rom = 31;
		23354: rom = 31;
		23355: rom = 31;
		23356: rom = 31;
		23357: rom = 31;
		23358: rom = 31;
		23359: rom = 31;
		23360: rom = 31;
		23361: rom = 31;
		23362: rom = 31;
		23363: rom = 31;
		23364: rom = 31;
		23365: rom = 31;
		23366: rom = 31;
		23367: rom = 31;
		23368: rom = 31;
		23369: rom = 31;
		23370: rom = 31;
		23371: rom = 31;
		23372: rom = 31;
		23373: rom = 0;
		23374: rom = 0;
		23375: rom = 0;
		23376: rom = 31;
		23377: rom = 0;
		23378: rom = 31;
		23379: rom = 31;
		23380: rom = 31;
		23381: rom = 0;
		23382: rom = 31;
		23383: rom = 0;
		23384: rom = 31;
		23385: rom = 0;
		23386: rom = 31;
		23387: rom = 0;
		23388: rom = 31;
		23389: rom = 31;
		23390: rom = 31;
		23391: rom = 0;
		23392: rom = 31;
		23393: rom = 0;
		23394: rom = 31;
		23395: rom = 0;
		23396: rom = 31;
		23397: rom = 0;
		23398: rom = 31;
		23399: rom = 31;
		23400: rom = 31;
		23401: rom = 31;
		23402: rom = 31;
		23403: rom = 31;
		23404: rom = 31;
		23405: rom = 31;
		23406: rom = 31;
		23407: rom = 31;
		23408: rom = 31;
		23409: rom = 31;
		23410: rom = 31;
		23411: rom = 31;
		23412: rom = 31;
		23413: rom = 31;
		23414: rom = 31;
		23415: rom = 31;
		23416: rom = 0;
		23417: rom = 0;
		23418: rom = 31;
		23424: rom = 31;
		23425: rom = 31;
		23426: rom = 31;
		23427: rom = 31;
		23428: rom = 31;
		23429: rom = 31;
		23430: rom = 31;
		23431: rom = 31;
		23432: rom = 31;
		23433: rom = 31;
		23434: rom = 31;
		23435: rom = 31;
		23436: rom = 31;
		23437: rom = 31;
		23438: rom = 31;
		23439: rom = 31;
		23440: rom = 31;
		23441: rom = 31;
		23442: rom = 31;
		23443: rom = 31;
		23444: rom = 31;
		23445: rom = 31;
		23446: rom = 31;
		23447: rom = 31;
		23448: rom = 31;
		23449: rom = 31;
		23450: rom = 31;
		23451: rom = 31;
		23452: rom = 31;
		23453: rom = 31;
		23454: rom = 31;
		23455: rom = 31;
		23456: rom = 31;
		23457: rom = 31;
		23458: rom = 31;
		23459: rom = 31;
		23460: rom = 31;
		23461: rom = 31;
		23462: rom = 31;
		23463: rom = 31;
		23464: rom = 31;
		23465: rom = 31;
		23466: rom = 31;
		23467: rom = 31;
		23468: rom = 31;
		23469: rom = 31;
		23470: rom = 31;
		23471: rom = 31;
		23472: rom = 31;
		23473: rom = 31;
		23474: rom = 31;
		23475: rom = 31;
		23476: rom = 31;
		23477: rom = 31;
		23478: rom = 31;
		23479: rom = 31;
		23480: rom = 31;
		23481: rom = 31;
		23482: rom = 31;
		23483: rom = 31;
		23484: rom = 31;
		23485: rom = 31;
		23486: rom = 31;
		23487: rom = 31;
		23488: rom = 31;
		23489: rom = 31;
		23490: rom = 31;
		23491: rom = 31;
		23492: rom = 31;
		23493: rom = 31;
		23494: rom = 31;
		23495: rom = 31;
		23496: rom = 31;
		23497: rom = 31;
		23498: rom = 31;
		23499: rom = 31;
		23500: rom = 31;
		23501: rom = 0;
		23502: rom = 31;
		23503: rom = 0;
		23504: rom = 0;
		23505: rom = 0;
		23506: rom = 31;
		23507: rom = 31;
		23508: rom = 0;
		23509: rom = 31;
		23510: rom = 0;
		23511: rom = 31;
		23512: rom = 0;
		23513: rom = 31;
		23514: rom = 0;
		23515: rom = 31;
		23516: rom = 0;
		23517: rom = 31;
		23518: rom = 31;
		23519: rom = 0;
		23520: rom = 31;
		23521: rom = 0;
		23522: rom = 31;
		23523: rom = 0;
		23524: rom = 31;
		23525: rom = 0;
		23526: rom = 31;
		23527: rom = 31;
		23528: rom = 0;
		23529: rom = 0;
		23530: rom = 0;
		23531: rom = 0;
		23532: rom = 0;
		23533: rom = 0;
		23534: rom = 0;
		23535: rom = 31;
		23536: rom = 31;
		23537: rom = 31;
		23538: rom = 31;
		23539: rom = 0;
		23540: rom = 31;
		23541: rom = 31;
		23542: rom = 31;
		23543: rom = 31;
		23544: rom = 31;
		23545: rom = 31;
		23546: rom = 31;
		23552: rom = 31;
		23553: rom = 31;
		23554: rom = 31;
		23555: rom = 31;
		23556: rom = 31;
		23557: rom = 31;
		23558: rom = 31;
		23559: rom = 31;
		23560: rom = 31;
		23561: rom = 31;
		23562: rom = 31;
		23563: rom = 31;
		23564: rom = 31;
		23565: rom = 31;
		23566: rom = 31;
		23567: rom = 31;
		23568: rom = 31;
		23569: rom = 31;
		23570: rom = 31;
		23571: rom = 31;
		23572: rom = 31;
		23573: rom = 31;
		23574: rom = 31;
		23575: rom = 31;
		23576: rom = 31;
		23577: rom = 31;
		23578: rom = 31;
		23579: rom = 31;
		23580: rom = 31;
		23581: rom = 31;
		23582: rom = 31;
		23583: rom = 31;
		23584: rom = 31;
		23585: rom = 31;
		23586: rom = 31;
		23587: rom = 31;
		23588: rom = 31;
		23589: rom = 31;
		23590: rom = 31;
		23591: rom = 31;
		23592: rom = 31;
		23593: rom = 31;
		23594: rom = 31;
		23595: rom = 31;
		23596: rom = 31;
		23597: rom = 31;
		23598: rom = 31;
		23599: rom = 31;
		23600: rom = 31;
		23601: rom = 31;
		23602: rom = 31;
		23603: rom = 31;
		23604: rom = 31;
		23605: rom = 31;
		23606: rom = 31;
		23607: rom = 31;
		23608: rom = 31;
		23609: rom = 31;
		23610: rom = 31;
		23611: rom = 31;
		23612: rom = 31;
		23613: rom = 31;
		23614: rom = 31;
		23615: rom = 31;
		23616: rom = 31;
		23617: rom = 31;
		23618: rom = 31;
		23619: rom = 31;
		23620: rom = 31;
		23621: rom = 31;
		23622: rom = 31;
		23623: rom = 31;
		23624: rom = 31;
		23625: rom = 31;
		23626: rom = 31;
		23627: rom = 31;
		23628: rom = 31;
		23629: rom = 31;
		23630: rom = 31;
		23631: rom = 31;
		23632: rom = 31;
		23633: rom = 31;
		23634: rom = 31;
		23635: rom = 31;
		23636: rom = 31;
		23637: rom = 0;
		23638: rom = 31;
		23639: rom = 0;
		23640: rom = 31;
		23641: rom = 0;
		23642: rom = 31;
		23643: rom = 0;
		23644: rom = 31;
		23645: rom = 31;
		23646: rom = 31;
		23647: rom = 0;
		23648: rom = 31;
		23649: rom = 0;
		23650: rom = 31;
		23651: rom = 0;
		23652: rom = 31;
		23653: rom = 0;
		23654: rom = 31;
		23655: rom = 31;
		23656: rom = 31;
		23657: rom = 31;
		23658: rom = 31;
		23659: rom = 31;
		23660: rom = 31;
		23661: rom = 31;
		23662: rom = 31;
		23663: rom = 31;
		23664: rom = 31;
		23665: rom = 31;
		23666: rom = 0;
		23667: rom = 31;
		23668: rom = 0;
		23669: rom = 31;
		23670: rom = 31;
		23671: rom = 0;
		23672: rom = 0;
		23673: rom = 0;
		23674: rom = 31;
		23680: rom = 31;
		23681: rom = 31;
		23682: rom = 31;
		23683: rom = 31;
		23684: rom = 31;
		23685: rom = 31;
		23686: rom = 31;
		23687: rom = 31;
		23688: rom = 31;
		23689: rom = 31;
		23690: rom = 31;
		23691: rom = 31;
		23692: rom = 31;
		23693: rom = 31;
		23694: rom = 31;
		23695: rom = 31;
		23696: rom = 31;
		23697: rom = 31;
		23698: rom = 31;
		23699: rom = 31;
		23700: rom = 31;
		23701: rom = 31;
		23702: rom = 31;
		23703: rom = 31;
		23704: rom = 31;
		23705: rom = 31;
		23706: rom = 31;
		23707: rom = 31;
		23708: rom = 31;
		23709: rom = 31;
		23710: rom = 31;
		23711: rom = 31;
		23712: rom = 31;
		23713: rom = 31;
		23714: rom = 31;
		23715: rom = 31;
		23716: rom = 31;
		23717: rom = 31;
		23718: rom = 31;
		23719: rom = 31;
		23720: rom = 31;
		23721: rom = 31;
		23722: rom = 31;
		23723: rom = 31;
		23724: rom = 31;
		23725: rom = 31;
		23726: rom = 31;
		23727: rom = 31;
		23728: rom = 31;
		23729: rom = 31;
		23730: rom = 31;
		23731: rom = 31;
		23732: rom = 31;
		23733: rom = 31;
		23734: rom = 31;
		23735: rom = 31;
		23736: rom = 31;
		23737: rom = 31;
		23738: rom = 31;
		23739: rom = 31;
		23740: rom = 31;
		23741: rom = 31;
		23742: rom = 31;
		23743: rom = 31;
		23744: rom = 31;
		23745: rom = 31;
		23746: rom = 31;
		23747: rom = 31;
		23748: rom = 31;
		23749: rom = 31;
		23750: rom = 31;
		23751: rom = 31;
		23752: rom = 31;
		23753: rom = 31;
		23754: rom = 31;
		23755: rom = 31;
		23756: rom = 31;
		23757: rom = 0;
		23758: rom = 31;
		23759: rom = 31;
		23760: rom = 31;
		23761: rom = 31;
		23762: rom = 31;
		23763: rom = 31;
		23764: rom = 0;
		23765: rom = 31;
		23766: rom = 0;
		23767: rom = 31;
		23768: rom = 0;
		23769: rom = 31;
		23770: rom = 0;
		23771: rom = 31;
		23772: rom = 0;
		23773: rom = 31;
		23774: rom = 31;
		23775: rom = 0;
		23776: rom = 31;
		23777: rom = 0;
		23778: rom = 31;
		23779: rom = 0;
		23780: rom = 31;
		23781: rom = 0;
		23782: rom = 31;
		23783: rom = 31;
		23784: rom = 0;
		23785: rom = 0;
		23786: rom = 0;
		23787: rom = 0;
		23788: rom = 0;
		23789: rom = 0;
		23790: rom = 0;
		23791: rom = 31;
		23792: rom = 31;
		23793: rom = 31;
		23794: rom = 31;
		23795: rom = 0;
		23796: rom = 31;
		23797: rom = 31;
		23798: rom = 0;
		23799: rom = 31;
		23800: rom = 0;
		23801: rom = 31;
		23802: rom = 31;
		23808: rom = 31;
		23809: rom = 31;
		23810: rom = 31;
		23811: rom = 31;
		23812: rom = 31;
		23813: rom = 31;
		23814: rom = 31;
		23815: rom = 31;
		23816: rom = 31;
		23817: rom = 31;
		23818: rom = 31;
		23819: rom = 31;
		23820: rom = 31;
		23821: rom = 31;
		23822: rom = 31;
		23823: rom = 31;
		23824: rom = 31;
		23825: rom = 31;
		23826: rom = 31;
		23827: rom = 31;
		23828: rom = 31;
		23829: rom = 31;
		23830: rom = 31;
		23831: rom = 31;
		23832: rom = 31;
		23833: rom = 31;
		23834: rom = 31;
		23835: rom = 31;
		23836: rom = 31;
		23837: rom = 31;
		23838: rom = 31;
		23839: rom = 31;
		23840: rom = 31;
		23841: rom = 31;
		23842: rom = 31;
		23843: rom = 31;
		23844: rom = 31;
		23845: rom = 31;
		23846: rom = 31;
		23847: rom = 31;
		23848: rom = 31;
		23849: rom = 31;
		23850: rom = 31;
		23851: rom = 31;
		23852: rom = 31;
		23853: rom = 31;
		23854: rom = 31;
		23855: rom = 31;
		23856: rom = 31;
		23857: rom = 31;
		23858: rom = 31;
		23859: rom = 31;
		23860: rom = 31;
		23861: rom = 31;
		23862: rom = 31;
		23863: rom = 31;
		23864: rom = 31;
		23865: rom = 31;
		23866: rom = 31;
		23867: rom = 31;
		23868: rom = 31;
		23869: rom = 31;
		23870: rom = 31;
		23871: rom = 31;
		23872: rom = 31;
		23873: rom = 31;
		23874: rom = 31;
		23875: rom = 31;
		23876: rom = 31;
		23877: rom = 31;
		23878: rom = 31;
		23879: rom = 31;
		23880: rom = 31;
		23881: rom = 31;
		23882: rom = 31;
		23883: rom = 31;
		23884: rom = 31;
		23885: rom = 0;
		23886: rom = 0;
		23887: rom = 0;
		23888: rom = 0;
		23889: rom = 0;
		23890: rom = 31;
		23891: rom = 31;
		23892: rom = 31;
		23893: rom = 0;
		23894: rom = 31;
		23895: rom = 0;
		23896: rom = 31;
		23897: rom = 0;
		23898: rom = 31;
		23899: rom = 0;
		23900: rom = 31;
		23901: rom = 31;
		23902: rom = 31;
		23903: rom = 0;
		23904: rom = 31;
		23905: rom = 0;
		23906: rom = 31;
		23907: rom = 0;
		23908: rom = 31;
		23909: rom = 0;
		23910: rom = 31;
		23911: rom = 31;
		23912: rom = 31;
		23913: rom = 31;
		23914: rom = 31;
		23915: rom = 31;
		23916: rom = 31;
		23917: rom = 31;
		23918: rom = 31;
		23919: rom = 31;
		23920: rom = 31;
		23921: rom = 31;
		23922: rom = 31;
		23923: rom = 31;
		23924: rom = 31;
		23925: rom = 31;
		23926: rom = 31;
		23927: rom = 0;
		23928: rom = 0;
		23929: rom = 0;
		23930: rom = 31;
		23936: rom = 31;
		23937: rom = 31;
		23938: rom = 31;
		23939: rom = 31;
		23940: rom = 31;
		23941: rom = 31;
		23942: rom = 31;
		23943: rom = 31;
		23944: rom = 31;
		23945: rom = 31;
		23946: rom = 31;
		23947: rom = 31;
		23948: rom = 31;
		23949: rom = 31;
		23950: rom = 31;
		23951: rom = 31;
		23952: rom = 31;
		23953: rom = 31;
		23954: rom = 31;
		23955: rom = 31;
		23956: rom = 31;
		23957: rom = 31;
		23958: rom = 31;
		23959: rom = 31;
		23960: rom = 31;
		23961: rom = 31;
		23962: rom = 31;
		23963: rom = 31;
		23964: rom = 31;
		23965: rom = 31;
		23966: rom = 31;
		23967: rom = 31;
		23968: rom = 31;
		23969: rom = 31;
		23970: rom = 31;
		23971: rom = 31;
		23972: rom = 31;
		23973: rom = 31;
		23974: rom = 31;
		23975: rom = 31;
		23976: rom = 31;
		23977: rom = 31;
		23978: rom = 31;
		23979: rom = 31;
		23980: rom = 31;
		23981: rom = 31;
		23982: rom = 31;
		23983: rom = 31;
		23984: rom = 31;
		23985: rom = 31;
		23986: rom = 31;
		23987: rom = 31;
		23988: rom = 31;
		23989: rom = 31;
		23990: rom = 31;
		23991: rom = 31;
		23992: rom = 31;
		23993: rom = 31;
		23994: rom = 31;
		23995: rom = 31;
		23996: rom = 31;
		23997: rom = 31;
		23998: rom = 31;
		23999: rom = 31;
		24000: rom = 31;
		24001: rom = 31;
		24002: rom = 31;
		24003: rom = 31;
		24004: rom = 31;
		24005: rom = 31;
		24006: rom = 31;
		24007: rom = 31;
		24008: rom = 31;
		24009: rom = 31;
		24010: rom = 31;
		24011: rom = 31;
		24012: rom = 31;
		24013: rom = 0;
		24014: rom = 31;
		24015: rom = 31;
		24016: rom = 31;
		24017: rom = 31;
		24018: rom = 31;
		24019: rom = 31;
		24020: rom = 0;
		24021: rom = 31;
		24022: rom = 0;
		24023: rom = 31;
		24024: rom = 0;
		24025: rom = 31;
		24026: rom = 0;
		24027: rom = 31;
		24028: rom = 0;
		24029: rom = 31;
		24030: rom = 31;
		24031: rom = 0;
		24032: rom = 31;
		24033: rom = 0;
		24034: rom = 31;
		24035: rom = 0;
		24036: rom = 31;
		24037: rom = 0;
		24038: rom = 31;
		24039: rom = 31;
		24040: rom = 0;
		24041: rom = 0;
		24042: rom = 0;
		24043: rom = 0;
		24044: rom = 0;
		24045: rom = 0;
		24046: rom = 0;
		24047: rom = 31;
		24048: rom = 31;
		24049: rom = 31;
		24050: rom = 31;
		24051: rom = 31;
		24052: rom = 31;
		24053: rom = 31;
		24054: rom = 31;
		24055: rom = 31;
		24056: rom = 31;
		24057: rom = 31;
		24058: rom = 31;
	endcase
end

endmodule
