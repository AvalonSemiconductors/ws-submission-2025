module avali_logo;
endmodule
