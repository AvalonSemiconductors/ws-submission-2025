VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__asig_5p0_fixed
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_fd_io__asig_5p0_fixed ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN ASIG5V
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1200.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.020 349.000 23.560 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 26.700 349.000 29.240 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 32.380 349.000 34.920 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 40.080 349.000 42.620 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 45.760 349.000 48.300 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 51.440 349.000 53.980 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 57.120 349.000 59.660 350.000 ;
    END
  END ASIG5V
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -0.160 65.540 0.000 349.785 ;
        RECT 75.000 65.540 75.160 349.785 ;
      LAYER Metal5 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1200.000000 ;
    PORT
      LAYER Metal5 ;
        RECT 25.000 20.000 50.000 45.000 ;
    END
  END PAD
  OBS
      LAYER Pwell ;
        RECT 3.790 329.755 19.670 344.755 ;
        RECT 20.970 329.755 36.850 344.755 ;
        RECT 38.150 329.755 54.030 344.755 ;
        RECT 55.330 329.755 71.210 344.755 ;
        RECT 3.790 310.015 19.670 325.015 ;
        RECT 20.970 310.015 36.850 325.015 ;
        RECT 38.150 310.015 54.030 325.015 ;
        RECT 55.330 310.015 71.210 325.015 ;
        RECT 3.790 290.275 19.670 305.275 ;
        RECT 20.970 290.275 36.850 305.275 ;
        RECT 38.150 290.275 54.030 305.275 ;
        RECT 55.330 290.275 71.210 305.275 ;
        RECT 3.790 270.535 19.670 285.535 ;
        RECT 20.970 270.535 36.850 285.535 ;
        RECT 38.150 270.535 54.030 285.535 ;
        RECT 55.330 270.535 71.210 285.535 ;
        RECT 3.790 250.795 19.670 265.795 ;
        RECT 20.970 250.795 36.850 265.795 ;
        RECT 38.150 250.795 54.030 265.795 ;
        RECT 55.330 250.795 71.210 265.795 ;
        RECT 3.790 231.055 19.670 246.055 ;
        RECT 20.970 231.055 36.850 246.055 ;
        RECT 38.150 231.055 54.030 246.055 ;
        RECT 55.330 231.055 71.210 246.055 ;
        RECT 3.790 211.315 19.670 226.315 ;
        RECT 20.970 211.315 36.850 226.315 ;
        RECT 38.150 211.315 54.030 226.315 ;
        RECT 55.330 211.315 71.210 226.315 ;
        RECT 3.790 191.575 19.670 206.575 ;
        RECT 20.970 191.575 36.850 206.575 ;
        RECT 38.150 191.575 54.030 206.575 ;
        RECT 55.330 191.575 71.210 206.575 ;
        RECT 3.790 171.835 19.670 186.835 ;
        RECT 20.970 171.835 36.850 186.835 ;
        RECT 38.150 171.835 54.030 186.835 ;
        RECT 55.330 171.835 71.210 186.835 ;
      LAYER Nwell ;
        RECT 11.840 164.355 63.160 167.135 ;
        RECT 11.840 144.635 14.620 164.355 ;
        RECT 60.380 144.635 63.160 164.355 ;
        RECT 11.840 141.855 63.160 144.635 ;
        RECT 6.590 137.080 68.410 140.360 ;
        RECT 6.590 107.860 9.870 137.080 ;
        RECT 65.130 107.860 68.410 137.080 ;
        RECT 6.590 104.580 68.410 107.860 ;
        RECT 9.850 70.755 65.150 100.115 ;
      LAYER Metal1 ;
        RECT 0.000 348.945 75.000 349.785 ;
        RECT 0.000 165.355 0.450 348.945 ;
        RECT 1.780 345.505 73.220 347.295 ;
        RECT 1.780 329.005 2.120 345.505 ;
        RECT 4.440 344.865 19.020 345.205 ;
        RECT 3.140 329.005 4.140 344.755 ;
        RECT 4.440 329.645 9.440 344.865 ;
        RECT 14.020 329.645 19.020 344.865 ;
        RECT 21.620 344.865 36.200 345.205 ;
        RECT 4.440 329.305 19.020 329.645 ;
        RECT 19.320 329.005 21.320 344.755 ;
        RECT 21.620 329.645 26.620 344.865 ;
        RECT 31.200 329.645 36.200 344.865 ;
        RECT 38.800 344.865 53.380 345.205 ;
        RECT 21.620 329.305 36.200 329.645 ;
        RECT 36.500 329.005 38.500 344.755 ;
        RECT 38.800 329.645 43.800 344.865 ;
        RECT 48.380 329.645 53.380 344.865 ;
        RECT 55.980 344.865 70.560 345.205 ;
        RECT 38.800 329.305 53.380 329.645 ;
        RECT 53.680 329.005 55.680 344.755 ;
        RECT 55.980 329.645 60.980 344.865 ;
        RECT 65.560 329.645 70.560 344.865 ;
        RECT 55.980 329.305 70.560 329.645 ;
        RECT 70.860 329.005 71.860 344.755 ;
        RECT 72.880 329.005 73.220 345.505 ;
        RECT 1.780 325.765 73.220 329.005 ;
        RECT 1.780 309.265 2.120 325.765 ;
        RECT 4.440 325.125 19.020 325.465 ;
        RECT 3.140 309.265 4.140 325.015 ;
        RECT 4.440 309.905 9.440 325.125 ;
        RECT 14.020 309.905 19.020 325.125 ;
        RECT 21.620 325.125 36.200 325.465 ;
        RECT 4.440 309.565 19.020 309.905 ;
        RECT 19.320 309.265 21.320 325.015 ;
        RECT 21.620 309.905 26.620 325.125 ;
        RECT 31.200 309.905 36.200 325.125 ;
        RECT 38.800 325.125 53.380 325.465 ;
        RECT 21.620 309.565 36.200 309.905 ;
        RECT 36.500 309.265 38.500 325.015 ;
        RECT 38.800 309.905 43.800 325.125 ;
        RECT 48.380 309.905 53.380 325.125 ;
        RECT 55.980 325.125 70.560 325.465 ;
        RECT 38.800 309.565 53.380 309.905 ;
        RECT 53.680 309.265 55.680 325.015 ;
        RECT 55.980 309.905 60.980 325.125 ;
        RECT 65.560 309.905 70.560 325.125 ;
        RECT 55.980 309.565 70.560 309.905 ;
        RECT 70.860 309.265 71.860 325.015 ;
        RECT 72.880 309.265 73.220 325.765 ;
        RECT 1.780 306.025 73.220 309.265 ;
        RECT 1.780 289.525 2.120 306.025 ;
        RECT 4.440 305.385 19.020 305.725 ;
        RECT 3.140 289.525 4.140 305.275 ;
        RECT 4.440 290.165 9.440 305.385 ;
        RECT 14.020 290.165 19.020 305.385 ;
        RECT 21.620 305.385 36.200 305.725 ;
        RECT 4.440 289.825 19.020 290.165 ;
        RECT 19.320 289.525 21.320 305.275 ;
        RECT 21.620 290.165 26.620 305.385 ;
        RECT 31.200 290.165 36.200 305.385 ;
        RECT 38.800 305.385 53.380 305.725 ;
        RECT 21.620 289.825 36.200 290.165 ;
        RECT 36.500 289.525 38.500 305.275 ;
        RECT 38.800 290.165 43.800 305.385 ;
        RECT 48.380 290.165 53.380 305.385 ;
        RECT 55.980 305.385 70.560 305.725 ;
        RECT 38.800 289.825 53.380 290.165 ;
        RECT 53.680 289.525 55.680 305.275 ;
        RECT 55.980 290.165 60.980 305.385 ;
        RECT 65.560 290.165 70.560 305.385 ;
        RECT 55.980 289.825 70.560 290.165 ;
        RECT 70.860 289.525 71.860 305.275 ;
        RECT 72.880 289.525 73.220 306.025 ;
        RECT 1.780 286.285 73.220 289.525 ;
        RECT 1.780 269.785 2.120 286.285 ;
        RECT 4.440 285.645 19.020 285.985 ;
        RECT 3.140 269.785 4.140 285.535 ;
        RECT 4.440 270.425 9.440 285.645 ;
        RECT 14.020 270.425 19.020 285.645 ;
        RECT 21.620 285.645 36.200 285.985 ;
        RECT 4.440 270.085 19.020 270.425 ;
        RECT 19.320 269.785 21.320 285.535 ;
        RECT 21.620 270.425 26.620 285.645 ;
        RECT 31.200 270.425 36.200 285.645 ;
        RECT 38.800 285.645 53.380 285.985 ;
        RECT 21.620 270.085 36.200 270.425 ;
        RECT 36.500 269.785 38.500 285.535 ;
        RECT 38.800 270.425 43.800 285.645 ;
        RECT 48.380 270.425 53.380 285.645 ;
        RECT 55.980 285.645 70.560 285.985 ;
        RECT 38.800 270.085 53.380 270.425 ;
        RECT 53.680 269.785 55.680 285.535 ;
        RECT 55.980 270.425 60.980 285.645 ;
        RECT 65.560 270.425 70.560 285.645 ;
        RECT 55.980 270.085 70.560 270.425 ;
        RECT 70.860 269.785 71.860 285.535 ;
        RECT 72.880 269.785 73.220 286.285 ;
        RECT 1.780 266.545 73.220 269.785 ;
        RECT 1.780 250.045 2.120 266.545 ;
        RECT 4.440 265.905 19.020 266.245 ;
        RECT 3.140 250.045 4.140 265.795 ;
        RECT 4.440 250.685 9.440 265.905 ;
        RECT 14.020 250.685 19.020 265.905 ;
        RECT 21.620 265.905 36.200 266.245 ;
        RECT 4.440 250.345 19.020 250.685 ;
        RECT 19.320 250.045 21.320 265.795 ;
        RECT 21.620 250.685 26.620 265.905 ;
        RECT 31.200 250.685 36.200 265.905 ;
        RECT 38.800 265.905 53.380 266.245 ;
        RECT 21.620 250.345 36.200 250.685 ;
        RECT 36.500 250.045 38.500 265.795 ;
        RECT 38.800 250.685 43.800 265.905 ;
        RECT 48.380 250.685 53.380 265.905 ;
        RECT 55.980 265.905 70.560 266.245 ;
        RECT 38.800 250.345 53.380 250.685 ;
        RECT 53.680 250.045 55.680 265.795 ;
        RECT 55.980 250.685 60.980 265.905 ;
        RECT 65.560 250.685 70.560 265.905 ;
        RECT 55.980 250.345 70.560 250.685 ;
        RECT 70.860 250.045 71.860 265.795 ;
        RECT 72.880 250.045 73.220 266.545 ;
        RECT 1.780 246.805 73.220 250.045 ;
        RECT 1.780 230.305 2.120 246.805 ;
        RECT 4.440 246.165 19.020 246.505 ;
        RECT 3.140 230.305 4.140 246.055 ;
        RECT 4.440 230.945 9.440 246.165 ;
        RECT 14.020 230.945 19.020 246.165 ;
        RECT 21.620 246.165 36.200 246.505 ;
        RECT 4.440 230.605 19.020 230.945 ;
        RECT 19.320 230.305 21.320 246.055 ;
        RECT 21.620 230.945 26.620 246.165 ;
        RECT 31.200 230.945 36.200 246.165 ;
        RECT 38.800 246.165 53.380 246.505 ;
        RECT 21.620 230.605 36.200 230.945 ;
        RECT 36.500 230.305 38.500 246.055 ;
        RECT 38.800 230.945 43.800 246.165 ;
        RECT 48.380 230.945 53.380 246.165 ;
        RECT 55.980 246.165 70.560 246.505 ;
        RECT 38.800 230.605 53.380 230.945 ;
        RECT 53.680 230.305 55.680 246.055 ;
        RECT 55.980 230.945 60.980 246.165 ;
        RECT 65.560 230.945 70.560 246.165 ;
        RECT 55.980 230.605 70.560 230.945 ;
        RECT 70.860 230.305 71.860 246.055 ;
        RECT 72.880 230.305 73.220 246.805 ;
        RECT 1.780 227.065 73.220 230.305 ;
        RECT 1.780 210.565 2.120 227.065 ;
        RECT 4.440 226.425 19.020 226.765 ;
        RECT 3.140 210.565 4.140 226.315 ;
        RECT 4.440 211.205 9.440 226.425 ;
        RECT 14.020 211.205 19.020 226.425 ;
        RECT 21.620 226.425 36.200 226.765 ;
        RECT 4.440 210.865 19.020 211.205 ;
        RECT 19.320 210.565 21.320 226.315 ;
        RECT 21.620 211.205 26.620 226.425 ;
        RECT 31.200 211.205 36.200 226.425 ;
        RECT 38.800 226.425 53.380 226.765 ;
        RECT 21.620 210.865 36.200 211.205 ;
        RECT 36.500 210.565 38.500 226.315 ;
        RECT 38.800 211.205 43.800 226.425 ;
        RECT 48.380 211.205 53.380 226.425 ;
        RECT 55.980 226.425 70.560 226.765 ;
        RECT 38.800 210.865 53.380 211.205 ;
        RECT 53.680 210.565 55.680 226.315 ;
        RECT 55.980 211.205 60.980 226.425 ;
        RECT 65.560 211.205 70.560 226.425 ;
        RECT 55.980 210.865 70.560 211.205 ;
        RECT 70.860 210.565 71.860 226.315 ;
        RECT 72.880 210.565 73.220 227.065 ;
        RECT 1.780 207.325 73.220 210.565 ;
        RECT 1.780 190.825 2.120 207.325 ;
        RECT 4.440 206.685 19.020 207.025 ;
        RECT 3.140 190.825 4.140 206.575 ;
        RECT 4.440 191.465 9.440 206.685 ;
        RECT 14.020 191.465 19.020 206.685 ;
        RECT 21.620 206.685 36.200 207.025 ;
        RECT 4.440 191.125 19.020 191.465 ;
        RECT 19.320 190.825 21.320 206.575 ;
        RECT 21.620 191.465 26.620 206.685 ;
        RECT 31.200 191.465 36.200 206.685 ;
        RECT 38.800 206.685 53.380 207.025 ;
        RECT 21.620 191.125 36.200 191.465 ;
        RECT 36.500 190.825 38.500 206.575 ;
        RECT 38.800 191.465 43.800 206.685 ;
        RECT 48.380 191.465 53.380 206.685 ;
        RECT 55.980 206.685 70.560 207.025 ;
        RECT 38.800 191.125 53.380 191.465 ;
        RECT 53.680 190.825 55.680 206.575 ;
        RECT 55.980 191.465 60.980 206.685 ;
        RECT 65.560 191.465 70.560 206.685 ;
        RECT 55.980 191.125 70.560 191.465 ;
        RECT 70.860 190.825 71.860 206.575 ;
        RECT 72.880 190.825 73.220 207.325 ;
        RECT 1.780 187.585 73.220 190.825 ;
        RECT 1.780 171.085 2.120 187.585 ;
        RECT 4.440 186.945 19.020 187.285 ;
        RECT 3.140 171.085 4.140 186.835 ;
        RECT 4.440 171.725 9.440 186.945 ;
        RECT 14.020 171.725 19.020 186.945 ;
        RECT 21.620 186.945 36.200 187.285 ;
        RECT 4.440 171.385 19.020 171.725 ;
        RECT 19.320 171.085 21.320 186.835 ;
        RECT 21.620 171.725 26.620 186.945 ;
        RECT 31.200 171.725 36.200 186.945 ;
        RECT 38.800 186.945 53.380 187.285 ;
        RECT 21.620 171.385 36.200 171.725 ;
        RECT 36.500 171.085 38.500 186.835 ;
        RECT 38.800 171.725 43.800 186.945 ;
        RECT 48.380 171.725 53.380 186.945 ;
        RECT 55.980 186.945 70.560 187.285 ;
        RECT 38.800 171.385 53.380 171.725 ;
        RECT 53.680 171.085 55.680 186.835 ;
        RECT 55.980 171.725 60.980 186.945 ;
        RECT 65.560 171.725 70.560 186.945 ;
        RECT 55.980 171.385 70.560 171.725 ;
        RECT 70.860 171.085 71.860 186.835 ;
        RECT 72.880 171.085 73.220 187.585 ;
        RECT 1.780 169.295 73.220 171.085 ;
        RECT 0.000 160.355 5.180 165.355 ;
        RECT 0.000 159.355 0.450 160.355 ;
        RECT 1.340 159.355 5.180 160.355 ;
        RECT 0.000 154.355 5.180 159.355 ;
        RECT 0.000 153.355 0.450 154.355 ;
        RECT 1.340 153.355 5.180 154.355 ;
        RECT 0.000 148.355 5.180 153.355 ;
        RECT 0.000 147.355 0.450 148.355 ;
        RECT 1.340 147.355 5.180 148.355 ;
        RECT 0.000 142.355 5.180 147.355 ;
        RECT 0.000 141.355 0.450 142.355 ;
        RECT 1.340 141.355 5.180 142.355 ;
        RECT 12.310 164.825 62.690 166.665 ;
        RECT 74.550 165.355 75.000 348.945 ;
        RECT 12.310 144.165 14.150 164.825 ;
        RECT 15.475 162.315 59.525 163.425 ;
        RECT 15.475 159.795 16.585 162.315 ;
        RECT 17.500 160.535 57.500 161.535 ;
        RECT 58.415 159.795 59.525 162.315 ;
        RECT 15.475 157.915 59.525 159.795 ;
        RECT 15.475 155.435 16.585 157.915 ;
        RECT 17.500 156.175 57.500 157.175 ;
        RECT 58.415 155.435 59.525 157.915 ;
        RECT 15.475 153.555 59.525 155.435 ;
        RECT 15.475 151.075 16.585 153.555 ;
        RECT 17.500 151.815 57.500 152.815 ;
        RECT 58.415 151.075 59.525 153.555 ;
        RECT 15.475 149.195 59.525 151.075 ;
        RECT 15.475 146.675 16.585 149.195 ;
        RECT 17.500 147.455 57.500 148.455 ;
        RECT 58.415 146.675 59.525 149.195 ;
        RECT 15.475 145.565 59.525 146.675 ;
        RECT 60.850 144.165 62.690 164.825 ;
        RECT 12.310 142.325 62.690 144.165 ;
        RECT 69.820 160.355 75.000 165.355 ;
        RECT 69.820 159.355 73.660 160.355 ;
        RECT 74.550 159.355 75.000 160.355 ;
        RECT 69.820 154.355 75.000 159.355 ;
        RECT 69.820 153.355 73.660 154.355 ;
        RECT 74.550 153.355 75.000 154.355 ;
        RECT 69.820 148.355 75.000 153.355 ;
        RECT 69.820 147.355 73.660 148.355 ;
        RECT 74.550 147.355 75.000 148.355 ;
        RECT 69.820 142.355 75.000 147.355 ;
        RECT 0.000 136.355 5.180 141.355 ;
        RECT 69.820 141.355 73.660 142.355 ;
        RECT 74.550 141.355 75.000 142.355 ;
        RECT 0.000 135.355 0.450 136.355 ;
        RECT 1.340 135.355 5.180 136.355 ;
        RECT 0.000 130.355 5.180 135.355 ;
        RECT 0.000 129.355 0.450 130.355 ;
        RECT 1.340 129.355 5.180 130.355 ;
        RECT 0.000 124.355 5.180 129.355 ;
        RECT 0.000 123.355 0.450 124.355 ;
        RECT 1.340 123.355 5.180 124.355 ;
        RECT 0.000 118.355 5.180 123.355 ;
        RECT 0.000 117.355 0.450 118.355 ;
        RECT 1.340 117.355 5.180 118.355 ;
        RECT 0.000 112.355 5.180 117.355 ;
        RECT 0.000 109.015 0.450 112.355 ;
        RECT 1.340 109.015 5.180 112.355 ;
        RECT 0.000 104.015 5.180 109.015 ;
        RECT 7.060 137.550 67.940 139.890 ;
        RECT 7.060 107.390 9.400 137.550 ;
        RECT 10.320 135.570 64.680 136.680 ;
        RECT 10.320 130.430 11.430 135.570 ;
        RECT 12.500 131.500 62.500 134.500 ;
        RECT 63.570 130.430 64.680 135.570 ;
        RECT 10.320 128.550 64.680 130.430 ;
        RECT 10.320 123.410 11.430 128.550 ;
        RECT 12.500 124.480 62.500 127.480 ;
        RECT 63.570 123.410 64.680 128.550 ;
        RECT 10.320 121.530 64.680 123.410 ;
        RECT 10.320 116.390 11.430 121.530 ;
        RECT 12.500 117.460 62.500 120.460 ;
        RECT 63.570 116.390 64.680 121.530 ;
        RECT 10.320 114.510 64.680 116.390 ;
        RECT 10.320 109.370 11.430 114.510 ;
        RECT 12.500 110.440 62.500 113.440 ;
        RECT 63.570 109.370 64.680 114.510 ;
        RECT 10.320 108.260 64.680 109.370 ;
        RECT 65.600 107.390 67.940 137.550 ;
        RECT 7.060 105.050 67.940 107.390 ;
        RECT 69.820 136.355 75.000 141.355 ;
        RECT 69.820 135.355 73.660 136.355 ;
        RECT 74.550 135.355 75.000 136.355 ;
        RECT 69.820 130.355 75.000 135.355 ;
        RECT 69.820 129.355 73.660 130.355 ;
        RECT 74.550 129.355 75.000 130.355 ;
        RECT 69.820 124.355 75.000 129.355 ;
        RECT 69.820 123.355 73.660 124.355 ;
        RECT 74.550 123.355 75.000 124.355 ;
        RECT 69.820 118.355 75.000 123.355 ;
        RECT 69.820 117.355 73.660 118.355 ;
        RECT 74.550 117.355 75.000 118.355 ;
        RECT 69.820 112.355 75.000 117.355 ;
        RECT 69.820 109.015 73.660 112.355 ;
        RECT 74.550 109.015 75.000 112.355 ;
        RECT 0.000 103.015 0.450 104.015 ;
        RECT 1.340 103.015 5.180 104.015 ;
        RECT 0.000 98.015 5.180 103.015 ;
        RECT 69.820 104.015 75.000 109.015 ;
        RECT 69.820 103.015 73.660 104.015 ;
        RECT 74.550 103.015 75.000 104.015 ;
        RECT 0.000 97.015 0.450 98.015 ;
        RECT 1.340 97.015 5.180 98.015 ;
        RECT 0.000 92.015 5.180 97.015 ;
        RECT 0.000 91.015 0.450 92.015 ;
        RECT 1.340 91.015 5.180 92.015 ;
        RECT 0.000 86.015 5.180 91.015 ;
        RECT 0.000 85.015 0.450 86.015 ;
        RECT 1.340 85.015 5.180 86.015 ;
        RECT 0.000 80.015 5.180 85.015 ;
        RECT 0.000 79.015 0.450 80.015 ;
        RECT 1.340 79.015 5.180 80.015 ;
        RECT 0.000 74.015 5.180 79.015 ;
        RECT 0.000 73.015 0.450 74.015 ;
        RECT 1.340 73.015 5.180 74.015 ;
        RECT 0.000 68.015 5.180 73.015 ;
        RECT 7.060 100.515 67.940 102.855 ;
        RECT 7.060 70.355 9.400 100.515 ;
        RECT 10.320 98.535 64.680 99.645 ;
        RECT 10.320 93.395 11.430 98.535 ;
        RECT 12.500 94.465 62.500 97.465 ;
        RECT 63.570 93.395 64.680 98.535 ;
        RECT 10.320 91.515 64.680 93.395 ;
        RECT 10.320 86.375 11.430 91.515 ;
        RECT 12.500 87.445 62.500 90.445 ;
        RECT 63.570 86.375 64.680 91.515 ;
        RECT 10.320 84.495 64.680 86.375 ;
        RECT 10.320 79.355 11.430 84.495 ;
        RECT 12.500 80.425 62.500 83.425 ;
        RECT 63.570 79.355 64.680 84.495 ;
        RECT 10.320 77.475 64.680 79.355 ;
        RECT 10.320 72.335 11.430 77.475 ;
        RECT 12.500 73.405 62.500 76.405 ;
        RECT 63.570 72.335 64.680 77.475 ;
        RECT 10.320 71.225 64.680 72.335 ;
        RECT 65.600 70.355 67.940 100.515 ;
        RECT 7.060 68.015 67.940 70.355 ;
        RECT 69.820 98.015 75.000 103.015 ;
        RECT 69.820 97.015 73.660 98.015 ;
        RECT 74.550 97.015 75.000 98.015 ;
        RECT 69.820 92.015 75.000 97.015 ;
        RECT 69.820 91.015 73.660 92.015 ;
        RECT 74.550 91.015 75.000 92.015 ;
        RECT 69.820 86.015 75.000 91.015 ;
        RECT 69.820 85.015 73.660 86.015 ;
        RECT 74.550 85.015 75.000 86.015 ;
        RECT 69.820 80.015 75.000 85.015 ;
        RECT 69.820 79.015 73.660 80.015 ;
        RECT 74.550 79.015 75.000 80.015 ;
        RECT 69.820 74.015 75.000 79.015 ;
        RECT 69.820 73.015 73.660 74.015 ;
        RECT 74.550 73.015 75.000 74.015 ;
        RECT 69.820 68.015 75.000 73.015 ;
        RECT 0.000 66.380 0.450 68.015 ;
        RECT 74.550 66.380 75.000 68.015 ;
        RECT 0.000 65.540 75.000 66.380 ;
      LAYER Metal2 ;
        RECT 0.000 318.000 0.450 325.000 ;
        RECT 0.000 246.000 0.450 253.000 ;
        RECT 1.140 68.015 3.680 348.390 ;
        RECT 4.670 340.790 6.290 345.195 ;
        RECT 4.130 334.210 6.370 340.790 ;
        RECT 4.670 329.315 6.290 334.210 ;
        RECT 3.980 254.000 4.980 317.000 ;
        RECT 5.520 246.495 6.520 329.315 ;
        RECT 4.670 230.615 6.520 246.495 ;
        RECT 5.520 228.820 6.520 230.615 ;
        RECT 4.130 214.180 6.520 228.820 ;
        RECT 4.670 212.790 6.520 214.180 ;
        RECT 4.130 206.210 6.520 212.790 ;
        RECT 4.670 196.820 6.520 206.210 ;
        RECT 4.130 182.180 6.520 196.820 ;
        RECT 4.670 180.820 6.520 182.180 ;
        RECT 4.130 166.180 6.520 180.820 ;
        RECT 5.520 164.820 6.520 166.180 ;
        RECT 4.130 150.180 6.520 164.820 ;
        RECT 5.520 148.820 6.520 150.180 ;
        RECT 4.130 134.180 6.520 148.820 ;
        RECT 5.520 124.790 6.520 134.180 ;
        RECT 4.130 118.210 6.520 124.790 ;
        RECT 5.520 68.015 6.520 118.210 ;
        RECT 6.820 68.015 9.360 348.390 ;
        RECT 9.660 68.015 12.200 348.390 ;
        RECT 12.500 68.015 15.040 348.390 ;
        RECT 15.340 65.325 17.880 350.000 ;
        RECT 18.180 68.015 20.720 348.390 ;
        RECT 21.020 65.325 23.560 349.000 ;
        RECT 23.860 68.015 26.400 348.390 ;
        RECT 26.700 65.325 29.240 349.000 ;
        RECT 29.540 68.015 32.080 348.390 ;
        RECT 32.380 65.325 34.920 349.000 ;
        RECT 35.220 68.015 37.350 348.390 ;
        RECT 37.650 68.015 39.780 348.390 ;
        RECT 40.080 65.325 42.620 349.000 ;
        RECT 42.920 68.015 45.460 348.390 ;
        RECT 45.760 65.325 48.300 349.000 ;
        RECT 48.600 68.015 51.140 348.390 ;
        RECT 51.440 65.325 53.980 349.000 ;
        RECT 54.280 68.015 56.820 348.390 ;
        RECT 57.120 65.325 59.660 349.000 ;
        RECT 59.960 68.015 62.500 348.390 ;
        RECT 62.800 68.015 65.340 348.390 ;
        RECT 65.640 325.650 68.180 348.390 ;
        RECT 65.640 246.000 66.640 325.000 ;
        RECT 67.180 244.820 68.180 325.650 ;
        RECT 65.790 244.815 68.180 244.820 ;
        RECT 65.640 68.015 68.180 244.815 ;
        RECT 68.480 68.015 71.020 348.390 ;
        RECT 71.320 68.015 73.860 348.390 ;
        RECT 74.550 318.000 75.000 325.000 ;
        RECT 74.550 246.000 75.000 253.000 ;
        RECT 3.500 62.000 71.500 65.325 ;
        RECT 3.500 2.000 7.500 62.000 ;
        RECT 8.840 2.000 10.540 62.000 ;
        RECT 10.840 2.000 12.540 62.000 ;
        RECT 12.840 2.000 14.540 62.000 ;
        RECT 14.840 2.000 16.540 62.000 ;
        RECT 16.840 2.000 18.540 62.000 ;
        RECT 18.840 2.000 20.540 62.000 ;
        RECT 20.840 2.000 22.540 62.000 ;
        RECT 22.840 2.000 24.540 62.000 ;
        RECT 24.840 2.000 26.540 62.000 ;
        RECT 26.840 2.000 28.540 62.000 ;
        RECT 28.840 2.000 30.540 62.000 ;
        RECT 30.840 2.000 32.540 62.000 ;
        RECT 32.840 2.000 34.540 62.000 ;
        RECT 34.840 2.000 36.540 62.000 ;
        RECT 36.840 2.000 38.540 62.000 ;
        RECT 38.840 2.000 40.540 62.000 ;
        RECT 40.840 2.000 42.540 62.000 ;
        RECT 42.840 2.000 44.540 62.000 ;
        RECT 44.840 2.000 46.540 62.000 ;
        RECT 46.840 2.000 48.540 62.000 ;
        RECT 48.840 2.000 50.540 62.000 ;
        RECT 50.840 2.000 52.540 62.000 ;
        RECT 52.840 2.000 54.540 62.000 ;
        RECT 54.840 2.000 56.540 62.000 ;
        RECT 56.840 2.000 58.540 62.000 ;
        RECT 58.840 2.000 60.540 62.000 ;
        RECT 60.840 2.000 62.540 62.000 ;
        RECT 62.840 2.000 64.540 62.000 ;
        RECT 64.840 2.000 66.540 62.000 ;
        RECT 67.500 2.000 71.500 62.000 ;
        RECT 3.500 0.000 71.500 2.000 ;
      LAYER Metal3 ;
        RECT 1.000 342.000 74.000 348.390 ;
        RECT 1.000 334.000 74.000 341.000 ;
        RECT 1.000 326.000 74.000 333.000 ;
        RECT 1.000 318.000 74.000 325.000 ;
        RECT 1.000 310.000 74.000 317.000 ;
        RECT 1.000 302.000 74.000 309.000 ;
        RECT 1.000 294.000 74.000 301.000 ;
        RECT 1.000 286.000 74.000 293.000 ;
        RECT 1.000 278.000 74.000 285.000 ;
        RECT 4.685 277.000 19.685 278.000 ;
        RECT 21.685 277.000 36.685 278.000 ;
        RECT 38.685 277.000 53.685 278.000 ;
        RECT 55.685 277.000 70.685 278.000 ;
        RECT 1.000 270.000 74.000 277.000 ;
        RECT 4.685 269.000 19.685 270.000 ;
        RECT 21.685 269.000 36.685 270.000 ;
        RECT 38.685 269.000 53.685 270.000 ;
        RECT 55.685 269.000 70.685 270.000 ;
        RECT 1.000 262.000 74.000 269.000 ;
        RECT 1.000 254.000 74.000 261.000 ;
        RECT 1.000 246.000 74.000 253.000 ;
        RECT 1.000 230.000 74.000 245.000 ;
        RECT 1.000 214.000 74.000 229.000 ;
        RECT 4.685 213.000 19.685 214.000 ;
        RECT 21.685 213.000 36.685 214.000 ;
        RECT 38.685 213.000 53.685 214.000 ;
        RECT 55.685 213.000 70.685 214.000 ;
        RECT 1.000 206.000 74.000 213.000 ;
        RECT 1.000 198.000 74.000 205.000 ;
        RECT 1.000 182.000 74.000 197.000 ;
        RECT 4.685 181.000 19.685 182.000 ;
        RECT 21.685 181.000 36.685 182.000 ;
        RECT 38.685 181.000 53.685 182.000 ;
        RECT 55.685 181.000 70.685 182.000 ;
        RECT 1.000 166.000 74.000 181.000 ;
        RECT 4.685 165.000 19.685 166.000 ;
        RECT 21.685 165.000 36.685 166.000 ;
        RECT 38.685 165.000 53.685 166.000 ;
        RECT 55.685 165.000 70.685 166.000 ;
        RECT 1.000 150.000 74.000 165.000 ;
        RECT 4.685 149.000 19.685 150.000 ;
        RECT 21.685 149.000 36.685 150.000 ;
        RECT 38.685 149.000 53.685 150.000 ;
        RECT 55.685 149.000 70.685 150.000 ;
        RECT 1.000 134.000 74.000 149.000 ;
        RECT 1.000 126.000 74.000 133.000 ;
        RECT 1.000 118.000 74.000 125.000 ;
        RECT 1.000 102.000 74.000 117.000 ;
        RECT 4.685 101.000 19.685 102.000 ;
        RECT 21.685 101.000 36.685 102.000 ;
        RECT 38.685 101.000 53.685 102.000 ;
        RECT 55.685 101.000 70.685 102.000 ;
        RECT 1.000 86.000 74.000 101.000 ;
        RECT 4.685 85.000 19.685 86.000 ;
        RECT 21.685 85.000 36.685 86.000 ;
        RECT 38.685 85.000 53.685 86.000 ;
        RECT 55.685 85.000 70.685 86.000 ;
        RECT 1.000 70.000 74.000 85.000 ;
        RECT 3.500 61.600 71.500 65.325 ;
        RECT 3.500 2.290 7.500 61.600 ;
        RECT 8.840 2.290 10.540 61.600 ;
        RECT 10.840 2.290 12.540 61.600 ;
        RECT 12.840 2.290 14.540 61.600 ;
        RECT 14.840 2.290 16.540 61.600 ;
        RECT 16.840 2.290 18.540 61.600 ;
        RECT 18.840 2.290 20.540 61.600 ;
        RECT 20.840 2.290 22.540 61.600 ;
        RECT 22.840 2.290 24.540 61.600 ;
        RECT 24.840 2.290 26.540 61.600 ;
        RECT 26.840 2.290 28.540 61.600 ;
        RECT 28.840 2.290 30.540 61.600 ;
        RECT 30.840 2.290 32.540 61.600 ;
        RECT 32.840 2.290 34.540 61.600 ;
        RECT 34.840 2.290 36.540 61.600 ;
        RECT 36.840 2.290 38.540 61.600 ;
        RECT 38.840 2.290 40.540 61.600 ;
        RECT 40.840 2.290 42.540 61.600 ;
        RECT 42.840 2.290 44.540 61.600 ;
        RECT 44.840 2.290 46.540 61.600 ;
        RECT 46.840 2.290 48.540 61.600 ;
        RECT 48.840 2.290 50.540 61.600 ;
        RECT 50.840 2.290 52.540 61.600 ;
        RECT 52.840 2.290 54.540 61.600 ;
        RECT 54.840 2.290 56.540 61.600 ;
        RECT 56.840 2.290 58.540 61.600 ;
        RECT 58.840 2.290 60.540 61.600 ;
        RECT 60.840 2.290 62.540 61.600 ;
        RECT 62.840 2.290 64.540 61.600 ;
        RECT 64.840 2.290 66.540 61.600 ;
        RECT 67.500 2.290 71.500 61.600 ;
        RECT 3.500 0.000 71.500 2.290 ;
      LAYER Metal4 ;
        RECT 1.000 342.000 74.000 348.390 ;
        RECT 1.000 334.000 74.000 341.000 ;
        RECT 1.000 326.000 74.000 333.000 ;
        RECT 1.000 318.000 74.000 325.000 ;
        RECT 1.000 310.000 74.000 317.000 ;
        RECT 1.000 302.000 74.000 309.000 ;
        RECT 1.000 294.000 74.000 301.000 ;
        RECT 1.000 286.000 74.000 293.000 ;
        RECT 1.000 278.000 74.000 285.000 ;
        RECT 4.685 277.000 19.685 278.000 ;
        RECT 21.685 277.000 36.685 278.000 ;
        RECT 38.685 277.000 53.685 278.000 ;
        RECT 55.685 277.000 70.685 278.000 ;
        RECT 1.000 270.000 74.000 277.000 ;
        RECT 4.685 269.000 19.685 270.000 ;
        RECT 21.685 269.000 36.685 270.000 ;
        RECT 38.685 269.000 53.685 270.000 ;
        RECT 55.685 269.000 70.685 270.000 ;
        RECT 1.000 262.000 74.000 269.000 ;
        RECT 1.000 254.000 74.000 261.000 ;
        RECT 1.000 246.000 74.000 253.000 ;
        RECT 1.000 230.000 74.000 245.000 ;
        RECT 1.000 214.000 74.000 229.000 ;
        RECT 4.685 213.000 19.685 214.000 ;
        RECT 21.685 213.000 36.685 214.000 ;
        RECT 38.685 213.000 53.685 214.000 ;
        RECT 55.685 213.000 70.685 214.000 ;
        RECT 1.000 206.000 74.000 213.000 ;
        RECT 1.000 198.000 74.000 205.000 ;
        RECT 1.000 182.000 74.000 197.000 ;
        RECT 4.685 181.000 19.685 182.000 ;
        RECT 21.685 181.000 36.685 182.000 ;
        RECT 38.685 181.000 53.685 182.000 ;
        RECT 55.685 181.000 70.685 182.000 ;
        RECT 1.000 166.000 74.000 181.000 ;
        RECT 4.685 165.000 19.685 166.000 ;
        RECT 21.685 165.000 36.685 166.000 ;
        RECT 38.685 165.000 53.685 166.000 ;
        RECT 55.685 165.000 70.685 166.000 ;
        RECT 1.000 150.000 74.000 165.000 ;
        RECT 4.685 149.000 19.685 150.000 ;
        RECT 21.685 149.000 36.685 150.000 ;
        RECT 38.685 149.000 53.685 150.000 ;
        RECT 55.685 149.000 70.685 150.000 ;
        RECT 1.000 134.000 74.000 149.000 ;
        RECT 1.000 126.000 74.000 133.000 ;
        RECT 1.000 118.000 74.000 125.000 ;
        RECT 1.000 102.000 74.000 117.000 ;
        RECT 4.685 101.000 19.685 102.000 ;
        RECT 21.685 101.000 36.685 102.000 ;
        RECT 38.685 101.000 53.685 102.000 ;
        RECT 55.685 101.000 70.685 102.000 ;
        RECT 1.000 86.000 74.000 101.000 ;
        RECT 4.685 85.000 19.685 86.000 ;
        RECT 21.685 85.000 36.685 86.000 ;
        RECT 38.685 85.000 53.685 86.000 ;
        RECT 55.685 85.000 70.685 86.000 ;
        RECT 1.000 70.000 74.000 85.000 ;
        RECT 3.500 61.600 71.500 65.325 ;
        RECT 3.500 2.290 7.500 61.600 ;
        RECT 8.840 2.290 10.540 61.600 ;
        RECT 10.840 2.290 12.540 61.600 ;
        RECT 12.840 2.290 14.540 61.600 ;
        RECT 14.840 2.290 16.540 61.600 ;
        RECT 16.840 2.290 18.540 61.600 ;
        RECT 18.840 2.290 20.540 61.600 ;
        RECT 20.840 2.290 22.540 61.600 ;
        RECT 22.840 2.290 24.540 61.600 ;
        RECT 24.840 2.290 26.540 61.600 ;
        RECT 26.840 2.290 28.540 61.600 ;
        RECT 28.840 2.290 30.540 61.600 ;
        RECT 30.840 2.290 32.540 61.600 ;
        RECT 32.840 2.290 34.540 61.600 ;
        RECT 34.840 2.290 36.540 61.600 ;
        RECT 36.840 2.290 38.540 61.600 ;
        RECT 38.840 2.290 40.540 61.600 ;
        RECT 40.840 2.290 42.540 61.600 ;
        RECT 42.840 2.290 44.540 61.600 ;
        RECT 44.840 2.290 46.540 61.600 ;
        RECT 46.840 2.290 48.540 61.600 ;
        RECT 48.840 2.290 50.540 61.600 ;
        RECT 50.840 2.290 52.540 61.600 ;
        RECT 52.840 2.290 54.540 61.600 ;
        RECT 54.840 2.290 56.540 61.600 ;
        RECT 56.840 2.290 58.540 61.600 ;
        RECT 58.840 2.290 60.540 61.600 ;
        RECT 60.840 2.290 62.540 61.600 ;
        RECT 62.840 2.290 64.540 61.600 ;
        RECT 64.840 2.290 66.540 61.600 ;
        RECT 67.500 2.290 71.500 61.600 ;
        RECT 3.500 0.000 71.500 2.290 ;
      LAYER Metal5 ;
        RECT 1.000 342.000 74.000 348.390 ;
        RECT 1.000 334.000 74.000 341.000 ;
        RECT 1.000 326.000 74.000 333.000 ;
        RECT 1.000 318.000 74.000 325.000 ;
        RECT 1.000 310.000 74.000 317.000 ;
        RECT 1.000 302.000 74.000 309.000 ;
        RECT 1.000 294.000 74.000 301.000 ;
        RECT 1.000 286.000 74.000 293.000 ;
        RECT 1.000 278.000 74.000 285.000 ;
        RECT 4.685 277.000 19.685 278.000 ;
        RECT 21.685 277.000 36.685 278.000 ;
        RECT 38.685 277.000 53.685 278.000 ;
        RECT 55.685 277.000 70.685 278.000 ;
        RECT 1.000 270.000 74.000 277.000 ;
        RECT 4.685 269.000 19.685 270.000 ;
        RECT 21.685 269.000 36.685 270.000 ;
        RECT 38.685 269.000 53.685 270.000 ;
        RECT 55.685 269.000 70.685 270.000 ;
        RECT 1.000 262.000 74.000 269.000 ;
        RECT 1.000 254.000 74.000 261.000 ;
        RECT 1.000 246.000 74.000 253.000 ;
        RECT 1.000 230.000 74.000 245.000 ;
        RECT 1.000 214.000 74.000 229.000 ;
        RECT 4.685 213.000 19.685 214.000 ;
        RECT 21.685 213.000 36.685 214.000 ;
        RECT 38.685 213.000 53.685 214.000 ;
        RECT 55.685 213.000 70.685 214.000 ;
        RECT 1.000 206.000 74.000 213.000 ;
        RECT 1.000 198.000 74.000 205.000 ;
        RECT 1.000 182.000 74.000 197.000 ;
        RECT 4.685 181.000 19.685 182.000 ;
        RECT 21.685 181.000 36.685 182.000 ;
        RECT 38.685 181.000 53.685 182.000 ;
        RECT 55.685 181.000 70.685 182.000 ;
        RECT 1.000 166.000 74.000 181.000 ;
        RECT 4.685 165.000 19.685 166.000 ;
        RECT 21.685 165.000 36.685 166.000 ;
        RECT 38.685 165.000 53.685 166.000 ;
        RECT 55.685 165.000 70.685 166.000 ;
        RECT 1.000 150.000 74.000 165.000 ;
        RECT 4.685 149.000 19.685 150.000 ;
        RECT 21.685 149.000 36.685 150.000 ;
        RECT 38.685 149.000 53.685 150.000 ;
        RECT 55.685 149.000 70.685 150.000 ;
        RECT 1.000 134.000 74.000 149.000 ;
        RECT 1.000 126.000 74.000 133.000 ;
        RECT 1.000 118.000 74.000 125.000 ;
        RECT 1.000 102.000 74.000 117.000 ;
        RECT 4.685 101.000 19.685 102.000 ;
        RECT 21.685 101.000 36.685 102.000 ;
        RECT 38.685 101.000 53.685 102.000 ;
        RECT 55.685 101.000 70.685 102.000 ;
        RECT 1.000 86.000 74.000 101.000 ;
        RECT 4.685 85.000 19.685 86.000 ;
        RECT 21.685 85.000 36.685 86.000 ;
        RECT 38.685 85.000 53.685 86.000 ;
        RECT 55.685 85.000 70.685 86.000 ;
        RECT 1.000 70.000 74.000 85.000 ;
        RECT 3.500 45.000 71.500 65.325 ;
        RECT 3.500 20.000 25.000 45.000 ;
        RECT 50.000 20.000 71.500 45.000 ;
        RECT 3.500 0.000 71.500 20.000 ;
  END
END gf180mcu_fd_io__asig_5p0_fixed
END LIBRARY

