magic
tech gf180mcuD
magscale 1 10
timestamp 1762867378
<< nwell >>
rect -324 -1656 324 1656
<< mvpmos >>
rect -60 -1400 60 1400
<< mvpdiff >>
rect -148 1387 -60 1400
rect -148 -1387 -135 1387
rect -89 -1387 -60 1387
rect -148 -1400 -60 -1387
rect 60 1387 148 1400
rect 60 -1387 89 1387
rect 135 -1387 148 1387
rect 60 -1400 148 -1387
<< mvpdiffc >>
rect -135 -1387 -89 1387
rect 89 -1387 135 1387
<< mvnsubdiff >>
rect -292 1552 292 1624
rect -292 1508 -220 1552
rect -292 -1508 -279 1508
rect -233 -1508 -220 1508
rect 220 1508 292 1552
rect -292 -1552 -220 -1508
rect 220 -1508 233 1508
rect 279 -1508 292 1508
rect 220 -1552 292 -1508
rect -292 -1624 292 -1552
<< mvnsubdiffcont >>
rect -279 -1508 -233 1508
rect 233 -1508 279 1508
<< polysilicon >>
rect -60 1479 60 1492
rect -60 1433 -47 1479
rect 47 1433 60 1479
rect -60 1400 60 1433
rect -60 -1433 60 -1400
rect -60 -1479 -47 -1433
rect 47 -1479 60 -1433
rect -60 -1492 60 -1479
<< polycontact >>
rect -47 1433 47 1479
rect -47 -1479 47 -1433
<< metal1 >>
rect -279 1565 279 1611
rect -279 1508 -233 1565
rect 233 1508 279 1565
rect -58 1479 58 1489
rect -58 1433 -47 1479
rect 47 1433 58 1479
rect -135 1387 -89 1398
rect -135 -1398 -89 -1387
rect 89 1387 135 1398
rect 89 -1398 135 -1387
rect -58 -1479 -47 -1433
rect 47 -1479 58 -1433
rect -58 -1489 58 -1479
rect -279 -1565 -233 -1508
rect 233 -1565 279 -1508
rect -279 -1611 279 -1565
<< properties >>
string FIXED_BBOX -256 -1588 256 1588
string gencell pfet_06v0
string library gf180mcu
string parameters w 14.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
