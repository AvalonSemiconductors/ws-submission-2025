VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO r2r_dac_buffered
  CLASS BLOCK ;
  FOREIGN r2r_dac_buffered ;
  ORIGIN 0.000 0.000 ;
  SIZE 324.855 BY 60.590 ;
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2400.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 257.680 56.845 258.665 60.590 ;
    END
  END OUT
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 56.845 58.670 60.585 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.700 56.845 53.690 60.585 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.720 56.845 48.710 60.585 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.740 56.845 43.730 60.585 ;
    END
  END D3
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.760 56.845 38.750 60.585 ;
    END
  END D4
  PIN D5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.780 56.845 33.770 60.585 ;
    END
  END D5
  PIN D6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.800 56.845 28.790 60.585 ;
    END
  END D6
  PIN D7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.820 56.845 23.810 60.585 ;
    END
  END D7
  PIN D8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.840 56.845 18.830 60.585 ;
    END
  END D8
  PIN D9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.860 56.845 13.850 60.585 ;
    END
  END D9
  PIN D10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.880 56.845 8.870 60.585 ;
    END
  END D10
  PIN D11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2.900 56.845 3.890 60.585 ;
    END
  END D11
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 323.795 0.005 324.855 60.590 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 0.000 1.060 60.585 ;
    END
  END VSS
  OBS
      LAYER Pwell ;
        RECT 1.675 51.380 56.450 58.360 ;
        RECT 56.455 51.380 64.565 58.360 ;
        RECT 1.675 47.325 64.565 51.380 ;
        RECT 1.675 12.680 11.330 47.325 ;
      LAYER Nwell ;
        RECT 11.330 23.375 323.225 46.665 ;
        RECT 11.330 12.680 17.560 23.375 ;
      LAYER Pwell ;
        RECT 17.560 12.680 323.225 23.375 ;
        RECT 1.675 0.000 323.225 12.680 ;
      LAYER Metal1 ;
        RECT 0.000 58.360 1.060 60.585 ;
        RECT 0.000 57.905 64.545 58.360 ;
        RECT 0.000 48.395 2.130 57.905 ;
        RECT 2.900 56.845 3.890 57.125 ;
        RECT 2.905 51.985 3.885 52.215 ;
        RECT 2.960 50.155 3.405 51.985 ;
        RECT 4.660 51.155 7.110 57.905 ;
        RECT 7.880 56.845 8.870 57.125 ;
        RECT 7.885 51.985 8.865 52.215 ;
        RECT 4.565 50.925 7.110 51.155 ;
        RECT 2.960 49.170 3.855 50.155 ;
        RECT 7.940 50.150 8.340 51.985 ;
        RECT 9.640 51.155 12.090 57.905 ;
        RECT 12.860 56.845 13.850 57.125 ;
        RECT 12.865 51.985 13.845 52.215 ;
        RECT 9.545 50.925 12.090 51.155 ;
        RECT 12.875 50.150 13.190 51.985 ;
        RECT 14.620 51.155 17.070 57.905 ;
        RECT 17.840 56.845 18.830 57.125 ;
        RECT 17.845 51.985 18.825 52.215 ;
        RECT 14.525 50.925 17.070 51.155 ;
        RECT 17.855 50.150 18.170 51.985 ;
        RECT 19.600 51.155 22.050 57.905 ;
        RECT 22.820 56.845 23.810 57.125 ;
        RECT 22.825 51.985 23.805 52.215 ;
        RECT 19.505 50.925 22.050 51.155 ;
        RECT 22.830 50.150 23.145 51.985 ;
        RECT 24.580 51.155 27.030 57.905 ;
        RECT 27.800 56.845 28.790 57.125 ;
        RECT 27.805 51.985 28.785 52.215 ;
        RECT 24.485 50.925 27.030 51.155 ;
        RECT 27.810 50.150 28.125 51.985 ;
        RECT 29.560 51.155 32.010 57.905 ;
        RECT 32.780 56.845 33.770 57.125 ;
        RECT 32.785 51.985 33.765 52.215 ;
        RECT 29.465 50.925 32.010 51.155 ;
        RECT 32.790 50.150 33.105 51.985 ;
        RECT 34.540 51.155 36.990 57.905 ;
        RECT 37.760 56.845 38.750 57.125 ;
        RECT 34.445 50.925 36.990 51.155 ;
        RECT 37.765 51.985 38.745 52.215 ;
        RECT 37.765 50.150 38.080 51.985 ;
        RECT 39.520 51.155 41.970 57.905 ;
        RECT 42.740 56.845 43.730 57.125 ;
        RECT 39.425 50.925 41.970 51.155 ;
        RECT 42.745 51.985 43.725 52.215 ;
        RECT 42.745 50.150 43.060 51.985 ;
        RECT 44.500 51.155 46.950 57.905 ;
        RECT 47.720 56.845 48.710 57.125 ;
        RECT 47.725 51.985 48.705 52.215 ;
        RECT 44.405 50.925 46.950 51.155 ;
        RECT 48.010 50.150 48.325 51.985 ;
        RECT 49.480 51.155 51.930 57.905 ;
        RECT 52.700 56.845 53.690 57.125 ;
        RECT 52.705 51.985 53.685 52.215 ;
        RECT 49.385 50.925 51.930 51.155 ;
        RECT 52.990 50.150 53.305 51.985 ;
        RECT 54.460 51.155 56.910 57.905 ;
        RECT 57.680 56.845 58.670 57.125 ;
        RECT 57.680 52.215 58.365 52.245 ;
        RECT 57.680 51.985 58.665 52.215 ;
        RECT 59.440 51.155 64.545 57.905 ;
        RECT 54.365 50.925 64.545 51.155 ;
        RECT 57.740 50.150 58.000 50.160 ;
        RECT 63.660 50.150 64.545 50.925 ;
        RECT 5.820 49.170 8.340 50.150 ;
        RECT 10.800 49.170 13.190 50.150 ;
        RECT 15.780 49.170 18.170 50.150 ;
        RECT 20.760 49.170 23.145 50.150 ;
        RECT 25.740 49.170 28.125 50.150 ;
        RECT 30.720 49.170 33.105 50.150 ;
        RECT 35.700 49.170 38.080 50.150 ;
        RECT 40.680 49.170 43.060 50.150 ;
        RECT 45.660 49.170 48.325 50.150 ;
        RECT 50.640 49.170 53.305 50.150 ;
        RECT 55.620 49.170 58.000 50.150 ;
        RECT 62.600 49.170 64.545 50.150 ;
        RECT 57.740 49.165 58.000 49.170 ;
        RECT 63.660 48.395 64.545 49.170 ;
        RECT 0.000 47.355 64.545 48.395 ;
        RECT 0.000 45.365 5.400 47.355 ;
        RECT 6.060 46.665 11.400 46.670 ;
        RECT 323.795 46.665 324.855 60.590 ;
        RECT 6.060 45.670 324.855 46.665 ;
        RECT 0.000 45.135 11.090 45.365 ;
        RECT 0.000 42.765 5.570 45.135 ;
        RECT 6.340 44.075 7.330 44.335 ;
        RECT 0.000 20.015 2.130 42.765 ;
        RECT 2.900 41.705 3.890 41.965 ;
        RECT 4.660 32.385 5.570 42.765 ;
        RECT 6.340 33.150 7.330 33.445 ;
        RECT 8.100 32.385 8.330 45.135 ;
        RECT 9.055 44.015 10.135 44.400 ;
        RECT 9.105 32.385 10.085 33.445 ;
        RECT 10.860 32.385 11.090 45.135 ;
        RECT 4.660 32.155 11.090 32.385 ;
        RECT 11.330 44.665 324.855 45.670 ;
        RECT 4.660 26.835 5.340 32.155 ;
        RECT 6.335 31.290 7.335 31.750 ;
        RECT 6.335 30.325 10.065 31.290 ;
        RECT 4.660 26.605 8.305 26.835 ;
        RECT 2.905 25.910 3.885 25.920 ;
        RECT 2.860 25.485 3.935 25.910 ;
        RECT 2.905 20.845 3.885 25.485 ;
        RECT 4.660 20.015 5.545 26.605 ;
        RECT 6.310 25.535 7.310 25.810 ;
        RECT 0.000 0.455 5.545 20.015 ;
        RECT 8.075 13.435 8.305 26.605 ;
        RECT 9.065 21.005 10.065 30.325 ;
        RECT 10.470 13.435 10.920 32.155 ;
        RECT 11.330 29.015 12.455 44.665 ;
        RECT 13.330 44.005 13.910 44.285 ;
        RECT 14.785 43.830 15.015 44.665 ;
        RECT 15.890 44.005 16.470 44.285 ;
        RECT 17.345 44.170 324.855 44.665 ;
        RECT 17.345 43.830 18.415 44.170 ;
        RECT 19.250 43.940 321.550 44.170 ;
        RECT 12.945 41.150 13.175 43.830 ;
        RECT 12.855 30.515 13.175 41.150 ;
        RECT 12.945 29.850 13.175 30.515 ;
        RECT 14.065 29.850 15.015 43.830 ;
        RECT 15.415 29.850 15.735 43.830 ;
        RECT 16.625 35.610 18.415 43.830 ;
        RECT 18.645 43.205 19.075 43.785 ;
        RECT 119.350 43.280 120.290 43.710 ;
        RECT 220.510 43.280 221.450 43.710 ;
        RECT 321.725 43.205 322.155 43.785 ;
        RECT 18.645 42.665 18.920 43.205 ;
        RECT 120.665 43.050 167.535 43.140 ;
        RECT 221.920 43.050 321.150 43.140 ;
        RECT 19.250 42.820 321.550 43.050 ;
        RECT 321.820 42.665 322.155 43.205 ;
        RECT 18.645 42.085 19.075 42.665 ;
        RECT 119.350 42.160 120.290 42.590 ;
        RECT 220.510 42.160 221.450 42.590 ;
        RECT 321.725 42.085 322.155 42.665 ;
        RECT 18.645 41.545 18.920 42.085 ;
        RECT 19.360 41.930 118.980 42.020 ;
        RECT 173.070 41.930 219.900 42.080 ;
        RECT 19.250 41.700 321.550 41.930 ;
        RECT 321.820 41.545 322.155 42.085 ;
        RECT 18.645 40.965 19.075 41.545 ;
        RECT 119.350 41.040 120.290 41.470 ;
        RECT 220.510 41.040 221.450 41.470 ;
        RECT 321.725 40.965 322.155 41.545 ;
        RECT 18.645 40.425 18.920 40.965 ;
        RECT 120.680 40.810 167.550 40.900 ;
        RECT 221.925 40.810 321.155 40.900 ;
        RECT 19.250 40.580 321.550 40.810 ;
        RECT 321.820 40.425 322.155 40.965 ;
        RECT 18.645 39.845 19.075 40.425 ;
        RECT 119.350 39.920 120.290 40.350 ;
        RECT 220.510 39.920 221.450 40.350 ;
        RECT 321.725 39.845 322.155 40.425 ;
        RECT 18.645 39.305 18.920 39.845 ;
        RECT 19.380 39.690 119.000 39.780 ;
        RECT 173.055 39.690 219.885 39.840 ;
        RECT 19.250 39.460 321.550 39.690 ;
        RECT 321.820 39.305 322.155 39.845 ;
        RECT 18.645 38.725 19.075 39.305 ;
        RECT 119.350 38.800 120.290 39.230 ;
        RECT 220.510 38.800 221.450 39.230 ;
        RECT 321.725 38.725 322.155 39.305 ;
        RECT 18.645 38.185 18.920 38.725 ;
        RECT 120.670 38.570 167.540 38.660 ;
        RECT 221.930 38.570 321.160 38.660 ;
        RECT 19.250 38.340 321.550 38.570 ;
        RECT 321.820 38.185 322.155 38.725 ;
        RECT 18.645 37.605 19.075 38.185 ;
        RECT 119.350 37.680 120.290 38.110 ;
        RECT 220.510 37.680 221.450 38.110 ;
        RECT 321.725 37.605 322.155 38.185 ;
        RECT 18.645 37.065 18.920 37.605 ;
        RECT 19.380 37.450 119.000 37.540 ;
        RECT 173.035 37.450 219.865 37.600 ;
        RECT 19.250 37.220 321.550 37.450 ;
        RECT 321.820 37.065 322.155 37.605 ;
        RECT 18.645 36.485 19.075 37.065 ;
        RECT 119.350 36.560 120.290 36.990 ;
        RECT 220.510 36.560 221.450 36.990 ;
        RECT 321.725 36.485 322.155 37.065 ;
        RECT 120.680 36.330 167.550 36.420 ;
        RECT 221.905 36.330 321.135 36.420 ;
        RECT 19.250 36.100 321.550 36.330 ;
        RECT 322.385 35.610 324.855 44.170 ;
        RECT 16.625 32.890 324.855 35.610 ;
        RECT 16.625 29.850 18.415 32.890 ;
        RECT 19.250 32.660 321.550 32.890 ;
        RECT 13.330 29.395 13.910 29.675 ;
        RECT 14.785 29.015 15.015 29.850 ;
        RECT 15.890 29.395 16.470 29.675 ;
        RECT 17.345 29.015 18.415 29.850 ;
        RECT 11.330 28.785 18.415 29.015 ;
        RECT 8.075 13.205 11.065 13.435 ;
        RECT 6.305 1.255 7.305 1.515 ;
        RECT 8.075 0.455 8.305 13.205 ;
        RECT 10.470 12.415 11.065 13.205 ;
        RECT 11.330 13.135 11.785 28.785 ;
        RECT 12.660 28.125 13.240 28.405 ;
        RECT 12.275 21.055 12.505 27.950 ;
        RECT 12.025 13.970 12.505 21.055 ;
        RECT 12.750 13.795 13.105 28.125 ;
        RECT 13.395 26.925 13.625 27.950 ;
        RECT 13.395 15.305 13.715 26.925 ;
        RECT 13.395 13.970 13.625 15.305 ;
        RECT 12.660 13.515 13.240 13.795 ;
        RECT 14.115 13.135 14.345 28.785 ;
        RECT 15.220 28.125 15.800 28.405 ;
        RECT 14.835 26.900 15.065 27.950 ;
        RECT 14.740 15.280 15.065 26.900 ;
        RECT 14.835 13.970 15.065 15.280 ;
        RECT 15.390 14.955 15.625 28.125 ;
        RECT 15.305 13.795 15.625 14.955 ;
        RECT 15.955 26.930 16.185 27.950 ;
        RECT 15.955 15.570 16.275 26.930 ;
        RECT 16.675 24.330 18.415 28.785 ;
        RECT 18.645 31.925 19.075 32.505 ;
        RECT 119.350 32.000 120.290 32.430 ;
        RECT 220.510 32.000 221.450 32.430 ;
        RECT 321.725 31.925 322.155 32.505 ;
        RECT 18.645 31.385 18.920 31.925 ;
        RECT 120.660 31.770 167.530 31.860 ;
        RECT 221.945 31.770 321.175 31.860 ;
        RECT 19.250 31.540 321.550 31.770 ;
        RECT 321.820 31.385 322.155 31.925 ;
        RECT 18.645 30.805 19.075 31.385 ;
        RECT 119.350 30.880 120.290 31.310 ;
        RECT 220.510 30.880 221.450 31.310 ;
        RECT 321.725 30.805 322.155 31.385 ;
        RECT 18.645 30.265 18.920 30.805 ;
        RECT 19.360 30.650 118.980 30.740 ;
        RECT 173.065 30.650 219.895 30.800 ;
        RECT 19.250 30.420 321.550 30.650 ;
        RECT 321.820 30.265 322.155 30.805 ;
        RECT 18.645 29.685 19.075 30.265 ;
        RECT 119.350 29.760 120.290 30.190 ;
        RECT 220.510 29.760 221.450 30.190 ;
        RECT 321.725 29.685 322.155 30.265 ;
        RECT 18.645 29.145 18.920 29.685 ;
        RECT 120.665 29.530 167.535 29.620 ;
        RECT 221.970 29.530 321.200 29.620 ;
        RECT 19.250 29.300 321.550 29.530 ;
        RECT 321.820 29.145 322.155 29.685 ;
        RECT 18.645 28.565 19.075 29.145 ;
        RECT 119.350 28.640 120.290 29.070 ;
        RECT 220.510 28.640 221.450 29.070 ;
        RECT 321.725 28.565 322.155 29.145 ;
        RECT 18.645 28.025 18.920 28.565 ;
        RECT 19.390 28.410 119.010 28.500 ;
        RECT 173.070 28.410 219.900 28.560 ;
        RECT 19.250 28.180 321.550 28.410 ;
        RECT 321.820 28.025 322.155 28.565 ;
        RECT 18.645 27.445 19.075 28.025 ;
        RECT 119.350 27.520 120.290 27.950 ;
        RECT 220.510 27.520 221.450 27.950 ;
        RECT 321.725 27.445 322.155 28.025 ;
        RECT 18.645 26.905 18.920 27.445 ;
        RECT 120.655 27.290 167.525 27.380 ;
        RECT 221.980 27.290 321.210 27.380 ;
        RECT 19.250 27.060 321.550 27.290 ;
        RECT 321.820 26.905 322.155 27.445 ;
        RECT 18.645 26.325 19.075 26.905 ;
        RECT 119.350 26.400 120.290 26.830 ;
        RECT 220.510 26.400 221.450 26.830 ;
        RECT 321.725 26.325 322.155 26.905 ;
        RECT 18.645 25.785 18.920 26.325 ;
        RECT 19.355 26.170 118.975 26.260 ;
        RECT 173.060 26.170 219.890 26.320 ;
        RECT 19.250 25.940 321.550 26.170 ;
        RECT 321.820 25.785 322.155 26.325 ;
        RECT 18.645 25.205 19.075 25.785 ;
        RECT 119.350 25.280 120.290 25.710 ;
        RECT 220.510 25.280 221.450 25.710 ;
        RECT 321.725 25.205 322.155 25.785 ;
        RECT 120.665 25.050 167.535 25.140 ;
        RECT 221.935 25.050 321.165 25.140 ;
        RECT 19.250 24.820 321.550 25.050 ;
        RECT 322.385 24.330 324.855 32.890 ;
        RECT 16.675 23.375 324.855 24.330 ;
        RECT 15.955 13.970 16.185 15.570 ;
        RECT 15.220 13.515 15.800 13.795 ;
        RECT 16.675 13.135 16.905 23.375 ;
        RECT 11.330 12.905 16.905 13.135 ;
        RECT 17.560 23.140 22.565 23.145 ;
        RECT 17.560 21.840 323.225 23.140 ;
        RECT 17.560 13.280 18.400 21.840 ;
        RECT 19.235 21.610 321.535 21.840 ;
        RECT 18.630 20.875 19.060 21.455 ;
        RECT 119.335 20.950 120.275 21.380 ;
        RECT 220.495 20.950 221.435 21.380 ;
        RECT 321.710 20.875 322.140 21.455 ;
        RECT 18.630 20.335 18.890 20.875 ;
        RECT 120.695 20.720 167.565 20.810 ;
        RECT 221.925 20.720 321.155 20.810 ;
        RECT 19.235 20.490 321.535 20.720 ;
        RECT 321.880 20.335 322.140 20.875 ;
        RECT 18.630 19.755 19.060 20.335 ;
        RECT 119.335 19.830 120.275 20.260 ;
        RECT 220.495 19.830 221.435 20.260 ;
        RECT 321.710 19.755 322.140 20.335 ;
        RECT 18.630 19.215 18.890 19.755 ;
        RECT 19.375 19.600 118.995 19.690 ;
        RECT 173.160 19.600 219.990 19.755 ;
        RECT 19.235 19.370 321.535 19.600 ;
        RECT 321.880 19.215 322.140 19.755 ;
        RECT 18.630 18.635 19.060 19.215 ;
        RECT 119.335 18.710 120.275 19.140 ;
        RECT 220.495 18.710 221.435 19.140 ;
        RECT 321.710 18.635 322.140 19.215 ;
        RECT 18.630 18.095 18.890 18.635 ;
        RECT 120.690 18.480 167.560 18.570 ;
        RECT 221.945 18.480 321.175 18.570 ;
        RECT 19.235 18.250 321.535 18.480 ;
        RECT 321.880 18.095 322.140 18.635 ;
        RECT 18.630 17.515 19.060 18.095 ;
        RECT 119.335 17.590 120.275 18.020 ;
        RECT 220.495 17.590 221.435 18.020 ;
        RECT 321.710 17.515 322.140 18.095 ;
        RECT 18.630 16.975 18.890 17.515 ;
        RECT 19.385 17.360 119.005 17.450 ;
        RECT 173.160 17.360 219.990 17.515 ;
        RECT 19.235 17.130 321.535 17.360 ;
        RECT 321.880 16.975 322.140 17.515 ;
        RECT 18.630 16.395 19.060 16.975 ;
        RECT 119.335 16.470 120.275 16.900 ;
        RECT 220.495 16.470 221.435 16.900 ;
        RECT 321.710 16.395 322.140 16.975 ;
        RECT 18.630 15.855 18.890 16.395 ;
        RECT 120.675 16.240 167.545 16.330 ;
        RECT 221.955 16.240 321.185 16.330 ;
        RECT 19.235 16.010 321.535 16.240 ;
        RECT 321.880 15.855 322.140 16.395 ;
        RECT 18.630 15.275 19.060 15.855 ;
        RECT 119.335 15.350 120.275 15.780 ;
        RECT 220.495 15.350 221.435 15.780 ;
        RECT 321.710 15.275 322.140 15.855 ;
        RECT 18.630 14.735 18.890 15.275 ;
        RECT 19.365 15.120 118.985 15.210 ;
        RECT 173.155 15.120 219.985 15.275 ;
        RECT 19.235 14.890 321.535 15.120 ;
        RECT 321.880 14.735 322.140 15.275 ;
        RECT 18.630 14.155 19.060 14.735 ;
        RECT 119.335 14.230 120.275 14.660 ;
        RECT 220.495 14.230 221.435 14.660 ;
        RECT 321.710 14.155 322.140 14.735 ;
        RECT 120.680 14.000 167.550 14.095 ;
        RECT 221.930 14.000 321.160 14.090 ;
        RECT 19.235 13.770 321.535 14.000 ;
        RECT 322.370 13.280 323.225 21.840 ;
        RECT 17.560 12.415 323.225 13.280 ;
        RECT 9.075 12.145 10.065 12.405 ;
        RECT 10.470 12.185 323.225 12.415 ;
        RECT 10.470 11.660 12.560 12.185 ;
        RECT 9.080 0.455 10.060 1.515 ;
        RECT 10.835 0.535 12.560 11.660 ;
        RECT 13.435 11.525 14.015 11.830 ;
        RECT 13.435 11.350 13.845 11.525 ;
        RECT 14.890 11.350 15.120 12.185 ;
        RECT 15.995 11.525 16.575 11.830 ;
        RECT 13.050 1.370 13.845 11.350 ;
        RECT 14.170 1.370 15.840 11.350 ;
        RECT 16.175 6.960 16.410 11.525 ;
        RECT 16.095 4.350 16.410 6.960 ;
        RECT 13.435 1.195 13.845 1.370 ;
        RECT 13.435 0.890 14.015 1.195 ;
        RECT 14.890 0.535 15.120 1.370 ;
        RECT 16.175 1.195 16.410 4.350 ;
        RECT 16.730 10.600 16.960 11.350 ;
        RECT 16.730 2.245 17.050 10.600 ;
        RECT 17.450 10.560 323.225 12.185 ;
        RECT 16.730 1.370 16.960 2.245 ;
        RECT 17.450 2.000 18.400 10.560 ;
        RECT 19.235 10.330 321.535 10.560 ;
        RECT 18.630 9.595 19.060 10.175 ;
        RECT 119.335 9.670 120.275 10.100 ;
        RECT 220.495 9.670 221.435 10.100 ;
        RECT 321.710 9.595 322.140 10.175 ;
        RECT 18.630 9.055 18.890 9.595 ;
        RECT 120.690 9.440 167.560 9.530 ;
        RECT 221.920 9.440 321.150 9.530 ;
        RECT 19.235 9.210 321.535 9.440 ;
        RECT 321.880 9.055 322.140 9.595 ;
        RECT 18.630 8.475 19.060 9.055 ;
        RECT 119.335 8.550 120.275 8.980 ;
        RECT 220.495 8.550 221.435 8.980 ;
        RECT 321.710 8.475 322.140 9.055 ;
        RECT 18.630 7.935 18.890 8.475 ;
        RECT 19.355 8.320 118.975 8.410 ;
        RECT 173.165 8.320 219.995 8.475 ;
        RECT 19.235 8.090 321.535 8.320 ;
        RECT 321.880 7.935 322.140 8.475 ;
        RECT 18.630 7.355 19.060 7.935 ;
        RECT 119.335 7.430 120.275 7.860 ;
        RECT 220.495 7.430 221.435 7.860 ;
        RECT 321.710 7.355 322.140 7.935 ;
        RECT 18.630 6.815 18.890 7.355 ;
        RECT 120.695 7.200 167.565 7.290 ;
        RECT 221.925 7.200 321.155 7.290 ;
        RECT 19.235 6.970 321.535 7.200 ;
        RECT 321.880 6.815 322.140 7.355 ;
        RECT 18.630 6.235 19.060 6.815 ;
        RECT 119.335 6.310 120.275 6.740 ;
        RECT 220.495 6.310 221.435 6.740 ;
        RECT 321.710 6.235 322.140 6.815 ;
        RECT 18.630 5.695 18.890 6.235 ;
        RECT 19.355 6.080 118.975 6.170 ;
        RECT 173.215 6.080 220.045 6.235 ;
        RECT 19.235 5.850 321.535 6.080 ;
        RECT 321.880 5.695 322.140 6.235 ;
        RECT 18.630 5.115 19.060 5.695 ;
        RECT 119.335 5.190 120.275 5.620 ;
        RECT 220.495 5.190 221.435 5.620 ;
        RECT 321.710 5.115 322.140 5.695 ;
        RECT 18.630 4.575 18.890 5.115 ;
        RECT 120.675 4.960 167.545 5.050 ;
        RECT 221.950 4.960 321.180 5.050 ;
        RECT 19.235 4.730 321.535 4.960 ;
        RECT 321.880 4.575 322.140 5.115 ;
        RECT 18.630 3.995 19.060 4.575 ;
        RECT 119.335 4.070 120.275 4.500 ;
        RECT 220.495 4.070 221.435 4.500 ;
        RECT 321.710 3.995 322.140 4.575 ;
        RECT 18.630 3.455 18.890 3.995 ;
        RECT 19.295 3.840 118.915 3.930 ;
        RECT 173.130 3.840 219.960 3.995 ;
        RECT 19.235 3.610 321.535 3.840 ;
        RECT 321.880 3.455 322.140 3.995 ;
        RECT 18.630 2.875 19.060 3.455 ;
        RECT 119.335 2.950 120.275 3.380 ;
        RECT 220.495 2.950 221.435 3.380 ;
        RECT 321.710 2.875 322.140 3.455 ;
        RECT 120.660 2.720 167.530 2.810 ;
        RECT 221.905 2.720 321.135 2.810 ;
        RECT 19.235 2.490 321.535 2.720 ;
        RECT 322.370 2.000 323.225 10.560 ;
        RECT 15.995 0.890 16.575 1.195 ;
        RECT 17.450 0.535 323.225 2.000 ;
        RECT 10.835 0.455 323.225 0.535 ;
        RECT 0.000 0.005 323.225 0.455 ;
        RECT 323.795 0.005 324.855 23.375 ;
        RECT 0.000 0.000 11.325 0.005 ;
        RECT 12.330 0.000 323.225 0.005 ;
      LAYER Metal2 ;
        RECT 0.000 0.000 1.060 60.585 ;
        RECT 257.675 56.845 257.680 57.550 ;
        RECT 257.675 53.805 258.660 56.845 ;
        RECT 57.620 51.920 58.365 52.265 ;
        RECT 2.890 41.685 3.895 50.255 ;
        RECT 57.620 49.105 58.050 51.920 ;
        RECT 6.320 44.050 7.340 46.690 ;
        RECT 18.525 44.735 322.225 45.350 ;
        RECT 18.525 44.420 18.930 44.735 ;
        RECT 9.040 43.995 18.930 44.420 ;
        RECT 13.325 43.990 18.930 43.995 ;
        RECT 6.335 30.760 7.335 33.475 ;
        RECT 12.750 30.470 13.215 41.200 ;
        RECT 12.750 28.995 13.100 30.470 ;
        RECT 13.380 29.695 13.925 29.735 ;
        RECT 15.330 29.695 15.745 43.990 ;
        RECT 18.525 29.695 18.930 43.990 ;
        RECT 13.380 29.370 18.930 29.695 ;
        RECT 13.380 29.355 13.925 29.370 ;
        RECT 12.750 28.635 13.725 28.995 ;
        RECT 12.650 25.910 13.080 28.060 ;
        RECT 2.860 25.485 13.080 25.910 ;
        RECT 12.650 25.150 13.080 25.485 ;
        RECT 13.360 26.985 13.725 28.635 ;
        RECT 9.070 21.335 13.075 21.760 ;
        RECT 9.070 12.135 10.065 21.335 ;
        RECT 11.955 11.960 12.370 21.055 ;
        RECT 12.650 17.100 13.075 21.335 ;
        RECT 12.650 14.965 13.080 17.100 ;
        RECT 13.360 15.245 15.120 26.985 ;
        RECT 15.915 19.975 16.290 26.970 ;
        RECT 18.525 25.080 18.930 29.370 ;
        RECT 19.290 25.820 119.030 44.325 ;
        RECT 119.350 25.225 120.290 44.735 ;
        RECT 120.590 24.950 167.590 43.395 ;
        RECT 172.975 25.880 219.980 44.370 ;
        RECT 220.510 25.230 221.450 44.735 ;
        RECT 221.800 24.950 321.335 43.395 ;
        RECT 321.820 25.040 322.225 44.735 ;
        RECT 120.590 22.410 321.335 24.950 ;
        RECT 18.295 19.975 18.910 21.525 ;
        RECT 15.915 17.185 18.910 19.975 ;
        RECT 15.915 15.530 16.290 17.185 ;
        RECT 12.650 14.495 15.685 14.965 ;
        RECT 15.215 13.820 15.685 14.495 ;
        RECT 15.170 13.480 15.840 13.820 ;
        RECT 11.955 11.545 13.385 11.960 ;
        RECT 12.970 6.940 13.385 11.545 ;
        RECT 16.685 10.390 17.060 10.640 ;
        RECT 18.295 10.390 18.910 17.185 ;
        RECT 16.685 7.600 18.910 10.390 ;
        RECT 12.970 6.465 16.405 6.940 ;
        RECT 16.010 4.370 16.405 6.465 ;
        RECT 16.685 2.205 17.060 7.600 ;
        RECT 18.295 2.115 18.910 7.600 ;
        RECT 19.255 3.535 118.965 22.040 ;
        RECT 119.335 2.115 120.275 21.555 ;
        RECT 120.590 2.415 167.590 22.410 ;
        RECT 173.095 3.500 220.100 21.980 ;
        RECT 220.495 2.115 221.435 21.550 ;
        RECT 221.800 2.415 321.335 22.410 ;
        RECT 321.845 2.115 322.250 21.525 ;
        RECT 6.305 1.155 7.310 1.545 ;
        RECT 18.295 1.500 322.250 2.115 ;
        RECT 122.250 1.155 123.200 1.190 ;
        RECT 6.305 0.540 123.200 1.155 ;
        RECT 122.250 0.515 123.200 0.540 ;
        RECT 323.795 0.005 324.855 60.590 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 1.060 60.585 ;
        RECT 257.675 41.925 258.660 55.040 ;
        RECT 257.675 37.175 262.260 41.925 ;
        RECT 122.280 1.190 123.280 4.245 ;
        RECT 122.250 0.540 123.280 1.190 ;
        RECT 122.250 0.515 123.200 0.540 ;
        RECT 323.795 0.005 324.855 60.590 ;
  END
END r2r_dac_buffered
END LIBRARY

