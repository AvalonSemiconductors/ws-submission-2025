magic
tech gf180mcuD
magscale 1 10
timestamp 1762910833
<< nwell >>
rect 298 9023 62677 9333
rect 298 5848 432 9023
rect 1559 7031 1669 9023
rect 42146 7312 42310 7398
rect 62600 7031 62677 9023
rect 1559 6767 62677 7031
rect 1559 5744 1669 6767
rect 1577 5712 1633 5744
rect 1458 4775 1624 5712
rect 62600 4775 62677 6767
rect 1458 4675 62677 4775
rect 1088 2703 1180 2758
rect 1458 2536 1544 4675
<< pwell >>
rect 1544 4557 62677 4675
rect 1544 2565 1621 4557
rect 62597 2565 62677 4557
rect 1544 2536 62677 2565
rect 298 2528 62677 2536
rect 298 16 453 2528
rect 1613 2301 62677 2528
rect 1613 309 1621 2301
rect 62401 392 62482 567
rect 62597 309 62677 2301
rect 1613 16 62677 309
rect 298 0 62677 16
<< polysilicon >>
rect 42146 7312 42310 7398
rect 1088 2703 1180 2758
<< metal1 >>
rect 298 8979 62677 9333
rect 298 5803 477 8979
rect 1547 8978 62677 8979
rect 603 6103 615 8230
rect 891 5970 989 8766
rect 1115 8754 1179 8766
rect 1115 5982 1127 8754
rect 1115 5970 1179 5982
rect 1403 5970 1501 8766
rect 1547 7076 1669 8978
rect 1715 8852 62509 8932
rect 1715 8840 32646 8852
rect 1715 8834 1902 8840
rect 21826 8834 32646 8840
rect 42012 8834 62509 8852
rect 1764 8739 1816 8745
rect 62407 8739 62459 8745
rect 22165 8616 31539 8628
rect 42416 8616 62262 8628
rect 32646 8404 42012 8416
rect 1904 8392 21828 8404
rect 22168 8168 31542 8180
rect 42417 8168 62263 8180
rect 32643 7956 42009 7968
rect 1908 7944 21832 7956
rect 22166 7720 31540 7732
rect 42418 7720 62264 7732
rect 32639 7508 42005 7520
rect 1908 7496 21832 7508
rect 22168 7272 31542 7284
rect 42413 7272 62259 7284
rect 1547 6722 1910 7076
rect 298 2581 343 5803
rect 1547 5757 1669 6722
rect 1715 6578 1910 6676
rect 21834 6722 32640 7076
rect 21834 6584 32640 6676
rect 21835 6578 32640 6584
rect 62555 7076 62677 8978
rect 42006 6722 62677 7076
rect 42006 6578 62509 6676
rect 582 5600 653 5625
rect 582 5042 589 5600
rect 641 5042 653 5600
rect 437 4199 487 4211
rect 437 2800 449 4199
rect 437 2794 487 2800
rect 582 2759 653 5042
rect 763 3061 775 5385
rect 980 3056 992 5380
rect 1110 2991 1157 5625
rect 1275 3114 1287 5386
rect 1413 4821 1669 5757
rect 22164 6360 31538 6372
rect 42421 6360 62267 6372
rect 32645 6148 42011 6160
rect 1904 6136 21828 6148
rect 22165 5912 31539 5924
rect 42426 5912 62272 5924
rect 32646 5700 42012 5712
rect 1910 5688 21834 5700
rect 22163 5464 31537 5476
rect 42428 5464 62274 5476
rect 32644 5252 42010 5264
rect 1903 5240 21827 5252
rect 22165 5016 31539 5028
rect 42419 5016 62265 5028
rect 62555 4821 62677 6722
rect 1413 4675 62677 4821
rect 1544 4628 2545 4629
rect 1544 4512 62677 4628
rect 1093 2759 1105 2991
rect 576 2707 668 2759
rect 1544 2610 1666 4512
rect 1712 4387 62506 4466
rect 1712 4374 32662 4387
rect 1712 4368 1901 4374
rect 21823 4368 32662 4374
rect 21823 4322 21825 4368
rect 42028 4368 62506 4387
rect 22171 4150 31545 4162
rect 42417 4150 62263 4162
rect 32664 3939 42030 3951
rect 1907 3926 21831 3938
rect 21823 3874 21831 3926
rect 22170 3702 31544 3714
rect 42421 3702 62267 3714
rect 32664 3491 42030 3503
rect 1909 3478 21833 3490
rect 21823 3426 21833 3478
rect 22167 3254 31541 3266
rect 42423 3254 62269 3266
rect 32663 3043 42029 3055
rect 1905 3030 21829 3042
rect 21823 2978 21829 3030
rect 22168 2807 31542 2819
rect 42418 2806 62264 2818
rect 297 61 498 2483
rect 719 2270 801 2305
rect 688 2258 801 2270
rect 699 1301 801 2258
rect 688 274 801 1301
rect 912 274 1010 2270
rect 1056 274 1154 2270
rect 1267 1392 1314 2305
rect 1544 2256 1899 2610
rect 1251 1380 1314 1392
rect 1303 882 1314 1380
rect 1251 870 1314 882
rect 719 239 801 274
rect 1267 239 1314 870
rect 1430 449 1442 2120
rect 1544 354 1666 2256
rect 1712 2112 1899 2210
rect 21823 2256 32659 2610
rect 21823 2112 32659 2210
rect 62552 2610 62677 4512
rect 42025 2256 62677 2610
rect 42025 2131 62506 2210
rect 42026 2112 62506 2131
rect 22170 1894 31544 1906
rect 42416 1894 62262 1906
rect 32665 1683 42031 1695
rect 1903 1670 21827 1682
rect 21823 1618 21827 1670
rect 22171 1446 31545 1458
rect 42417 1446 62263 1458
rect 32675 1235 42041 1247
rect 1903 1222 21827 1234
rect 21823 1170 21827 1222
rect 22167 998 31541 1010
rect 42422 998 62268 1010
rect 32658 787 42024 799
rect 1891 774 21815 786
rect 22164 550 31538 562
rect 42413 550 62259 562
rect 62552 354 62677 2256
rect 1544 61 62677 354
rect 297 1 62677 61
rect 498 0 62677 1
<< via1 >>
rect 710 8804 802 8856
rect 1222 8804 1314 8856
rect 615 6103 667 8230
rect 1127 5982 1179 8754
rect 1902 8788 21826 8840
rect 32646 8788 42012 8852
rect 1764 7309 1816 8739
rect 21914 8656 22078 8742
rect 42146 8656 42310 8742
rect 22165 8564 31539 8616
rect 42416 8564 62262 8616
rect 21914 8432 22078 8518
rect 42146 8432 42310 8518
rect 1904 8340 21828 8392
rect 32646 8340 42012 8404
rect 21914 8208 22078 8294
rect 42146 8208 42310 8294
rect 22168 8116 31542 8168
rect 42417 8116 62263 8168
rect 21914 7984 22078 8070
rect 42146 7984 42310 8070
rect 1908 7892 21832 7944
rect 32643 7892 42009 7956
rect 21914 7760 22078 7846
rect 42146 7760 42310 7846
rect 22166 7668 31540 7720
rect 42418 7668 62264 7720
rect 21914 7536 22078 7622
rect 42146 7536 42310 7622
rect 1908 7444 21832 7496
rect 32639 7444 42005 7508
rect 21914 7312 22078 7398
rect 42146 7312 42310 7398
rect 62407 7309 62459 8739
rect 22168 7220 31542 7272
rect 42413 7220 62259 7272
rect 710 5883 802 5935
rect 1222 5883 1314 5935
rect 1910 6584 21834 7115
rect 1910 6532 21835 6584
rect 32640 6532 42006 7116
rect 589 5042 641 5600
rect 449 2800 501 4199
rect 711 3061 763 5385
rect 992 3056 1044 5380
rect 1223 3114 1275 5386
rect 1764 5053 1816 6489
rect 21914 6400 22078 6486
rect 42146 6400 42310 6486
rect 22164 6308 31538 6360
rect 42421 6308 62267 6360
rect 21914 6176 22078 6262
rect 42146 6176 42310 6262
rect 1904 6084 21828 6136
rect 32645 6084 42011 6148
rect 21914 5952 22078 6038
rect 42146 5952 42310 6038
rect 22165 5860 31539 5912
rect 42426 5860 62272 5912
rect 21914 5728 22078 5814
rect 42146 5728 42310 5814
rect 1910 5636 21834 5688
rect 32646 5636 42012 5700
rect 21914 5504 22078 5590
rect 42146 5504 42310 5590
rect 22163 5412 31537 5464
rect 42428 5412 62274 5464
rect 21914 5280 22078 5366
rect 42146 5280 42310 5366
rect 1903 5188 21827 5240
rect 32644 5188 42010 5252
rect 21914 5056 22078 5142
rect 42146 5056 42310 5142
rect 62407 5053 62459 6489
rect 22165 4964 31539 5016
rect 42419 4964 62265 5016
rect 1105 2759 1157 2991
rect 1088 2703 1180 2759
rect 1901 4322 21823 4374
rect 32662 4322 42028 4387
rect 1758 2843 1810 4279
rect 21911 4190 22075 4276
rect 42143 4190 42307 4276
rect 22171 4098 31545 4150
rect 42417 4098 62263 4150
rect 21911 3966 22075 4052
rect 42143 3966 42307 4052
rect 1907 3874 21823 3926
rect 32664 3874 42030 3939
rect 21911 3742 22075 3828
rect 42143 3742 42307 3828
rect 22170 3650 31544 3702
rect 42421 3650 62267 3702
rect 21911 3518 22075 3604
rect 42143 3518 42307 3604
rect 1909 3426 21823 3478
rect 32664 3426 42030 3491
rect 21911 3294 22075 3380
rect 42143 3294 42307 3380
rect 22167 3202 31541 3254
rect 42423 3202 62269 3254
rect 21911 3070 22075 3156
rect 42143 3070 42307 3156
rect 1905 2978 21823 3030
rect 32663 2978 42029 3043
rect 21911 2846 22075 2932
rect 42143 2846 42307 2932
rect 62408 2843 62460 4279
rect 22168 2755 31542 2807
rect 42418 2754 62264 2806
rect 647 1301 699 2258
rect 1251 882 1303 1380
rect 1378 449 1430 2120
rect 1899 2066 21823 2649
rect 32659 2131 42025 2650
rect 32659 2066 42026 2131
rect 1758 587 1810 2023
rect 21911 1934 22075 2020
rect 42143 1934 42307 2020
rect 22170 1842 31544 1894
rect 42416 1842 62262 1894
rect 21911 1710 22075 1796
rect 42143 1710 42307 1796
rect 1903 1618 21823 1670
rect 32665 1618 42031 1683
rect 21911 1486 22075 1572
rect 42143 1486 42307 1572
rect 22171 1394 31545 1446
rect 42417 1394 62263 1446
rect 21911 1262 22075 1348
rect 42143 1262 42307 1348
rect 1903 1170 21823 1222
rect 32675 1170 42041 1235
rect 21911 1038 22075 1124
rect 42143 1038 42307 1124
rect 22167 946 31541 998
rect 42422 946 62268 998
rect 21911 814 22075 900
rect 42143 814 42307 900
rect 1891 722 21815 774
rect 32658 722 42024 787
rect 21911 590 22075 676
rect 42143 590 42307 676
rect 62408 587 62460 2023
rect 22164 498 31538 550
rect 42413 498 62259 550
<< metal2 >>
rect 1737 8947 62477 9070
rect 1737 8884 1818 8947
rect 0 8856 1818 8884
rect 0 8804 710 8856
rect 802 8804 1222 8856
rect 1314 8804 1818 8856
rect 0 8799 1818 8804
rect 697 8798 1818 8799
rect 1098 8754 1181 8798
rect 582 8230 675 8240
rect 582 6103 615 8230
rect 667 6103 675 8230
rect 582 6094 675 6103
rect 582 5799 652 6094
rect 1098 5982 1127 8754
rect 1179 5982 1181 8754
rect 708 5939 817 5947
rect 1098 5939 1181 5982
rect 1737 8739 1818 8798
rect 1737 7309 1764 8739
rect 1816 7309 1818 8739
rect 1737 6489 1818 7309
rect 1737 5939 1764 6489
rect 708 5935 1764 5939
rect 708 5883 710 5935
rect 802 5883 1222 5935
rect 1314 5883 1764 5935
rect 708 5874 1764 5883
rect 708 5871 817 5874
rect 582 5727 777 5799
rect 562 5600 648 5612
rect 562 5182 589 5600
rect 0 5097 589 5182
rect 562 5042 589 5097
rect 641 5042 648 5600
rect 562 5030 648 5042
rect 704 5397 777 5727
rect 704 5385 1056 5397
rect 0 4267 647 4352
rect 423 4199 506 4211
rect 423 2800 449 4199
rect 501 2800 506 4199
rect 562 3420 647 4267
rect 562 2993 648 3420
rect 704 3061 711 5385
rect 763 5380 1056 5385
rect 763 3061 992 5380
rect 704 3056 992 3061
rect 1044 3056 1056 5380
rect 1215 5386 1290 5394
rect 1215 3114 1223 5386
rect 1275 3995 1290 5386
rect 1737 5053 1764 5874
rect 1816 5053 1818 6489
rect 1890 8840 21838 8865
rect 1890 8788 1902 8840
rect 21826 8788 21838 8840
rect 1890 8392 21838 8788
rect 1890 8340 1904 8392
rect 21828 8340 21838 8392
rect 1890 7944 21838 8340
rect 1890 7892 1908 7944
rect 21832 7892 21838 7944
rect 1890 7496 21838 7892
rect 1890 7444 1908 7496
rect 21832 7444 21838 7496
rect 1890 7115 21838 7444
rect 1890 6532 1910 7115
rect 21834 6584 21838 7115
rect 21835 6532 21838 6584
rect 1890 6136 21838 6532
rect 1890 6084 1904 6136
rect 21828 6084 21838 6136
rect 1890 5688 21838 6084
rect 1890 5636 1910 5688
rect 21834 5636 21838 5688
rect 1890 5240 21838 5636
rect 1890 5188 1903 5240
rect 21827 5188 21838 5240
rect 1890 5164 21838 5188
rect 21902 8742 22090 8947
rect 21902 8656 21914 8742
rect 22078 8656 22090 8742
rect 32627 8852 42028 8874
rect 32627 8788 32646 8852
rect 42012 8788 42028 8852
rect 21902 8518 22090 8656
rect 21902 8432 21914 8518
rect 22078 8432 22090 8518
rect 21902 8294 22090 8432
rect 21902 8208 21914 8294
rect 22078 8208 22090 8294
rect 21902 8070 22090 8208
rect 21902 7984 21914 8070
rect 22078 7984 22090 8070
rect 21902 7846 22090 7984
rect 21902 7760 21914 7846
rect 22078 7760 22090 7846
rect 21902 7622 22090 7760
rect 21902 7536 21914 7622
rect 22078 7536 22090 7622
rect 21902 7398 22090 7536
rect 21902 7312 21914 7398
rect 22078 7312 22090 7398
rect 21902 6486 22090 7312
rect 21902 6400 21914 6486
rect 22078 6400 22090 6486
rect 21902 6262 22090 6400
rect 21902 6176 21914 6262
rect 22078 6176 22090 6262
rect 21902 6038 22090 6176
rect 21902 5952 21914 6038
rect 22078 5952 22090 6038
rect 21902 5814 22090 5952
rect 21902 5728 21914 5814
rect 22078 5728 22090 5814
rect 21902 5590 22090 5728
rect 21902 5504 21914 5590
rect 22078 5504 22090 5590
rect 21902 5366 22090 5504
rect 21902 5280 21914 5366
rect 22078 5280 22090 5366
rect 1737 5016 1818 5053
rect 21902 5142 22090 5280
rect 21902 5056 21914 5142
rect 22078 5056 22090 5142
rect 21902 5045 22090 5056
rect 22150 8616 31550 8679
rect 22150 8564 22165 8616
rect 31539 8564 31550 8616
rect 22150 8168 31550 8564
rect 22150 8116 22168 8168
rect 31542 8116 31550 8168
rect 22150 7720 31550 8116
rect 22150 7668 22166 7720
rect 31540 7668 31550 7720
rect 22150 7272 31550 7668
rect 22150 7220 22168 7272
rect 31542 7220 31550 7272
rect 22150 6360 31550 7220
rect 22150 6308 22164 6360
rect 31538 6308 31550 6360
rect 22150 5912 31550 6308
rect 22150 5860 22165 5912
rect 31539 5860 31550 5912
rect 22150 5464 31550 5860
rect 22150 5412 22163 5464
rect 31537 5412 31550 5464
rect 22150 5016 31550 5412
rect 32627 8404 42028 8788
rect 32627 8340 32646 8404
rect 42012 8340 42028 8404
rect 32627 7956 42028 8340
rect 32627 7892 32643 7956
rect 42009 7892 42028 7956
rect 32627 7508 42028 7892
rect 32627 7444 32639 7508
rect 42005 7444 42028 7508
rect 32627 7116 42028 7444
rect 32627 6532 32640 7116
rect 42006 6532 42028 7116
rect 32627 6148 42028 6532
rect 32627 6084 32645 6148
rect 42011 6084 42028 6148
rect 32627 5700 42028 6084
rect 32627 5636 32646 5700
rect 42012 5636 42028 5700
rect 32627 5252 42028 5636
rect 32627 5188 32644 5252
rect 42010 5188 42028 5252
rect 32627 5176 42028 5188
rect 42134 8742 42322 8947
rect 42134 8656 42146 8742
rect 42310 8656 42322 8742
rect 62396 8739 62477 8947
rect 42134 8518 42322 8656
rect 42134 8432 42146 8518
rect 42310 8432 42322 8518
rect 42134 8294 42322 8432
rect 42134 8208 42146 8294
rect 42310 8208 42322 8294
rect 42134 8070 42322 8208
rect 42134 7984 42146 8070
rect 42310 7984 42322 8070
rect 42134 7846 42322 7984
rect 42134 7760 42146 7846
rect 42310 7760 42322 7846
rect 42134 7622 42322 7760
rect 42134 7536 42146 7622
rect 42310 7536 42322 7622
rect 42134 7398 42322 7536
rect 42134 7312 42146 7398
rect 42310 7312 42322 7398
rect 42134 6486 42322 7312
rect 42134 6400 42146 6486
rect 42310 6400 42322 6486
rect 42134 6262 42322 6400
rect 42134 6176 42146 6262
rect 42310 6176 42322 6262
rect 42134 6038 42322 6176
rect 42134 5952 42146 6038
rect 42310 5952 42322 6038
rect 42134 5814 42322 5952
rect 42134 5728 42146 5814
rect 42310 5728 42322 5814
rect 42134 5590 42322 5728
rect 42134 5504 42146 5590
rect 42310 5504 42322 5590
rect 42134 5366 42322 5504
rect 42134 5280 42146 5366
rect 42310 5280 42322 5366
rect 42134 5142 42322 5280
rect 42134 5056 42146 5142
rect 42310 5056 42322 5142
rect 42134 5046 42322 5056
rect 42392 8616 62299 8679
rect 42392 8564 42416 8616
rect 62262 8564 62299 8616
rect 42392 8168 62299 8564
rect 42392 8116 42417 8168
rect 62263 8116 62299 8168
rect 42392 7720 62299 8116
rect 42392 7668 42418 7720
rect 62264 7668 62299 7720
rect 42392 7272 62299 7668
rect 42392 7220 42413 7272
rect 62259 7220 62299 7272
rect 42392 6360 62299 7220
rect 42392 6308 42421 6360
rect 62267 6308 62299 6360
rect 42392 5912 62299 6308
rect 42392 5860 42426 5912
rect 62272 5860 62299 5912
rect 42392 5464 62299 5860
rect 42392 5412 42428 5464
rect 62274 5412 62299 5464
rect 22150 4964 22165 5016
rect 31539 4990 31550 5016
rect 42392 5016 62299 5412
rect 42392 4990 42419 5016
rect 31539 4964 42419 4990
rect 62265 4964 62299 5016
rect 62396 7309 62407 8739
rect 62459 7309 62477 8739
rect 62396 6489 62477 7309
rect 62396 5053 62407 6489
rect 62459 5053 62477 6489
rect 62396 5008 62477 5053
rect 22150 4482 62299 4964
rect 1883 4374 21825 4408
rect 1883 4322 1901 4374
rect 21823 4322 21825 4374
rect 1691 4279 1814 4305
rect 1691 3995 1758 4279
rect 1275 3437 1758 3995
rect 1275 3114 1290 3437
rect 1215 3106 1290 3114
rect 704 3049 1056 3056
rect 562 2991 1169 2993
rect 562 2899 1105 2991
rect 423 2392 506 2800
rect 1075 2764 1105 2899
rect 1066 2759 1105 2764
rect 1157 2764 1169 2991
rect 1691 2843 1758 3437
rect 1810 2843 1814 4279
rect 1157 2759 1200 2764
rect 1066 2703 1088 2759
rect 1180 2703 1200 2759
rect 1066 2696 1200 2703
rect 423 2309 709 2392
rect 626 2258 709 2309
rect 626 1301 647 2258
rect 699 1388 709 2258
rect 1369 2120 1444 2128
rect 699 1380 1313 1388
rect 699 1301 1251 1380
rect 626 1293 1251 1301
rect 1234 882 1251 1293
rect 1303 882 1313 1380
rect 1234 874 1313 882
rect 1369 449 1378 2120
rect 1430 2078 1444 2120
rect 1691 2078 1814 2843
rect 1430 2023 1814 2078
rect 1430 1520 1758 2023
rect 1430 449 1444 1520
rect 1369 441 1444 449
rect 1691 587 1758 1520
rect 1810 587 1814 2023
rect 1883 3926 21825 4322
rect 1883 3874 1907 3926
rect 21823 3874 21825 3926
rect 1883 3478 21825 3874
rect 1883 3426 1909 3478
rect 21823 3426 21825 3478
rect 1883 3030 21825 3426
rect 1883 2978 1905 3030
rect 21823 2978 21825 3030
rect 1883 2649 21825 2978
rect 1883 2066 1899 2649
rect 21823 2066 21825 2649
rect 1883 1670 21825 2066
rect 1883 1618 1903 1670
rect 21823 1618 21825 1670
rect 1883 1222 21825 1618
rect 1883 1170 1903 1222
rect 21823 1170 21825 1222
rect 1883 774 21825 1170
rect 1883 722 1891 774
rect 21815 722 21825 774
rect 1883 707 21825 722
rect 21899 4276 22087 4311
rect 21899 4190 21911 4276
rect 22075 4190 22087 4276
rect 21899 4052 22087 4190
rect 21899 3966 21911 4052
rect 22075 3966 22087 4052
rect 21899 3828 22087 3966
rect 21899 3742 21911 3828
rect 22075 3742 22087 3828
rect 21899 3604 22087 3742
rect 21899 3518 21911 3604
rect 22075 3518 22087 3604
rect 21899 3380 22087 3518
rect 21899 3294 21911 3380
rect 22075 3294 22087 3380
rect 21899 3156 22087 3294
rect 21899 3070 21911 3156
rect 22075 3070 22087 3156
rect 21899 2932 22087 3070
rect 21899 2846 21911 2932
rect 22075 2846 22087 2932
rect 21899 2020 22087 2846
rect 21899 1934 21911 2020
rect 22075 1934 22087 2020
rect 21899 1796 22087 1934
rect 21899 1710 21911 1796
rect 22075 1710 22087 1796
rect 21899 1572 22087 1710
rect 21899 1486 21911 1572
rect 22075 1486 22087 1572
rect 21899 1348 22087 1486
rect 21899 1262 21911 1348
rect 22075 1262 22087 1348
rect 21899 1124 22087 1262
rect 21899 1038 21911 1124
rect 22075 1038 22087 1124
rect 21899 900 22087 1038
rect 21899 814 21911 900
rect 22075 814 22087 900
rect 1691 423 1814 587
rect 21899 676 22087 814
rect 21899 590 21911 676
rect 22075 590 22087 676
rect 21899 423 22087 590
rect 22150 4150 31550 4482
rect 22150 4098 22171 4150
rect 31545 4098 31550 4150
rect 22150 3702 31550 4098
rect 22150 3650 22170 3702
rect 31544 3650 31550 3702
rect 22150 3254 31550 3650
rect 22150 3202 22167 3254
rect 31541 3202 31550 3254
rect 22150 2807 31550 3202
rect 22150 2755 22168 2807
rect 31542 2755 31550 2807
rect 22150 1894 31550 2755
rect 22150 1842 22170 1894
rect 31544 1842 31550 1894
rect 22150 1446 31550 1842
rect 22150 1394 22171 1446
rect 31545 1394 31550 1446
rect 22150 998 31550 1394
rect 22150 946 22167 998
rect 31541 946 31550 998
rect 22150 550 31550 946
rect 32651 4387 42052 4396
rect 32651 4322 32662 4387
rect 42028 4322 42052 4387
rect 32651 3939 42052 4322
rect 32651 3874 32664 3939
rect 42030 3874 42052 3939
rect 32651 3491 42052 3874
rect 32651 3426 32664 3491
rect 42030 3426 42052 3491
rect 32651 3043 42052 3426
rect 32651 2978 32663 3043
rect 42029 2978 42052 3043
rect 32651 2650 42052 2978
rect 32651 2066 32659 2650
rect 42025 2131 42052 2650
rect 42026 2066 42052 2131
rect 32651 1683 42052 2066
rect 32651 1618 32665 1683
rect 42031 1618 42052 1683
rect 32651 1235 42052 1618
rect 32651 1170 32675 1235
rect 42041 1170 42052 1235
rect 32651 787 42052 1170
rect 32651 722 32658 787
rect 42024 722 42052 787
rect 32651 700 42052 722
rect 42131 4276 42319 4310
rect 42131 4190 42143 4276
rect 42307 4190 42319 4276
rect 42131 4052 42319 4190
rect 42131 3966 42143 4052
rect 42307 3966 42319 4052
rect 42131 3828 42319 3966
rect 42131 3742 42143 3828
rect 42307 3742 42319 3828
rect 42131 3604 42319 3742
rect 42131 3518 42143 3604
rect 42307 3518 42319 3604
rect 42131 3380 42319 3518
rect 42131 3294 42143 3380
rect 42307 3294 42319 3380
rect 42131 3156 42319 3294
rect 42131 3070 42143 3156
rect 42307 3070 42319 3156
rect 42131 2932 42319 3070
rect 42131 2846 42143 2932
rect 42307 2846 42319 2932
rect 42131 2020 42319 2846
rect 42131 1934 42143 2020
rect 42307 1934 42319 2020
rect 42131 1796 42319 1934
rect 42131 1710 42143 1796
rect 42307 1710 42319 1796
rect 42131 1572 42319 1710
rect 42131 1486 42143 1572
rect 42307 1486 42319 1572
rect 42131 1348 42319 1486
rect 42131 1262 42143 1348
rect 42307 1262 42319 1348
rect 42131 1124 42319 1262
rect 42131 1038 42143 1124
rect 42307 1038 42319 1124
rect 42131 900 42319 1038
rect 42131 814 42143 900
rect 42307 814 42319 900
rect 22150 498 22164 550
rect 31538 498 31550 550
rect 22150 483 31550 498
rect 42131 676 42319 814
rect 42131 590 42143 676
rect 42307 590 42319 676
rect 42131 423 42319 590
rect 42392 4150 62299 4482
rect 42392 4098 42417 4150
rect 62263 4098 62299 4150
rect 42392 3702 62299 4098
rect 42392 3650 42421 3702
rect 62267 3650 62299 3702
rect 42392 3254 62299 3650
rect 42392 3202 42423 3254
rect 62269 3202 62299 3254
rect 42392 2806 62299 3202
rect 42392 2754 42418 2806
rect 62264 2754 62299 2806
rect 42392 1894 62299 2754
rect 42392 1842 42416 1894
rect 62262 1842 62299 1894
rect 42392 1446 62299 1842
rect 42392 1394 42417 1446
rect 62263 1394 62299 1446
rect 42392 998 62299 1394
rect 42392 946 42422 998
rect 62268 946 62299 998
rect 42392 550 62299 946
rect 42392 498 42413 550
rect 62259 498 62299 550
rect 42392 483 62299 498
rect 62401 4279 62482 4305
rect 62401 2843 62408 4279
rect 62460 2843 62482 4279
rect 62401 2023 62482 2843
rect 62401 587 62408 2023
rect 62460 587 62482 2023
rect 62401 423 62482 587
rect 1691 300 62482 423
use pfet_06v0_5JTQE2  XM1
timestamp 1762867378
transform 0 1 32112 -1 0 8027
box -996 -30488 996 30488
use pfet_06v0_E9HJGY  XM2
timestamp 1762867378
transform 1 0 1268 0 1 7368
box -324 -1656 324 1656
use nfet_06v0_AQU3CZ  XM3
timestamp 1762867098
transform 0 1 32109 -1 0 3561
box -996 -30488 996 30488
use pfet_06v0_E9HJGY  XM9
timestamp 1762867378
transform 1 0 756 0 1 7368
box -324 -1656 324 1656
use pfet_06v0_5JTQE2  XM10
timestamp 1762867378
transform 0 1 32112 -1 0 5771
box -996 -30488 996 30488
use pfet_06v0_E9HJGY  XM11
timestamp 1762867378
transform 1 0 622 0 1 4192
box -324 -1656 324 1656
use pfet_06v0_E9HJGY  XM12
timestamp 1762867378
transform 1 0 1134 0 1 4192
box -324 -1656 324 1656
use nfet_06v0_6KT3L3  XM13
timestamp 1762867378
transform 1 0 777 0 1 1272
box -324 -1256 324 1256
use nfet_06v0_6KT3L3  XM14
timestamp 1762867378
transform 1 0 1289 0 1 1272
box -324 -1256 324 1256
use nfet_06v0_AQU3CZ  XM15
timestamp 1762867098
transform 0 1 32109 -1 0 1305
box -996 -30488 996 30488
<< labels >>
flabel metal2 0 4267 286 4352 0 FreeSans 200 0 0 0 PLUS
port 1 nsew signal input
flabel metal2 0 5097 286 5182 0 FreeSans 200 0 0 0 MINUS
port 2 nsew signal input
flabel metal2 0 8799 286 8884 0 FreeSans 200 0 0 0 ADJ
port 3 nsew signal input
flabel metal1 298 9122 62677 9333 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 1613 0 62677 211 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal2 42392 483 62299 8679 0 FreeSans 200 0 0 0 OUT
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 62677 9333
<< end >>
