magic
tech gf180mcuD
magscale 1 10
timestamp 1763836631
<< nwell >>
rect 2266 4675 64645 9333
rect 2266 2536 3512 4675
<< pwell >>
rect 335 10276 11290 11672
rect 11291 10276 12913 11672
rect 335 9465 12913 10276
rect 335 2536 2266 9465
rect 3512 2536 64645 4675
rect 335 0 64645 2536
<< mvnmos >>
rect 3845 4173 23845 4293
rect 24077 4173 44077 4293
rect 44309 4173 64309 4293
rect 3845 3949 23845 4069
rect 24077 3949 44077 4069
rect 44309 3949 64309 4069
rect 3845 3725 23845 3845
rect 24077 3725 44077 3845
rect 44309 3725 64309 3845
rect 3845 3501 23845 3621
rect 24077 3501 44077 3621
rect 44309 3501 64309 3621
rect 3845 3277 23845 3397
rect 24077 3277 44077 3397
rect 44309 3277 64309 3397
rect 3845 3053 23845 3173
rect 24077 3053 44077 3173
rect 44309 3053 64309 3173
rect 3845 2829 23845 2949
rect 24077 2829 44077 2949
rect 44309 2829 64309 2949
rect 2685 272 2805 2272
rect 3197 272 3317 2272
rect 3845 1917 23845 2037
rect 24077 1917 44077 2037
rect 44309 1917 64309 2037
rect 3845 1693 23845 1813
rect 24077 1693 44077 1813
rect 44309 1693 64309 1813
rect 3845 1469 23845 1589
rect 24077 1469 44077 1589
rect 44309 1469 64309 1589
rect 3845 1245 23845 1365
rect 24077 1245 44077 1365
rect 44309 1245 64309 1365
rect 3845 1021 23845 1141
rect 24077 1021 44077 1141
rect 44309 1021 64309 1141
rect 3845 797 23845 917
rect 24077 797 44077 917
rect 44309 797 64309 917
rect 3845 573 23845 693
rect 24077 573 44077 693
rect 44309 573 64309 693
<< mvpmos >>
rect 2664 5968 2784 8768
rect 3176 5968 3296 8768
rect 3848 8639 23848 8759
rect 24080 8639 44080 8759
rect 44312 8639 64312 8759
rect 3848 8415 23848 8535
rect 24080 8415 44080 8535
rect 44312 8415 64312 8535
rect 3848 8191 23848 8311
rect 24080 8191 44080 8311
rect 44312 8191 64312 8311
rect 3848 7967 23848 8087
rect 24080 7967 44080 8087
rect 44312 7967 64312 8087
rect 3848 7743 23848 7863
rect 24080 7743 44080 7863
rect 44312 7743 64312 7863
rect 3848 7519 23848 7639
rect 24080 7519 44080 7639
rect 44312 7519 64312 7639
rect 3848 7295 23848 7415
rect 24080 7295 44080 7415
rect 44312 7295 64312 7415
rect 3848 6383 23848 6503
rect 24080 6383 44080 6503
rect 44312 6383 64312 6503
rect 3848 6159 23848 6279
rect 24080 6159 44080 6279
rect 44312 6159 64312 6279
rect 3848 5935 23848 6055
rect 24080 5935 44080 6055
rect 44312 5935 64312 6055
rect 2530 2792 2650 5592
rect 3042 2792 3162 5592
rect 3848 5711 23848 5831
rect 24080 5711 44080 5831
rect 44312 5711 64312 5831
rect 3848 5487 23848 5607
rect 24080 5487 44080 5607
rect 44312 5487 64312 5607
rect 3848 5263 23848 5383
rect 24080 5263 44080 5383
rect 44312 5263 64312 5383
rect 3848 5039 23848 5159
rect 24080 5039 44080 5159
rect 44312 5039 64312 5159
<< mvndiff >>
rect 3845 4368 23845 4381
rect 3845 4322 3858 4368
rect 23832 4322 23845 4368
rect 3845 4293 23845 4322
rect 24077 4368 44077 4381
rect 24077 4322 24090 4368
rect 44064 4322 44077 4368
rect 24077 4293 44077 4322
rect 44309 4368 64309 4381
rect 44309 4322 44322 4368
rect 64296 4322 64309 4368
rect 44309 4293 64309 4322
rect 3845 4144 23845 4173
rect 3845 4098 3858 4144
rect 23832 4098 23845 4144
rect 3845 4069 23845 4098
rect 24077 4144 44077 4173
rect 24077 4098 24090 4144
rect 44064 4098 44077 4144
rect 24077 4069 44077 4098
rect 44309 4144 64309 4173
rect 44309 4098 44322 4144
rect 64296 4098 64309 4144
rect 44309 4069 64309 4098
rect 3845 3920 23845 3949
rect 3845 3874 3858 3920
rect 23832 3874 23845 3920
rect 3845 3845 23845 3874
rect 24077 3920 44077 3949
rect 24077 3874 24090 3920
rect 44064 3874 44077 3920
rect 24077 3845 44077 3874
rect 44309 3920 64309 3949
rect 44309 3874 44322 3920
rect 64296 3874 64309 3920
rect 44309 3845 64309 3874
rect 3845 3696 23845 3725
rect 3845 3650 3858 3696
rect 23832 3650 23845 3696
rect 3845 3621 23845 3650
rect 24077 3696 44077 3725
rect 24077 3650 24090 3696
rect 44064 3650 44077 3696
rect 24077 3621 44077 3650
rect 44309 3696 64309 3725
rect 44309 3650 44322 3696
rect 64296 3650 64309 3696
rect 44309 3621 64309 3650
rect 3845 3472 23845 3501
rect 3845 3426 3858 3472
rect 23832 3426 23845 3472
rect 3845 3397 23845 3426
rect 24077 3472 44077 3501
rect 24077 3426 24090 3472
rect 44064 3426 44077 3472
rect 24077 3397 44077 3426
rect 44309 3472 64309 3501
rect 44309 3426 44322 3472
rect 64296 3426 64309 3472
rect 44309 3397 64309 3426
rect 3845 3248 23845 3277
rect 3845 3202 3858 3248
rect 23832 3202 23845 3248
rect 3845 3173 23845 3202
rect 24077 3248 44077 3277
rect 24077 3202 24090 3248
rect 44064 3202 44077 3248
rect 24077 3173 44077 3202
rect 44309 3248 64309 3277
rect 44309 3202 44322 3248
rect 64296 3202 64309 3248
rect 44309 3173 64309 3202
rect 3845 3024 23845 3053
rect 3845 2978 3858 3024
rect 23832 2978 23845 3024
rect 3845 2949 23845 2978
rect 24077 3024 44077 3053
rect 24077 2978 24090 3024
rect 44064 2978 44077 3024
rect 24077 2949 44077 2978
rect 44309 3024 64309 3053
rect 44309 2978 44322 3024
rect 64296 2978 64309 3024
rect 44309 2949 64309 2978
rect 3845 2800 23845 2829
rect 3845 2754 3858 2800
rect 23832 2754 23845 2800
rect 3845 2741 23845 2754
rect 24077 2800 44077 2829
rect 24077 2754 24090 2800
rect 44064 2754 44077 2800
rect 24077 2741 44077 2754
rect 44309 2800 64309 2829
rect 44309 2754 44322 2800
rect 64296 2754 64309 2800
rect 44309 2741 64309 2754
rect 2597 2259 2685 2272
rect 2597 285 2610 2259
rect 2656 285 2685 2259
rect 2597 272 2685 285
rect 2805 2259 2893 2272
rect 2805 285 2834 2259
rect 2880 285 2893 2259
rect 2805 272 2893 285
rect 3109 2259 3197 2272
rect 3109 285 3122 2259
rect 3168 285 3197 2259
rect 3109 272 3197 285
rect 3317 2259 3405 2272
rect 3317 285 3346 2259
rect 3392 285 3405 2259
rect 3317 272 3405 285
rect 3845 2112 23845 2125
rect 3845 2066 3858 2112
rect 23832 2066 23845 2112
rect 3845 2037 23845 2066
rect 24077 2112 44077 2125
rect 24077 2066 24090 2112
rect 44064 2066 44077 2112
rect 24077 2037 44077 2066
rect 44309 2112 64309 2125
rect 44309 2066 44322 2112
rect 64296 2066 64309 2112
rect 44309 2037 64309 2066
rect 3845 1888 23845 1917
rect 3845 1842 3858 1888
rect 23832 1842 23845 1888
rect 3845 1813 23845 1842
rect 24077 1888 44077 1917
rect 24077 1842 24090 1888
rect 44064 1842 44077 1888
rect 24077 1813 44077 1842
rect 44309 1888 64309 1917
rect 44309 1842 44322 1888
rect 64296 1842 64309 1888
rect 44309 1813 64309 1842
rect 3845 1664 23845 1693
rect 3845 1618 3858 1664
rect 23832 1618 23845 1664
rect 3845 1589 23845 1618
rect 24077 1664 44077 1693
rect 24077 1618 24090 1664
rect 44064 1618 44077 1664
rect 24077 1589 44077 1618
rect 44309 1664 64309 1693
rect 44309 1618 44322 1664
rect 64296 1618 64309 1664
rect 44309 1589 64309 1618
rect 3845 1440 23845 1469
rect 3845 1394 3858 1440
rect 23832 1394 23845 1440
rect 3845 1365 23845 1394
rect 24077 1440 44077 1469
rect 24077 1394 24090 1440
rect 44064 1394 44077 1440
rect 24077 1365 44077 1394
rect 44309 1440 64309 1469
rect 44309 1394 44322 1440
rect 64296 1394 64309 1440
rect 44309 1365 64309 1394
rect 3845 1216 23845 1245
rect 3845 1170 3858 1216
rect 23832 1170 23845 1216
rect 3845 1141 23845 1170
rect 24077 1216 44077 1245
rect 24077 1170 24090 1216
rect 44064 1170 44077 1216
rect 24077 1141 44077 1170
rect 44309 1216 64309 1245
rect 44309 1170 44322 1216
rect 64296 1170 64309 1216
rect 44309 1141 64309 1170
rect 3845 992 23845 1021
rect 3845 946 3858 992
rect 23832 946 23845 992
rect 3845 917 23845 946
rect 24077 992 44077 1021
rect 24077 946 24090 992
rect 44064 946 44077 992
rect 24077 917 44077 946
rect 44309 992 64309 1021
rect 44309 946 44322 992
rect 64296 946 64309 992
rect 44309 917 64309 946
rect 3845 768 23845 797
rect 3845 722 3858 768
rect 23832 722 23845 768
rect 3845 693 23845 722
rect 24077 768 44077 797
rect 24077 722 24090 768
rect 44064 722 44077 768
rect 24077 693 44077 722
rect 44309 768 64309 797
rect 44309 722 44322 768
rect 64296 722 64309 768
rect 44309 693 64309 722
rect 3845 544 23845 573
rect 3845 498 3858 544
rect 23832 498 23845 544
rect 3845 485 23845 498
rect 24077 544 44077 573
rect 24077 498 24090 544
rect 44064 498 44077 544
rect 24077 485 44077 498
rect 44309 544 64309 573
rect 44309 498 44322 544
rect 64296 498 64309 544
rect 44309 485 64309 498
<< mvpdiff >>
rect 2576 8755 2664 8768
rect 2576 5981 2589 8755
rect 2635 5981 2664 8755
rect 2576 5968 2664 5981
rect 2784 8755 2872 8768
rect 2784 5981 2813 8755
rect 2859 5981 2872 8755
rect 2784 5968 2872 5981
rect 3088 8755 3176 8768
rect 3088 5981 3101 8755
rect 3147 5981 3176 8755
rect 3088 5968 3176 5981
rect 3296 8755 3384 8768
rect 3296 5981 3325 8755
rect 3371 5981 3384 8755
rect 3296 5968 3384 5981
rect 3848 8834 23848 8847
rect 3848 8788 3861 8834
rect 23835 8788 23848 8834
rect 3848 8759 23848 8788
rect 24080 8834 44080 8847
rect 24080 8788 24093 8834
rect 44067 8788 44080 8834
rect 24080 8759 44080 8788
rect 44312 8834 64312 8847
rect 44312 8788 44325 8834
rect 64299 8788 64312 8834
rect 44312 8759 64312 8788
rect 3848 8610 23848 8639
rect 3848 8564 3861 8610
rect 23835 8564 23848 8610
rect 3848 8535 23848 8564
rect 24080 8610 44080 8639
rect 24080 8564 24093 8610
rect 44067 8564 44080 8610
rect 24080 8535 44080 8564
rect 44312 8610 64312 8639
rect 44312 8564 44325 8610
rect 64299 8564 64312 8610
rect 44312 8535 64312 8564
rect 3848 8386 23848 8415
rect 3848 8340 3861 8386
rect 23835 8340 23848 8386
rect 3848 8311 23848 8340
rect 24080 8386 44080 8415
rect 24080 8340 24093 8386
rect 44067 8340 44080 8386
rect 24080 8311 44080 8340
rect 44312 8386 64312 8415
rect 44312 8340 44325 8386
rect 64299 8340 64312 8386
rect 44312 8311 64312 8340
rect 3848 8162 23848 8191
rect 3848 8116 3861 8162
rect 23835 8116 23848 8162
rect 3848 8087 23848 8116
rect 24080 8162 44080 8191
rect 24080 8116 24093 8162
rect 44067 8116 44080 8162
rect 24080 8087 44080 8116
rect 44312 8162 64312 8191
rect 44312 8116 44325 8162
rect 64299 8116 64312 8162
rect 44312 8087 64312 8116
rect 3848 7938 23848 7967
rect 3848 7892 3861 7938
rect 23835 7892 23848 7938
rect 3848 7863 23848 7892
rect 24080 7938 44080 7967
rect 24080 7892 24093 7938
rect 44067 7892 44080 7938
rect 24080 7863 44080 7892
rect 44312 7938 64312 7967
rect 44312 7892 44325 7938
rect 64299 7892 64312 7938
rect 44312 7863 64312 7892
rect 3848 7714 23848 7743
rect 3848 7668 3861 7714
rect 23835 7668 23848 7714
rect 3848 7639 23848 7668
rect 24080 7714 44080 7743
rect 24080 7668 24093 7714
rect 44067 7668 44080 7714
rect 24080 7639 44080 7668
rect 44312 7714 64312 7743
rect 44312 7668 44325 7714
rect 64299 7668 64312 7714
rect 44312 7639 64312 7668
rect 3848 7490 23848 7519
rect 3848 7444 3861 7490
rect 23835 7444 23848 7490
rect 3848 7415 23848 7444
rect 24080 7490 44080 7519
rect 24080 7444 24093 7490
rect 44067 7444 44080 7490
rect 24080 7415 44080 7444
rect 44312 7490 64312 7519
rect 44312 7444 44325 7490
rect 64299 7444 64312 7490
rect 44312 7415 64312 7444
rect 3848 7266 23848 7295
rect 3848 7220 3861 7266
rect 23835 7220 23848 7266
rect 3848 7207 23848 7220
rect 24080 7266 44080 7295
rect 24080 7220 24093 7266
rect 44067 7220 44080 7266
rect 24080 7207 44080 7220
rect 44312 7266 64312 7295
rect 44312 7220 44325 7266
rect 64299 7220 64312 7266
rect 44312 7207 64312 7220
rect 3848 6578 23848 6591
rect 3848 6532 3861 6578
rect 23835 6532 23848 6578
rect 3848 6503 23848 6532
rect 24080 6578 44080 6591
rect 24080 6532 24093 6578
rect 44067 6532 44080 6578
rect 24080 6503 44080 6532
rect 44312 6578 64312 6591
rect 44312 6532 44325 6578
rect 64299 6532 64312 6578
rect 44312 6503 64312 6532
rect 3848 6354 23848 6383
rect 3848 6308 3861 6354
rect 23835 6308 23848 6354
rect 3848 6279 23848 6308
rect 24080 6354 44080 6383
rect 24080 6308 24093 6354
rect 44067 6308 44080 6354
rect 24080 6279 44080 6308
rect 44312 6354 64312 6383
rect 44312 6308 44325 6354
rect 64299 6308 64312 6354
rect 44312 6279 64312 6308
rect 3848 6130 23848 6159
rect 3848 6084 3861 6130
rect 23835 6084 23848 6130
rect 3848 6055 23848 6084
rect 24080 6130 44080 6159
rect 24080 6084 24093 6130
rect 44067 6084 44080 6130
rect 24080 6055 44080 6084
rect 44312 6130 64312 6159
rect 44312 6084 44325 6130
rect 64299 6084 64312 6130
rect 44312 6055 64312 6084
rect 3848 5906 23848 5935
rect 3848 5860 3861 5906
rect 23835 5860 23848 5906
rect 3848 5831 23848 5860
rect 24080 5906 44080 5935
rect 24080 5860 24093 5906
rect 44067 5860 44080 5906
rect 24080 5831 44080 5860
rect 44312 5906 64312 5935
rect 44312 5860 44325 5906
rect 64299 5860 64312 5906
rect 44312 5831 64312 5860
rect 2442 5579 2530 5592
rect 2442 2805 2455 5579
rect 2501 2805 2530 5579
rect 2442 2792 2530 2805
rect 2650 5579 2738 5592
rect 2650 2805 2679 5579
rect 2725 2805 2738 5579
rect 2650 2792 2738 2805
rect 2954 5579 3042 5592
rect 2954 2805 2967 5579
rect 3013 2805 3042 5579
rect 2954 2792 3042 2805
rect 3162 5579 3250 5592
rect 3162 2805 3191 5579
rect 3237 2805 3250 5579
rect 3162 2792 3250 2805
rect 3848 5682 23848 5711
rect 3848 5636 3861 5682
rect 23835 5636 23848 5682
rect 3848 5607 23848 5636
rect 24080 5682 44080 5711
rect 24080 5636 24093 5682
rect 44067 5636 44080 5682
rect 24080 5607 44080 5636
rect 44312 5682 64312 5711
rect 44312 5636 44325 5682
rect 64299 5636 64312 5682
rect 44312 5607 64312 5636
rect 3848 5458 23848 5487
rect 3848 5412 3861 5458
rect 23835 5412 23848 5458
rect 3848 5383 23848 5412
rect 24080 5458 44080 5487
rect 24080 5412 24093 5458
rect 44067 5412 44080 5458
rect 24080 5383 44080 5412
rect 44312 5458 64312 5487
rect 44312 5412 44325 5458
rect 64299 5412 64312 5458
rect 44312 5383 64312 5412
rect 3848 5234 23848 5263
rect 3848 5188 3861 5234
rect 23835 5188 23848 5234
rect 3848 5159 23848 5188
rect 24080 5234 44080 5263
rect 24080 5188 24093 5234
rect 44067 5188 44080 5234
rect 24080 5159 44080 5188
rect 44312 5234 64312 5263
rect 44312 5188 44325 5234
rect 64299 5188 64312 5234
rect 44312 5159 64312 5188
rect 3848 5010 23848 5039
rect 3848 4964 3861 5010
rect 23835 4964 23848 5010
rect 3848 4951 23848 4964
rect 24080 5010 44080 5039
rect 24080 4964 24093 5010
rect 44067 4964 44080 5010
rect 24080 4951 44080 4964
rect 44312 5010 64312 5039
rect 44312 4964 44325 5010
rect 64299 4964 64312 5010
rect 44312 4951 64312 4964
<< mvndiffc >>
rect 3858 4322 23832 4368
rect 24090 4322 44064 4368
rect 44322 4322 64296 4368
rect 3858 4098 23832 4144
rect 24090 4098 44064 4144
rect 44322 4098 64296 4144
rect 3858 3874 23832 3920
rect 24090 3874 44064 3920
rect 44322 3874 64296 3920
rect 3858 3650 23832 3696
rect 24090 3650 44064 3696
rect 44322 3650 64296 3696
rect 3858 3426 23832 3472
rect 24090 3426 44064 3472
rect 44322 3426 64296 3472
rect 3858 3202 23832 3248
rect 24090 3202 44064 3248
rect 44322 3202 64296 3248
rect 3858 2978 23832 3024
rect 24090 2978 44064 3024
rect 44322 2978 64296 3024
rect 3858 2754 23832 2800
rect 24090 2754 44064 2800
rect 44322 2754 64296 2800
rect 2610 285 2656 2259
rect 2834 285 2880 2259
rect 3122 285 3168 2259
rect 3346 285 3392 2259
rect 3858 2066 23832 2112
rect 24090 2066 44064 2112
rect 44322 2066 64296 2112
rect 3858 1842 23832 1888
rect 24090 1842 44064 1888
rect 44322 1842 64296 1888
rect 3858 1618 23832 1664
rect 24090 1618 44064 1664
rect 44322 1618 64296 1664
rect 3858 1394 23832 1440
rect 24090 1394 44064 1440
rect 44322 1394 64296 1440
rect 3858 1170 23832 1216
rect 24090 1170 44064 1216
rect 44322 1170 64296 1216
rect 3858 946 23832 992
rect 24090 946 44064 992
rect 44322 946 64296 992
rect 3858 722 23832 768
rect 24090 722 44064 768
rect 44322 722 64296 768
rect 3858 498 23832 544
rect 24090 498 44064 544
rect 44322 498 64296 544
<< mvpdiffc >>
rect 2589 5981 2635 8755
rect 2813 5981 2859 8755
rect 3101 5981 3147 8755
rect 3325 5981 3371 8755
rect 3861 8788 23835 8834
rect 24093 8788 44067 8834
rect 44325 8788 64299 8834
rect 3861 8564 23835 8610
rect 24093 8564 44067 8610
rect 44325 8564 64299 8610
rect 3861 8340 23835 8386
rect 24093 8340 44067 8386
rect 44325 8340 64299 8386
rect 3861 8116 23835 8162
rect 24093 8116 44067 8162
rect 44325 8116 64299 8162
rect 3861 7892 23835 7938
rect 24093 7892 44067 7938
rect 44325 7892 64299 7938
rect 3861 7668 23835 7714
rect 24093 7668 44067 7714
rect 44325 7668 64299 7714
rect 3861 7444 23835 7490
rect 24093 7444 44067 7490
rect 44325 7444 64299 7490
rect 3861 7220 23835 7266
rect 24093 7220 44067 7266
rect 44325 7220 64299 7266
rect 3861 6532 23835 6578
rect 24093 6532 44067 6578
rect 44325 6532 64299 6578
rect 3861 6308 23835 6354
rect 24093 6308 44067 6354
rect 44325 6308 64299 6354
rect 3861 6084 23835 6130
rect 24093 6084 44067 6130
rect 44325 6084 64299 6130
rect 3861 5860 23835 5906
rect 24093 5860 44067 5906
rect 44325 5860 64299 5906
rect 2455 2805 2501 5579
rect 2679 2805 2725 5579
rect 2967 2805 3013 5579
rect 3191 2805 3237 5579
rect 3861 5636 23835 5682
rect 24093 5636 44067 5682
rect 44325 5636 64299 5682
rect 3861 5412 23835 5458
rect 24093 5412 44067 5458
rect 44325 5412 64299 5458
rect 3861 5188 23835 5234
rect 24093 5188 44067 5234
rect 44325 5188 64299 5234
rect 3861 4964 23835 5010
rect 24093 4964 44067 5010
rect 44325 4964 64299 5010
<< mvpsubdiff >>
rect 367 11568 991 11640
rect 367 11524 439 11568
rect 367 10288 380 11524
rect 426 10288 439 11524
rect 919 11524 991 11568
rect 367 10244 439 10288
rect 919 10288 932 11524
rect 978 10288 991 11524
rect 919 10244 991 10288
rect 1363 11568 1987 11640
rect 1363 11524 1435 11568
rect 1363 10288 1376 11524
rect 1422 10288 1435 11524
rect 1915 11524 1987 11568
rect 1363 10244 1435 10288
rect 1915 10288 1928 11524
rect 1974 10288 1987 11524
rect 1915 10244 1987 10288
rect 2359 11568 2983 11640
rect 2359 11524 2431 11568
rect 2359 10288 2372 11524
rect 2418 10288 2431 11524
rect 2911 11524 2983 11568
rect 2359 10244 2431 10288
rect 2911 10288 2924 11524
rect 2970 10288 2983 11524
rect 2911 10244 2983 10288
rect 3355 11568 3979 11640
rect 3355 11524 3427 11568
rect 3355 10288 3368 11524
rect 3414 10288 3427 11524
rect 3907 11524 3979 11568
rect 3355 10244 3427 10288
rect 3907 10288 3920 11524
rect 3966 10288 3979 11524
rect 3907 10244 3979 10288
rect 4351 11568 4975 11640
rect 4351 11524 4423 11568
rect 4351 10288 4364 11524
rect 4410 10288 4423 11524
rect 4903 11524 4975 11568
rect 4351 10244 4423 10288
rect 4903 10288 4916 11524
rect 4962 10288 4975 11524
rect 4903 10244 4975 10288
rect 5347 11568 5971 11640
rect 5347 11524 5419 11568
rect 5347 10288 5360 11524
rect 5406 10288 5419 11524
rect 5899 11524 5971 11568
rect 5347 10244 5419 10288
rect 5899 10288 5912 11524
rect 5958 10288 5971 11524
rect 5899 10244 5971 10288
rect 6343 11568 6967 11640
rect 6343 11524 6415 11568
rect 6343 10288 6356 11524
rect 6402 10288 6415 11524
rect 6895 11524 6967 11568
rect 6343 10244 6415 10288
rect 6895 10288 6908 11524
rect 6954 10288 6967 11524
rect 6895 10244 6967 10288
rect 7339 11568 7963 11640
rect 7339 11524 7411 11568
rect 7339 10288 7352 11524
rect 7398 10288 7411 11524
rect 7891 11524 7963 11568
rect 7339 10244 7411 10288
rect 7891 10288 7904 11524
rect 7950 10288 7963 11524
rect 7891 10244 7963 10288
rect 8335 11568 8959 11640
rect 8335 11524 8407 11568
rect 8335 10288 8348 11524
rect 8394 10288 8407 11524
rect 8887 11524 8959 11568
rect 8335 10244 8407 10288
rect 8887 10288 8900 11524
rect 8946 10288 8959 11524
rect 8887 10244 8959 10288
rect 9331 11568 9955 11640
rect 9331 11524 9403 11568
rect 9331 10288 9344 11524
rect 9390 10288 9403 11524
rect 9883 11524 9955 11568
rect 9331 10244 9403 10288
rect 9883 10288 9896 11524
rect 9942 10288 9955 11524
rect 9883 10244 9955 10288
rect 10327 11568 10951 11640
rect 10327 11524 10399 11568
rect 10327 10288 10340 11524
rect 10386 10288 10399 11524
rect 10879 11524 10951 11568
rect 10327 10244 10399 10288
rect 10879 10288 10892 11524
rect 10938 10288 10951 11524
rect 10879 10244 10951 10288
rect 11323 11568 11947 11640
rect 11323 11524 11395 11568
rect 11323 10288 11336 11524
rect 11382 10288 11395 11524
rect 11875 11524 11947 11568
rect 11323 10244 11395 10288
rect 11875 10288 11888 11524
rect 11934 10288 11947 11524
rect 11875 10244 11947 10288
rect 367 10231 12791 10244
rect 367 10185 924 10231
rect 1319 10185 1920 10231
rect 2315 10185 2916 10231
rect 3311 10185 3912 10231
rect 4307 10185 4908 10231
rect 5303 10185 5904 10231
rect 6299 10185 6900 10231
rect 7295 10185 7896 10231
rect 8291 10185 8892 10231
rect 9287 10185 9888 10231
rect 10283 10185 10884 10231
rect 11279 10185 11439 10231
rect 12675 10185 12791 10231
rect 367 10172 12791 10185
rect 367 9692 439 10172
rect 1363 9692 1435 10172
rect 2359 9692 2431 10172
rect 3355 9692 3427 10172
rect 4351 9692 4423 10172
rect 5347 9692 5419 10172
rect 6343 9692 6415 10172
rect 7339 9692 7411 10172
rect 8335 9692 8407 10172
rect 9331 9692 9403 10172
rect 10327 9692 10399 10172
rect 11323 9692 11395 10172
rect 12719 9692 12791 10172
rect 367 9679 12791 9692
rect 367 9633 483 9679
rect 1319 9633 1479 9679
rect 2315 9633 2475 9679
rect 3311 9633 3471 9679
rect 4307 9633 4467 9679
rect 5303 9633 5463 9679
rect 6299 9633 6459 9679
rect 7295 9633 7455 9679
rect 8291 9633 8451 9679
rect 9287 9633 9447 9679
rect 10283 9633 10443 9679
rect 11279 9633 11439 9679
rect 12675 9633 12791 9679
rect 367 9620 12791 9633
rect 1055 9014 2231 9086
rect 1055 8970 1127 9014
rect 1055 8612 1068 8970
rect 367 8540 1068 8612
rect 367 8496 439 8540
rect 367 4060 380 8496
rect 426 4060 439 8496
rect 919 8496 1068 8540
rect 367 4016 439 4060
rect 919 4060 932 8496
rect 978 6534 1068 8496
rect 1114 6534 1127 8970
rect 1607 8970 1679 9014
rect 978 6490 1127 6534
rect 1607 6534 1620 8970
rect 1666 6534 1679 8970
rect 2159 8970 2231 9014
rect 1607 6490 1679 6534
rect 2159 6534 2172 8970
rect 2218 6534 2231 8970
rect 2159 6490 2231 6534
rect 978 6418 2231 6490
rect 978 5380 991 6418
rect 978 5308 1674 5380
rect 978 5264 1122 5308
rect 978 4060 1063 5264
rect 919 4016 1063 4060
rect 367 3944 1063 4016
rect 1050 148 1063 3944
rect 1109 148 1122 5264
rect 1602 2700 1674 5308
rect 1602 2628 2226 2700
rect 1602 2584 1674 2628
rect 1050 104 1122 148
rect 1602 148 1615 2584
rect 1661 148 1674 2584
rect 2154 2584 2226 2628
rect 1602 104 1674 148
rect 2154 148 2167 2584
rect 2213 148 2226 2584
rect 3621 4512 64533 4525
rect 3621 4466 3737 4512
rect 64417 4466 64533 4512
rect 3621 4453 64533 4466
rect 3621 2669 3693 4453
rect 64461 2669 64533 4453
rect 3621 2656 64533 2669
rect 3621 2610 3737 2656
rect 64417 2610 64533 2656
rect 3621 2598 64533 2610
rect 3548 2597 64533 2598
rect 3548 2496 3937 2597
rect 2154 104 2226 148
rect 1050 32 2226 104
rect 2453 2424 3937 2496
rect 2453 2380 2525 2424
rect 2453 164 2466 2380
rect 2512 164 2525 2380
rect 2965 2380 3037 2424
rect 2453 120 2525 164
rect 2965 164 2978 2380
rect 3024 164 3037 2380
rect 3477 2380 3937 2424
rect 2965 120 3037 164
rect 3477 164 3490 2380
rect 3536 2269 3937 2380
rect 3536 2256 64533 2269
rect 3536 2210 3737 2256
rect 64417 2210 64533 2256
rect 3536 2197 64533 2210
rect 3536 413 3693 2197
rect 64461 413 64533 2197
rect 3536 400 64533 413
rect 3536 354 3737 400
rect 64417 354 64533 400
rect 3536 341 64533 354
rect 3536 164 3549 341
rect 3477 120 3549 164
rect 2453 48 3549 120
<< mvnsubdiff >>
rect 2432 8991 3528 8992
rect 2432 8978 64536 8991
rect 2432 8932 3740 8978
rect 64420 8932 64536 8978
rect 2432 8920 64536 8932
rect 2432 8876 2504 8920
rect 2432 5860 2445 8876
rect 2491 5860 2504 8876
rect 2944 8876 3016 8920
rect 2432 5816 2504 5860
rect 2944 5860 2957 8876
rect 3003 5860 3016 8876
rect 3456 8919 64536 8920
rect 3456 8876 3696 8919
rect 2944 5816 3016 5860
rect 3456 5860 3469 8876
rect 3515 7135 3696 8876
rect 64464 7135 64536 8919
rect 3515 7122 64536 7135
rect 3515 7076 3740 7122
rect 64420 7076 64536 7122
rect 3515 7063 64536 7076
rect 3515 6735 3624 7063
rect 3515 6722 64536 6735
rect 3515 6676 3740 6722
rect 64420 6676 64536 6722
rect 3515 6663 64536 6676
rect 3515 5860 3696 6663
rect 3456 5816 3696 5860
rect 2298 5744 3696 5816
rect 2298 5700 2370 5744
rect 2298 2684 2311 5700
rect 2357 2684 2370 5700
rect 2810 5700 2882 5744
rect 2298 2640 2370 2684
rect 2810 2684 2823 5700
rect 2869 2684 2882 5700
rect 3322 5700 3394 5744
rect 2810 2640 2882 2684
rect 3322 2684 3335 5700
rect 3381 2684 3394 5700
rect 3624 4879 3696 5744
rect 64464 4879 64536 6663
rect 3624 4866 64536 4879
rect 3624 4820 3740 4866
rect 64420 4820 64536 4866
rect 3624 4807 64536 4820
rect 3322 2640 3394 2684
rect 2298 2568 3394 2640
<< mvpsubdiffcont >>
rect 380 10288 426 11524
rect 932 10288 978 11524
rect 1376 10288 1422 11524
rect 1928 10288 1974 11524
rect 2372 10288 2418 11524
rect 2924 10288 2970 11524
rect 3368 10288 3414 11524
rect 3920 10288 3966 11524
rect 4364 10288 4410 11524
rect 4916 10288 4962 11524
rect 5360 10288 5406 11524
rect 5912 10288 5958 11524
rect 6356 10288 6402 11524
rect 6908 10288 6954 11524
rect 7352 10288 7398 11524
rect 7904 10288 7950 11524
rect 8348 10288 8394 11524
rect 8900 10288 8946 11524
rect 9344 10288 9390 11524
rect 9896 10288 9942 11524
rect 10340 10288 10386 11524
rect 10892 10288 10938 11524
rect 11336 10288 11382 11524
rect 11888 10288 11934 11524
rect 924 10185 1319 10231
rect 1920 10185 2315 10231
rect 2916 10185 3311 10231
rect 3912 10185 4307 10231
rect 4908 10185 5303 10231
rect 5904 10185 6299 10231
rect 6900 10185 7295 10231
rect 7896 10185 8291 10231
rect 8892 10185 9287 10231
rect 9888 10185 10283 10231
rect 10884 10185 11279 10231
rect 11439 10185 12675 10231
rect 483 9633 1319 9679
rect 1479 9633 2315 9679
rect 2475 9633 3311 9679
rect 3471 9633 4307 9679
rect 4467 9633 5303 9679
rect 5463 9633 6299 9679
rect 6459 9633 7295 9679
rect 7455 9633 8291 9679
rect 8451 9633 9287 9679
rect 9447 9633 10283 9679
rect 10443 9633 11279 9679
rect 11439 9633 12675 9679
rect 380 4060 426 8496
rect 932 4060 978 8496
rect 1068 6534 1114 8970
rect 1620 6534 1666 8970
rect 2172 6534 2218 8970
rect 1063 148 1109 5264
rect 1615 148 1661 2584
rect 2167 148 2213 2584
rect 3737 4466 64417 4512
rect 3737 2610 64417 2656
rect 2466 164 2512 2380
rect 2978 164 3024 2380
rect 3490 164 3536 2380
rect 3737 2210 64417 2256
rect 3737 354 64417 400
<< mvnsubdiffcont >>
rect 3740 8932 64420 8978
rect 2445 5860 2491 8876
rect 2957 5860 3003 8876
rect 3469 5860 3515 8876
rect 3740 7076 64420 7122
rect 3740 6676 64420 6722
rect 2311 2684 2357 5700
rect 2823 2684 2869 5700
rect 3335 2684 3381 5700
rect 3740 4820 64420 4866
<< polysilicon >>
rect 579 11415 779 11428
rect 579 11369 592 11415
rect 766 11369 779 11415
rect 579 11306 779 11369
rect 579 10443 779 10506
rect 579 10397 592 10443
rect 766 10397 779 10443
rect 579 10384 779 10397
rect 1575 11415 1775 11428
rect 1575 11369 1588 11415
rect 1762 11369 1775 11415
rect 1575 11306 1775 11369
rect 1575 10443 1775 10506
rect 1575 10397 1588 10443
rect 1762 10397 1775 10443
rect 1575 10384 1775 10397
rect 2571 11415 2771 11428
rect 2571 11369 2584 11415
rect 2758 11369 2771 11415
rect 2571 11306 2771 11369
rect 2571 10443 2771 10506
rect 2571 10397 2584 10443
rect 2758 10397 2771 10443
rect 2571 10384 2771 10397
rect 3567 11415 3767 11428
rect 3567 11369 3580 11415
rect 3754 11369 3767 11415
rect 3567 11306 3767 11369
rect 3567 10443 3767 10506
rect 3567 10397 3580 10443
rect 3754 10397 3767 10443
rect 3567 10384 3767 10397
rect 4563 11415 4763 11428
rect 4563 11369 4576 11415
rect 4750 11369 4763 11415
rect 4563 11306 4763 11369
rect 4563 10443 4763 10506
rect 4563 10397 4576 10443
rect 4750 10397 4763 10443
rect 4563 10384 4763 10397
rect 5559 11415 5759 11428
rect 5559 11369 5572 11415
rect 5746 11369 5759 11415
rect 5559 11306 5759 11369
rect 5559 10443 5759 10506
rect 5559 10397 5572 10443
rect 5746 10397 5759 10443
rect 5559 10384 5759 10397
rect 6555 11415 6755 11428
rect 6555 11369 6568 11415
rect 6742 11369 6755 11415
rect 6555 11306 6755 11369
rect 6555 10443 6755 10506
rect 6555 10397 6568 10443
rect 6742 10397 6755 10443
rect 6555 10384 6755 10397
rect 7551 11415 7751 11428
rect 7551 11369 7564 11415
rect 7738 11369 7751 11415
rect 7551 11306 7751 11369
rect 7551 10443 7751 10506
rect 7551 10397 7564 10443
rect 7738 10397 7751 10443
rect 7551 10384 7751 10397
rect 8547 11415 8747 11428
rect 8547 11369 8560 11415
rect 8734 11369 8747 11415
rect 8547 11306 8747 11369
rect 8547 10443 8747 10506
rect 8547 10397 8560 10443
rect 8734 10397 8747 10443
rect 8547 10384 8747 10397
rect 9543 11415 9743 11428
rect 9543 11369 9556 11415
rect 9730 11369 9743 11415
rect 9543 11306 9743 11369
rect 9543 10443 9743 10506
rect 9543 10397 9556 10443
rect 9730 10397 9743 10443
rect 9543 10384 9743 10397
rect 10539 11415 10739 11428
rect 10539 11369 10552 11415
rect 10726 11369 10739 11415
rect 10539 11306 10739 11369
rect 10539 10443 10739 10506
rect 10539 10397 10552 10443
rect 10726 10397 10739 10443
rect 10539 10384 10739 10397
rect 11535 11415 11735 11428
rect 11535 11369 11548 11415
rect 11722 11369 11735 11415
rect 11535 11306 11735 11369
rect 11535 10443 11735 10506
rect 11535 10397 11548 10443
rect 11722 10397 11735 10443
rect 11535 10384 11735 10397
rect 579 10019 701 10032
rect 579 9845 592 10019
rect 638 9845 701 10019
rect 579 9832 701 9845
rect 1101 10019 1223 10032
rect 1101 9845 1164 10019
rect 1210 9845 1223 10019
rect 1101 9832 1223 9845
rect 1575 10019 1697 10032
rect 1575 9845 1588 10019
rect 1634 9845 1697 10019
rect 1575 9832 1697 9845
rect 2097 10019 2219 10032
rect 2097 9845 2160 10019
rect 2206 9845 2219 10019
rect 2097 9832 2219 9845
rect 2571 10019 2693 10032
rect 2571 9845 2584 10019
rect 2630 9845 2693 10019
rect 2571 9832 2693 9845
rect 3093 10019 3215 10032
rect 3093 9845 3156 10019
rect 3202 9845 3215 10019
rect 3093 9832 3215 9845
rect 3567 10019 3689 10032
rect 3567 9845 3580 10019
rect 3626 9845 3689 10019
rect 3567 9832 3689 9845
rect 4089 10019 4211 10032
rect 4089 9845 4152 10019
rect 4198 9845 4211 10019
rect 4089 9832 4211 9845
rect 4563 10019 4685 10032
rect 4563 9845 4576 10019
rect 4622 9845 4685 10019
rect 4563 9832 4685 9845
rect 5085 10019 5207 10032
rect 5085 9845 5148 10019
rect 5194 9845 5207 10019
rect 5085 9832 5207 9845
rect 5559 10019 5681 10032
rect 5559 9845 5572 10019
rect 5618 9845 5681 10019
rect 5559 9832 5681 9845
rect 6081 10019 6203 10032
rect 6081 9845 6144 10019
rect 6190 9845 6203 10019
rect 6081 9832 6203 9845
rect 6555 10019 6677 10032
rect 6555 9845 6568 10019
rect 6614 9845 6677 10019
rect 6555 9832 6677 9845
rect 7077 10019 7199 10032
rect 7077 9845 7140 10019
rect 7186 9845 7199 10019
rect 7077 9832 7199 9845
rect 7551 10019 7673 10032
rect 7551 9845 7564 10019
rect 7610 9845 7673 10019
rect 7551 9832 7673 9845
rect 8073 10019 8195 10032
rect 8073 9845 8136 10019
rect 8182 9845 8195 10019
rect 8073 9832 8195 9845
rect 8547 10019 8669 10032
rect 8547 9845 8560 10019
rect 8606 9845 8669 10019
rect 8547 9832 8669 9845
rect 9069 10019 9191 10032
rect 9069 9845 9132 10019
rect 9178 9845 9191 10019
rect 9069 9832 9191 9845
rect 9543 10019 9665 10032
rect 9543 9845 9556 10019
rect 9602 9845 9665 10019
rect 9543 9832 9665 9845
rect 10065 10019 10187 10032
rect 10065 9845 10128 10019
rect 10174 9845 10187 10019
rect 10065 9832 10187 9845
rect 10539 10019 10661 10032
rect 10539 9845 10552 10019
rect 10598 9845 10661 10019
rect 10539 9832 10661 9845
rect 11061 10019 11183 10032
rect 11061 9845 11124 10019
rect 11170 9845 11183 10019
rect 11061 9832 11183 9845
rect 11535 10019 11657 10032
rect 11535 9845 11548 10019
rect 11594 9845 11657 10019
rect 11535 9832 11657 9845
rect 12457 10019 12579 10032
rect 12457 9845 12520 10019
rect 12566 9845 12579 10019
rect 12457 9832 12579 9845
rect 579 8387 779 8400
rect 579 8341 592 8387
rect 766 8341 779 8387
rect 579 8278 779 8341
rect 579 4215 779 4278
rect 579 4169 592 4215
rect 766 4169 779 4215
rect 579 4156 779 4169
rect 1267 8861 1467 8874
rect 1267 8815 1280 8861
rect 1454 8815 1467 8861
rect 1267 8752 1467 8815
rect 1267 6689 1467 6752
rect 1267 6643 1280 6689
rect 1454 6643 1467 6689
rect 1267 6630 1467 6643
rect 1819 8861 2019 8874
rect 1819 8815 1832 8861
rect 2006 8815 2019 8861
rect 1819 8752 2019 8815
rect 1819 6689 2019 6752
rect 1819 6643 1832 6689
rect 2006 6643 2019 6689
rect 1819 6630 2019 6643
rect 2664 8847 2784 8860
rect 2664 8801 2677 8847
rect 2771 8801 2784 8847
rect 2664 8768 2784 8801
rect 2664 5935 2784 5968
rect 2664 5889 2677 5935
rect 2771 5889 2784 5935
rect 2664 5876 2784 5889
rect 3176 8847 3296 8860
rect 3176 8801 3189 8847
rect 3283 8801 3296 8847
rect 3176 8768 3296 8801
rect 3176 5935 3296 5968
rect 3176 5889 3189 5935
rect 3283 5889 3296 5935
rect 3176 5876 3296 5889
rect 3756 8746 3848 8759
rect 3756 8652 3769 8746
rect 3815 8652 3848 8746
rect 3756 8639 3848 8652
rect 23848 8742 24080 8759
rect 23848 8656 23881 8742
rect 23927 8656 24001 8742
rect 24047 8656 24080 8742
rect 23848 8639 24080 8656
rect 44080 8742 44312 8759
rect 44080 8656 44113 8742
rect 44159 8656 44233 8742
rect 44279 8656 44312 8742
rect 44080 8639 44312 8656
rect 64312 8746 64404 8759
rect 64312 8652 64345 8746
rect 64391 8652 64404 8746
rect 64312 8639 64404 8652
rect 3756 8522 3848 8535
rect 3756 8428 3769 8522
rect 3815 8428 3848 8522
rect 3756 8415 3848 8428
rect 23848 8518 24080 8535
rect 23848 8432 23881 8518
rect 23927 8432 24001 8518
rect 24047 8432 24080 8518
rect 23848 8415 24080 8432
rect 44080 8518 44312 8535
rect 44080 8432 44113 8518
rect 44159 8432 44233 8518
rect 44279 8432 44312 8518
rect 44080 8415 44312 8432
rect 64312 8522 64404 8535
rect 64312 8428 64345 8522
rect 64391 8428 64404 8522
rect 64312 8415 64404 8428
rect 3756 8298 3848 8311
rect 3756 8204 3769 8298
rect 3815 8204 3848 8298
rect 3756 8191 3848 8204
rect 23848 8294 24080 8311
rect 23848 8208 23881 8294
rect 23927 8208 24001 8294
rect 24047 8208 24080 8294
rect 23848 8191 24080 8208
rect 44080 8294 44312 8311
rect 44080 8208 44113 8294
rect 44159 8208 44233 8294
rect 44279 8208 44312 8294
rect 44080 8191 44312 8208
rect 64312 8298 64404 8311
rect 64312 8204 64345 8298
rect 64391 8204 64404 8298
rect 64312 8191 64404 8204
rect 3756 8074 3848 8087
rect 3756 7980 3769 8074
rect 3815 7980 3848 8074
rect 3756 7967 3848 7980
rect 23848 8070 24080 8087
rect 23848 7984 23881 8070
rect 23927 7984 24001 8070
rect 24047 7984 24080 8070
rect 23848 7967 24080 7984
rect 44080 8070 44312 8087
rect 44080 7984 44113 8070
rect 44159 7984 44233 8070
rect 44279 7984 44312 8070
rect 44080 7967 44312 7984
rect 64312 8074 64404 8087
rect 64312 7980 64345 8074
rect 64391 7980 64404 8074
rect 64312 7967 64404 7980
rect 3756 7850 3848 7863
rect 3756 7756 3769 7850
rect 3815 7756 3848 7850
rect 3756 7743 3848 7756
rect 23848 7846 24080 7863
rect 23848 7760 23881 7846
rect 23927 7760 24001 7846
rect 24047 7760 24080 7846
rect 23848 7743 24080 7760
rect 44080 7846 44312 7863
rect 44080 7760 44113 7846
rect 44159 7760 44233 7846
rect 44279 7760 44312 7846
rect 44080 7743 44312 7760
rect 64312 7850 64404 7863
rect 64312 7756 64345 7850
rect 64391 7756 64404 7850
rect 64312 7743 64404 7756
rect 3756 7626 3848 7639
rect 3756 7532 3769 7626
rect 3815 7532 3848 7626
rect 3756 7519 3848 7532
rect 23848 7622 24080 7639
rect 23848 7536 23881 7622
rect 23927 7536 24001 7622
rect 24047 7536 24080 7622
rect 23848 7519 24080 7536
rect 44080 7622 44312 7639
rect 44080 7536 44113 7622
rect 44159 7536 44233 7622
rect 44279 7536 44312 7622
rect 44080 7519 44312 7536
rect 64312 7626 64404 7639
rect 64312 7532 64345 7626
rect 64391 7532 64404 7626
rect 64312 7519 64404 7532
rect 3756 7402 3848 7415
rect 3756 7308 3769 7402
rect 3815 7308 3848 7402
rect 3756 7295 3848 7308
rect 23848 7398 24080 7415
rect 23848 7312 23881 7398
rect 23927 7312 24001 7398
rect 24047 7312 24080 7398
rect 23848 7295 24080 7312
rect 44080 7398 44312 7415
rect 44080 7312 44113 7398
rect 44159 7312 44233 7398
rect 44279 7312 44312 7398
rect 44080 7295 44312 7312
rect 64312 7402 64404 7415
rect 64312 7308 64345 7402
rect 64391 7308 64404 7402
rect 64312 7295 64404 7308
rect 3756 6490 3848 6503
rect 3756 6396 3769 6490
rect 3815 6396 3848 6490
rect 3756 6383 3848 6396
rect 23848 6486 24080 6503
rect 23848 6400 23881 6486
rect 23927 6400 24001 6486
rect 24047 6400 24080 6486
rect 23848 6383 24080 6400
rect 44080 6486 44312 6503
rect 44080 6400 44113 6486
rect 44159 6400 44233 6486
rect 44279 6400 44312 6486
rect 44080 6383 44312 6400
rect 64312 6490 64404 6503
rect 64312 6396 64345 6490
rect 64391 6396 64404 6490
rect 64312 6383 64404 6396
rect 3756 6266 3848 6279
rect 3756 6172 3769 6266
rect 3815 6172 3848 6266
rect 3756 6159 3848 6172
rect 23848 6262 24080 6279
rect 23848 6176 23881 6262
rect 23927 6176 24001 6262
rect 24047 6176 24080 6262
rect 23848 6159 24080 6176
rect 44080 6262 44312 6279
rect 44080 6176 44113 6262
rect 44159 6176 44233 6262
rect 44279 6176 44312 6262
rect 44080 6159 44312 6176
rect 64312 6266 64404 6279
rect 64312 6172 64345 6266
rect 64391 6172 64404 6266
rect 64312 6159 64404 6172
rect 3756 6042 3848 6055
rect 3756 5948 3769 6042
rect 3815 5948 3848 6042
rect 3756 5935 3848 5948
rect 23848 6038 24080 6055
rect 23848 5952 23881 6038
rect 23927 5952 24001 6038
rect 24047 5952 24080 6038
rect 23848 5935 24080 5952
rect 44080 6038 44312 6055
rect 44080 5952 44113 6038
rect 44159 5952 44233 6038
rect 44279 5952 44312 6038
rect 44080 5935 44312 5952
rect 64312 6042 64404 6055
rect 64312 5948 64345 6042
rect 64391 5948 64404 6042
rect 64312 5935 64404 5948
rect 1262 5155 1462 5168
rect 1262 5109 1275 5155
rect 1449 5109 1462 5155
rect 1262 5046 1462 5109
rect 1262 303 1462 366
rect 1262 257 1275 303
rect 1449 257 1462 303
rect 1262 244 1462 257
rect 1814 2475 2014 2488
rect 1814 2429 1827 2475
rect 2001 2429 2014 2475
rect 1814 2366 2014 2429
rect 1814 303 2014 366
rect 1814 257 1827 303
rect 2001 257 2014 303
rect 1814 244 2014 257
rect 2530 5671 2650 5684
rect 2530 5625 2543 5671
rect 2637 5625 2650 5671
rect 2530 5592 2650 5625
rect 2530 2759 2650 2792
rect 2530 2713 2543 2759
rect 2637 2713 2650 2759
rect 2530 2700 2650 2713
rect 3042 5671 3162 5684
rect 3042 5625 3055 5671
rect 3149 5625 3162 5671
rect 3042 5592 3162 5625
rect 3042 2759 3162 2792
rect 3042 2713 3055 2759
rect 3149 2713 3162 2759
rect 3042 2700 3162 2713
rect 3756 5818 3848 5831
rect 3756 5724 3769 5818
rect 3815 5724 3848 5818
rect 3756 5711 3848 5724
rect 23848 5814 24080 5831
rect 23848 5728 23881 5814
rect 23927 5728 24001 5814
rect 24047 5728 24080 5814
rect 23848 5711 24080 5728
rect 44080 5814 44312 5831
rect 44080 5728 44113 5814
rect 44159 5728 44233 5814
rect 44279 5728 44312 5814
rect 44080 5711 44312 5728
rect 64312 5818 64404 5831
rect 64312 5724 64345 5818
rect 64391 5724 64404 5818
rect 64312 5711 64404 5724
rect 3756 5594 3848 5607
rect 3756 5500 3769 5594
rect 3815 5500 3848 5594
rect 3756 5487 3848 5500
rect 23848 5590 24080 5607
rect 23848 5504 23881 5590
rect 23927 5504 24001 5590
rect 24047 5504 24080 5590
rect 23848 5487 24080 5504
rect 44080 5590 44312 5607
rect 44080 5504 44113 5590
rect 44159 5504 44233 5590
rect 44279 5504 44312 5590
rect 44080 5487 44312 5504
rect 64312 5594 64404 5607
rect 64312 5500 64345 5594
rect 64391 5500 64404 5594
rect 64312 5487 64404 5500
rect 3756 5370 3848 5383
rect 3756 5276 3769 5370
rect 3815 5276 3848 5370
rect 3756 5263 3848 5276
rect 23848 5366 24080 5383
rect 23848 5280 23881 5366
rect 23927 5280 24001 5366
rect 24047 5280 24080 5366
rect 23848 5263 24080 5280
rect 44080 5366 44312 5383
rect 44080 5280 44113 5366
rect 44159 5280 44233 5366
rect 44279 5280 44312 5366
rect 44080 5263 44312 5280
rect 64312 5370 64404 5383
rect 64312 5276 64345 5370
rect 64391 5276 64404 5370
rect 64312 5263 64404 5276
rect 3756 5146 3848 5159
rect 3756 5052 3769 5146
rect 3815 5052 3848 5146
rect 3756 5039 3848 5052
rect 23848 5142 24080 5159
rect 23848 5056 23881 5142
rect 23927 5056 24001 5142
rect 24047 5056 24080 5142
rect 23848 5039 24080 5056
rect 44080 5142 44312 5159
rect 44080 5056 44113 5142
rect 44159 5056 44233 5142
rect 44279 5056 44312 5142
rect 44080 5039 44312 5056
rect 64312 5146 64404 5159
rect 64312 5052 64345 5146
rect 64391 5052 64404 5146
rect 64312 5039 64404 5052
rect 3753 4280 3845 4293
rect 3753 4186 3766 4280
rect 3812 4186 3845 4280
rect 3753 4173 3845 4186
rect 23845 4276 24077 4293
rect 23845 4190 23878 4276
rect 23924 4190 23998 4276
rect 24044 4190 24077 4276
rect 23845 4173 24077 4190
rect 44077 4276 44309 4293
rect 44077 4190 44110 4276
rect 44156 4190 44230 4276
rect 44276 4190 44309 4276
rect 44077 4173 44309 4190
rect 64309 4280 64401 4293
rect 64309 4186 64342 4280
rect 64388 4186 64401 4280
rect 64309 4173 64401 4186
rect 3753 4056 3845 4069
rect 3753 3962 3766 4056
rect 3812 3962 3845 4056
rect 3753 3949 3845 3962
rect 23845 4052 24077 4069
rect 23845 3966 23878 4052
rect 23924 3966 23998 4052
rect 24044 3966 24077 4052
rect 23845 3949 24077 3966
rect 44077 4052 44309 4069
rect 44077 3966 44110 4052
rect 44156 3966 44230 4052
rect 44276 3966 44309 4052
rect 44077 3949 44309 3966
rect 64309 4056 64401 4069
rect 64309 3962 64342 4056
rect 64388 3962 64401 4056
rect 64309 3949 64401 3962
rect 3753 3832 3845 3845
rect 3753 3738 3766 3832
rect 3812 3738 3845 3832
rect 3753 3725 3845 3738
rect 23845 3828 24077 3845
rect 23845 3742 23878 3828
rect 23924 3742 23998 3828
rect 24044 3742 24077 3828
rect 23845 3725 24077 3742
rect 44077 3828 44309 3845
rect 44077 3742 44110 3828
rect 44156 3742 44230 3828
rect 44276 3742 44309 3828
rect 44077 3725 44309 3742
rect 64309 3832 64401 3845
rect 64309 3738 64342 3832
rect 64388 3738 64401 3832
rect 64309 3725 64401 3738
rect 3753 3608 3845 3621
rect 3753 3514 3766 3608
rect 3812 3514 3845 3608
rect 3753 3501 3845 3514
rect 23845 3604 24077 3621
rect 23845 3518 23878 3604
rect 23924 3518 23998 3604
rect 24044 3518 24077 3604
rect 23845 3501 24077 3518
rect 44077 3604 44309 3621
rect 44077 3518 44110 3604
rect 44156 3518 44230 3604
rect 44276 3518 44309 3604
rect 44077 3501 44309 3518
rect 64309 3608 64401 3621
rect 64309 3514 64342 3608
rect 64388 3514 64401 3608
rect 64309 3501 64401 3514
rect 3753 3384 3845 3397
rect 3753 3290 3766 3384
rect 3812 3290 3845 3384
rect 3753 3277 3845 3290
rect 23845 3380 24077 3397
rect 23845 3294 23878 3380
rect 23924 3294 23998 3380
rect 24044 3294 24077 3380
rect 23845 3277 24077 3294
rect 44077 3380 44309 3397
rect 44077 3294 44110 3380
rect 44156 3294 44230 3380
rect 44276 3294 44309 3380
rect 44077 3277 44309 3294
rect 64309 3384 64401 3397
rect 64309 3290 64342 3384
rect 64388 3290 64401 3384
rect 64309 3277 64401 3290
rect 3753 3160 3845 3173
rect 3753 3066 3766 3160
rect 3812 3066 3845 3160
rect 3753 3053 3845 3066
rect 23845 3156 24077 3173
rect 23845 3070 23878 3156
rect 23924 3070 23998 3156
rect 24044 3070 24077 3156
rect 23845 3053 24077 3070
rect 44077 3156 44309 3173
rect 44077 3070 44110 3156
rect 44156 3070 44230 3156
rect 44276 3070 44309 3156
rect 44077 3053 44309 3070
rect 64309 3160 64401 3173
rect 64309 3066 64342 3160
rect 64388 3066 64401 3160
rect 64309 3053 64401 3066
rect 3753 2936 3845 2949
rect 3753 2842 3766 2936
rect 3812 2842 3845 2936
rect 3753 2829 3845 2842
rect 23845 2932 24077 2949
rect 23845 2846 23878 2932
rect 23924 2846 23998 2932
rect 24044 2846 24077 2932
rect 23845 2829 24077 2846
rect 44077 2932 44309 2949
rect 44077 2846 44110 2932
rect 44156 2846 44230 2932
rect 44276 2846 44309 2932
rect 44077 2829 44309 2846
rect 64309 2936 64401 2949
rect 64309 2842 64342 2936
rect 64388 2842 64401 2936
rect 64309 2829 64401 2842
rect 2685 2351 2805 2364
rect 2685 2305 2698 2351
rect 2792 2305 2805 2351
rect 2685 2272 2805 2305
rect 2685 239 2805 272
rect 2685 193 2698 239
rect 2792 193 2805 239
rect 2685 180 2805 193
rect 3197 2351 3317 2364
rect 3197 2305 3210 2351
rect 3304 2305 3317 2351
rect 3197 2272 3317 2305
rect 3197 239 3317 272
rect 3197 193 3210 239
rect 3304 193 3317 239
rect 3197 180 3317 193
rect 3753 2024 3845 2037
rect 3753 1930 3766 2024
rect 3812 1930 3845 2024
rect 3753 1917 3845 1930
rect 23845 2020 24077 2037
rect 23845 1934 23878 2020
rect 23924 1934 23998 2020
rect 24044 1934 24077 2020
rect 23845 1917 24077 1934
rect 44077 2020 44309 2037
rect 44077 1934 44110 2020
rect 44156 1934 44230 2020
rect 44276 1934 44309 2020
rect 44077 1917 44309 1934
rect 64309 2024 64401 2037
rect 64309 1930 64342 2024
rect 64388 1930 64401 2024
rect 64309 1917 64401 1930
rect 3753 1800 3845 1813
rect 3753 1706 3766 1800
rect 3812 1706 3845 1800
rect 3753 1693 3845 1706
rect 23845 1796 24077 1813
rect 23845 1710 23878 1796
rect 23924 1710 23998 1796
rect 24044 1710 24077 1796
rect 23845 1693 24077 1710
rect 44077 1796 44309 1813
rect 44077 1710 44110 1796
rect 44156 1710 44230 1796
rect 44276 1710 44309 1796
rect 44077 1693 44309 1710
rect 64309 1800 64401 1813
rect 64309 1706 64342 1800
rect 64388 1706 64401 1800
rect 64309 1693 64401 1706
rect 3753 1576 3845 1589
rect 3753 1482 3766 1576
rect 3812 1482 3845 1576
rect 3753 1469 3845 1482
rect 23845 1572 24077 1589
rect 23845 1486 23878 1572
rect 23924 1486 23998 1572
rect 24044 1486 24077 1572
rect 23845 1469 24077 1486
rect 44077 1572 44309 1589
rect 44077 1486 44110 1572
rect 44156 1486 44230 1572
rect 44276 1486 44309 1572
rect 44077 1469 44309 1486
rect 64309 1576 64401 1589
rect 64309 1482 64342 1576
rect 64388 1482 64401 1576
rect 64309 1469 64401 1482
rect 3753 1352 3845 1365
rect 3753 1258 3766 1352
rect 3812 1258 3845 1352
rect 3753 1245 3845 1258
rect 23845 1348 24077 1365
rect 23845 1262 23878 1348
rect 23924 1262 23998 1348
rect 24044 1262 24077 1348
rect 23845 1245 24077 1262
rect 44077 1348 44309 1365
rect 44077 1262 44110 1348
rect 44156 1262 44230 1348
rect 44276 1262 44309 1348
rect 44077 1245 44309 1262
rect 64309 1352 64401 1365
rect 64309 1258 64342 1352
rect 64388 1258 64401 1352
rect 64309 1245 64401 1258
rect 3753 1128 3845 1141
rect 3753 1034 3766 1128
rect 3812 1034 3845 1128
rect 3753 1021 3845 1034
rect 23845 1124 24077 1141
rect 23845 1038 23878 1124
rect 23924 1038 23998 1124
rect 24044 1038 24077 1124
rect 23845 1021 24077 1038
rect 44077 1124 44309 1141
rect 44077 1038 44110 1124
rect 44156 1038 44230 1124
rect 44276 1038 44309 1124
rect 44077 1021 44309 1038
rect 64309 1128 64401 1141
rect 64309 1034 64342 1128
rect 64388 1034 64401 1128
rect 64309 1021 64401 1034
rect 3753 904 3845 917
rect 3753 810 3766 904
rect 3812 810 3845 904
rect 3753 797 3845 810
rect 23845 900 24077 917
rect 23845 814 23878 900
rect 23924 814 23998 900
rect 24044 814 24077 900
rect 23845 797 24077 814
rect 44077 900 44309 917
rect 44077 814 44110 900
rect 44156 814 44230 900
rect 44276 814 44309 900
rect 44077 797 44309 814
rect 64309 904 64401 917
rect 64309 810 64342 904
rect 64388 810 64401 904
rect 64309 797 64401 810
rect 3753 680 3845 693
rect 3753 586 3766 680
rect 3812 586 3845 680
rect 3753 573 3845 586
rect 23845 676 24077 693
rect 23845 590 23878 676
rect 23924 590 23998 676
rect 24044 590 24077 676
rect 23845 573 24077 590
rect 44077 676 44309 693
rect 44077 590 44110 676
rect 44156 590 44230 676
rect 44276 590 44309 676
rect 44077 573 44309 590
rect 64309 680 64401 693
rect 64309 586 64342 680
rect 64388 586 64401 680
rect 64309 573 64401 586
<< polycontact >>
rect 592 11369 766 11415
rect 592 10397 766 10443
rect 1588 11369 1762 11415
rect 1588 10397 1762 10443
rect 2584 11369 2758 11415
rect 2584 10397 2758 10443
rect 3580 11369 3754 11415
rect 3580 10397 3754 10443
rect 4576 11369 4750 11415
rect 4576 10397 4750 10443
rect 5572 11369 5746 11415
rect 5572 10397 5746 10443
rect 6568 11369 6742 11415
rect 6568 10397 6742 10443
rect 7564 11369 7738 11415
rect 7564 10397 7738 10443
rect 8560 11369 8734 11415
rect 8560 10397 8734 10443
rect 9556 11369 9730 11415
rect 9556 10397 9730 10443
rect 10552 11369 10726 11415
rect 10552 10397 10726 10443
rect 11548 11369 11722 11415
rect 11548 10397 11722 10443
rect 592 9845 638 10019
rect 1164 9845 1210 10019
rect 1588 9845 1634 10019
rect 2160 9845 2206 10019
rect 2584 9845 2630 10019
rect 3156 9845 3202 10019
rect 3580 9845 3626 10019
rect 4152 9845 4198 10019
rect 4576 9845 4622 10019
rect 5148 9845 5194 10019
rect 5572 9845 5618 10019
rect 6144 9845 6190 10019
rect 6568 9845 6614 10019
rect 7140 9845 7186 10019
rect 7564 9845 7610 10019
rect 8136 9845 8182 10019
rect 8560 9845 8606 10019
rect 9132 9845 9178 10019
rect 9556 9845 9602 10019
rect 10128 9845 10174 10019
rect 10552 9845 10598 10019
rect 11124 9845 11170 10019
rect 11548 9845 11594 10019
rect 12520 9845 12566 10019
rect 592 8341 766 8387
rect 592 4169 766 4215
rect 1280 8815 1454 8861
rect 1280 6643 1454 6689
rect 1832 8815 2006 8861
rect 1832 6643 2006 6689
rect 2677 8801 2771 8847
rect 2677 5889 2771 5935
rect 3189 8801 3283 8847
rect 3189 5889 3283 5935
rect 3769 8652 3815 8746
rect 23881 8656 23927 8742
rect 24001 8656 24047 8742
rect 44113 8656 44159 8742
rect 44233 8656 44279 8742
rect 64345 8652 64391 8746
rect 3769 8428 3815 8522
rect 23881 8432 23927 8518
rect 24001 8432 24047 8518
rect 44113 8432 44159 8518
rect 44233 8432 44279 8518
rect 64345 8428 64391 8522
rect 3769 8204 3815 8298
rect 23881 8208 23927 8294
rect 24001 8208 24047 8294
rect 44113 8208 44159 8294
rect 44233 8208 44279 8294
rect 64345 8204 64391 8298
rect 3769 7980 3815 8074
rect 23881 7984 23927 8070
rect 24001 7984 24047 8070
rect 44113 7984 44159 8070
rect 44233 7984 44279 8070
rect 64345 7980 64391 8074
rect 3769 7756 3815 7850
rect 23881 7760 23927 7846
rect 24001 7760 24047 7846
rect 44113 7760 44159 7846
rect 44233 7760 44279 7846
rect 64345 7756 64391 7850
rect 3769 7532 3815 7626
rect 23881 7536 23927 7622
rect 24001 7536 24047 7622
rect 44113 7536 44159 7622
rect 44233 7536 44279 7622
rect 64345 7532 64391 7626
rect 3769 7308 3815 7402
rect 23881 7312 23927 7398
rect 24001 7312 24047 7398
rect 44113 7312 44159 7398
rect 44233 7312 44279 7398
rect 64345 7308 64391 7402
rect 3769 6396 3815 6490
rect 23881 6400 23927 6486
rect 24001 6400 24047 6486
rect 44113 6400 44159 6486
rect 44233 6400 44279 6486
rect 64345 6396 64391 6490
rect 3769 6172 3815 6266
rect 23881 6176 23927 6262
rect 24001 6176 24047 6262
rect 44113 6176 44159 6262
rect 44233 6176 44279 6262
rect 64345 6172 64391 6266
rect 3769 5948 3815 6042
rect 23881 5952 23927 6038
rect 24001 5952 24047 6038
rect 44113 5952 44159 6038
rect 44233 5952 44279 6038
rect 64345 5948 64391 6042
rect 1275 5109 1449 5155
rect 1275 257 1449 303
rect 1827 2429 2001 2475
rect 1827 257 2001 303
rect 2543 5625 2637 5671
rect 2543 2713 2637 2759
rect 3055 5625 3149 5671
rect 3055 2713 3149 2759
rect 3769 5724 3815 5818
rect 23881 5728 23927 5814
rect 24001 5728 24047 5814
rect 44113 5728 44159 5814
rect 44233 5728 44279 5814
rect 64345 5724 64391 5818
rect 3769 5500 3815 5594
rect 23881 5504 23927 5590
rect 24001 5504 24047 5590
rect 44113 5504 44159 5590
rect 44233 5504 44279 5590
rect 64345 5500 64391 5594
rect 3769 5276 3815 5370
rect 23881 5280 23927 5366
rect 24001 5280 24047 5366
rect 44113 5280 44159 5366
rect 44233 5280 44279 5366
rect 64345 5276 64391 5370
rect 3769 5052 3815 5146
rect 23881 5056 23927 5142
rect 24001 5056 24047 5142
rect 44113 5056 44159 5142
rect 44233 5056 44279 5142
rect 64345 5052 64391 5146
rect 3766 4186 3812 4280
rect 23878 4190 23924 4276
rect 23998 4190 24044 4276
rect 44110 4190 44156 4276
rect 44230 4190 44276 4276
rect 64342 4186 64388 4280
rect 3766 3962 3812 4056
rect 23878 3966 23924 4052
rect 23998 3966 24044 4052
rect 44110 3966 44156 4052
rect 44230 3966 44276 4052
rect 64342 3962 64388 4056
rect 3766 3738 3812 3832
rect 23878 3742 23924 3828
rect 23998 3742 24044 3828
rect 44110 3742 44156 3828
rect 44230 3742 44276 3828
rect 64342 3738 64388 3832
rect 3766 3514 3812 3608
rect 23878 3518 23924 3604
rect 23998 3518 24044 3604
rect 44110 3518 44156 3604
rect 44230 3518 44276 3604
rect 64342 3514 64388 3608
rect 3766 3290 3812 3384
rect 23878 3294 23924 3380
rect 23998 3294 24044 3380
rect 44110 3294 44156 3380
rect 44230 3294 44276 3380
rect 64342 3290 64388 3384
rect 3766 3066 3812 3160
rect 23878 3070 23924 3156
rect 23998 3070 24044 3156
rect 44110 3070 44156 3156
rect 44230 3070 44276 3156
rect 64342 3066 64388 3160
rect 3766 2842 3812 2936
rect 23878 2846 23924 2932
rect 23998 2846 24044 2932
rect 44110 2846 44156 2932
rect 44230 2846 44276 2932
rect 64342 2842 64388 2936
rect 2698 2305 2792 2351
rect 2698 193 2792 239
rect 3210 2305 3304 2351
rect 3210 193 3304 239
rect 3766 1930 3812 2024
rect 23878 1934 23924 2020
rect 23998 1934 24044 2020
rect 44110 1934 44156 2020
rect 44230 1934 44276 2020
rect 64342 1930 64388 2024
rect 3766 1706 3812 1800
rect 23878 1710 23924 1796
rect 23998 1710 24044 1796
rect 44110 1710 44156 1796
rect 44230 1710 44276 1796
rect 64342 1706 64388 1800
rect 3766 1482 3812 1576
rect 23878 1486 23924 1572
rect 23998 1486 24044 1572
rect 44110 1486 44156 1572
rect 44230 1486 44276 1572
rect 64342 1482 64388 1576
rect 3766 1258 3812 1352
rect 23878 1262 23924 1348
rect 23998 1262 24044 1348
rect 44110 1262 44156 1348
rect 44230 1262 44276 1348
rect 64342 1258 64388 1352
rect 3766 1034 3812 1128
rect 23878 1038 23924 1124
rect 23998 1038 24044 1124
rect 44110 1038 44156 1124
rect 44230 1038 44276 1124
rect 64342 1034 64388 1128
rect 3766 810 3812 904
rect 23878 814 23924 900
rect 23998 814 24044 900
rect 44110 814 44156 900
rect 44230 814 44276 900
rect 64342 810 64388 904
rect 3766 586 3812 680
rect 23878 590 23924 676
rect 23998 590 24044 676
rect 44110 590 44156 676
rect 44230 590 44276 676
rect 64342 586 64388 680
<< mvnhighres >>
rect 579 10506 779 11306
rect 1575 10506 1775 11306
rect 2571 10506 2771 11306
rect 3567 10506 3767 11306
rect 4563 10506 4763 11306
rect 5559 10506 5759 11306
rect 6555 10506 6755 11306
rect 7551 10506 7751 11306
rect 8547 10506 8747 11306
rect 9543 10506 9743 11306
rect 10539 10506 10739 11306
rect 11535 10506 11735 11306
rect 701 9832 1101 10032
rect 1697 9832 2097 10032
rect 2693 9832 3093 10032
rect 3689 9832 4089 10032
rect 4685 9832 5085 10032
rect 5681 9832 6081 10032
rect 6677 9832 7077 10032
rect 7673 9832 8073 10032
rect 8669 9832 9069 10032
rect 9665 9832 10065 10032
rect 10661 9832 11061 10032
rect 11657 9832 12457 10032
rect 579 4278 779 8278
rect 1267 6752 1467 8752
rect 1819 6752 2019 8752
rect 1262 366 1462 5046
rect 1814 366 2014 2366
<< metal1 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 11672 212 12102
rect 64759 12100 64971 12118
rect 201 11581 12909 11672
rect 201 11524 426 11581
rect 201 10288 380 11524
rect 932 11524 1422 11581
rect 580 11423 778 11425
rect 580 11369 592 11423
rect 766 11369 778 11423
rect 581 10397 592 10443
rect 766 10397 777 10443
rect 201 9679 426 10288
rect 592 10031 681 10397
rect 978 10288 1376 11524
rect 1928 11524 2418 11581
rect 1576 11423 1774 11425
rect 1576 11369 1588 11423
rect 1762 11369 1774 11423
rect 1577 10397 1588 10443
rect 1762 10397 1773 10443
rect 932 10231 1422 10288
rect 913 10185 924 10231
rect 1319 10185 1422 10231
rect 592 10022 771 10031
rect 1588 10030 1668 10397
rect 1974 10288 2372 11524
rect 2924 11524 3414 11581
rect 2572 11423 2770 11425
rect 2572 11369 2584 11423
rect 2758 11369 2770 11423
rect 2573 10397 2584 10443
rect 2758 10397 2769 10443
rect 1928 10231 2418 10288
rect 1909 10185 1920 10231
rect 2315 10185 2418 10231
rect 2575 10030 2638 10397
rect 2970 10288 3368 11524
rect 3920 11524 4410 11581
rect 3568 11423 3766 11425
rect 3568 11369 3580 11423
rect 3754 11369 3766 11423
rect 3569 10397 3580 10443
rect 3754 10397 3765 10443
rect 2924 10231 3414 10288
rect 2905 10185 2916 10231
rect 3311 10185 3414 10231
rect 3571 10030 3634 10397
rect 3966 10288 4364 11524
rect 4916 11524 5406 11581
rect 4564 11423 4762 11425
rect 4564 11369 4576 11423
rect 4750 11369 4762 11423
rect 4565 10397 4576 10443
rect 4750 10397 4761 10443
rect 3920 10231 4410 10288
rect 3901 10185 3912 10231
rect 4307 10185 4410 10231
rect 4566 10030 4629 10397
rect 4962 10288 5360 11524
rect 5912 11524 6402 11581
rect 5560 11423 5758 11425
rect 5560 11369 5572 11423
rect 5746 11369 5758 11423
rect 5561 10397 5572 10443
rect 5746 10397 5757 10443
rect 4916 10231 5406 10288
rect 4897 10185 4908 10231
rect 5303 10185 5406 10231
rect 5562 10030 5625 10397
rect 5958 10288 6356 11524
rect 6908 11524 7398 11581
rect 6556 11423 6754 11425
rect 6556 11369 6568 11423
rect 6742 11369 6754 11423
rect 6557 10397 6568 10443
rect 6742 10397 6753 10443
rect 5912 10231 6402 10288
rect 5893 10185 5904 10231
rect 6299 10185 6402 10231
rect 6558 10030 6621 10397
rect 6954 10288 7352 11524
rect 7904 11524 8394 11581
rect 7552 11423 7750 11425
rect 7552 11369 7564 11423
rect 7738 11369 7750 11423
rect 6908 10231 7398 10288
rect 6889 10185 6900 10231
rect 7295 10185 7398 10231
rect 7553 10397 7564 10443
rect 7738 10397 7749 10443
rect 7553 10030 7616 10397
rect 7950 10288 8348 11524
rect 8900 11524 9390 11581
rect 8548 11423 8746 11425
rect 8548 11369 8560 11423
rect 8734 11369 8746 11423
rect 7904 10231 8394 10288
rect 7885 10185 7896 10231
rect 8291 10185 8394 10231
rect 8549 10397 8560 10443
rect 8734 10397 8745 10443
rect 8549 10030 8612 10397
rect 8946 10288 9344 11524
rect 9896 11524 10386 11581
rect 9544 11423 9742 11425
rect 9544 11369 9556 11423
rect 9730 11369 9742 11423
rect 9545 10397 9556 10443
rect 9730 10397 9741 10443
rect 8900 10231 9390 10288
rect 8881 10185 8892 10231
rect 9287 10185 9390 10231
rect 9602 10030 9665 10397
rect 9942 10288 10340 11524
rect 10892 11524 11382 11581
rect 10540 11423 10738 11425
rect 10540 11369 10552 11423
rect 10726 11369 10738 11423
rect 10541 10397 10552 10443
rect 10726 10397 10737 10443
rect 9896 10231 10386 10288
rect 9877 10185 9888 10231
rect 10283 10185 10386 10231
rect 10598 10030 10661 10397
rect 10938 10288 11336 11524
rect 11888 11524 12909 11581
rect 11536 11423 11734 11425
rect 11536 11369 11548 11423
rect 11722 11369 11734 11423
rect 11536 10397 11548 10449
rect 11661 10443 11673 10449
rect 11722 10397 11733 10443
rect 10892 10231 11382 10288
rect 11934 10288 12909 11524
rect 11888 10231 12909 10288
rect 10873 10185 10884 10231
rect 11279 10185 11439 10231
rect 12675 10185 12909 10231
rect 11548 10030 11600 10032
rect 12732 10030 12909 10185
rect 592 10019 601 10022
rect 592 9842 601 9845
rect 762 9842 771 10022
rect 592 9834 771 9842
rect 1164 10019 1668 10030
rect 1210 9845 1588 10019
rect 1634 9845 1668 10019
rect 1164 9834 1668 9845
rect 2160 10019 2638 10030
rect 2206 9845 2584 10019
rect 2630 9845 2638 10019
rect 2160 9834 2638 9845
rect 3156 10019 3634 10030
rect 3202 9845 3580 10019
rect 3626 9845 3634 10019
rect 3156 9834 3634 9845
rect 4152 10019 4629 10030
rect 4198 9845 4576 10019
rect 4622 9845 4629 10019
rect 4152 9834 4629 9845
rect 5148 10019 5625 10030
rect 5194 9845 5572 10019
rect 5618 9845 5625 10019
rect 5148 9834 5625 9845
rect 6144 10019 6621 10030
rect 6190 9845 6568 10019
rect 6614 9845 6621 10019
rect 6144 9834 6621 9845
rect 7140 10019 7616 10030
rect 7186 9845 7564 10019
rect 7610 9845 7616 10019
rect 7140 9834 7616 9845
rect 8136 10019 8612 10030
rect 8182 9845 8560 10019
rect 8606 9845 8612 10019
rect 8136 9834 8612 9845
rect 9132 10019 9665 10030
rect 9178 9845 9556 10019
rect 9602 9845 9665 10019
rect 9132 9834 9665 9845
rect 10128 10019 10661 10030
rect 10174 9845 10552 10019
rect 10598 9845 10661 10019
rect 10128 9834 10661 9845
rect 11124 10020 11600 10030
rect 11124 10019 11548 10020
rect 11170 9845 11548 10019
rect 11124 9834 11600 9845
rect 12520 10019 12909 10030
rect 12566 9845 12909 10019
rect 12520 9834 12909 9845
rect 11548 9833 11600 9834
rect 12732 9679 12909 9834
rect 201 9633 483 9679
rect 1319 9633 1479 9679
rect 2315 9633 2475 9679
rect 3311 9633 3471 9679
rect 4307 9633 4467 9679
rect 5303 9633 5463 9679
rect 6299 9633 6459 9679
rect 7295 9633 7455 9679
rect 8291 9633 8451 9679
rect 9287 9633 9447 9679
rect 10283 9633 10443 9679
rect 11279 9633 11439 9679
rect 12675 9633 12909 9679
rect 201 9471 12909 9633
rect 201 9073 1080 9471
rect 1212 9333 2280 9334
rect 64759 9333 64773 12100
rect 1212 9326 64773 9333
rect 1212 9148 1272 9326
rect 1462 9148 64773 9326
rect 1212 9134 64773 9148
rect 201 9027 2218 9073
rect 201 8970 1114 9027
rect 201 8553 1068 8970
rect 201 8496 426 8553
rect 201 4060 380 8496
rect 932 8496 1068 8553
rect 580 8341 592 8393
rect 766 8341 778 8393
rect 581 5182 777 5184
rect 572 5180 787 5182
rect 572 5100 584 5180
rect 775 5100 787 5180
rect 572 5097 787 5100
rect 581 4215 777 5097
rect 581 4169 592 4215
rect 766 4169 777 4215
rect 201 4003 426 4060
rect 978 6534 1068 8496
rect 1620 8970 1666 9027
rect 1268 8815 1280 8867
rect 1454 8815 1466 8867
rect 1268 6630 1280 6689
rect 1454 6630 1466 6689
rect 978 6477 1114 6534
rect 2172 8970 2218 9027
rect 1811 8867 2027 8880
rect 1811 8815 1823 8867
rect 2014 8815 2027 8867
rect 1811 8803 2027 8815
rect 1620 6477 1666 6534
rect 1821 6643 1832 6689
rect 2006 6643 2017 6689
rect 1821 6477 2017 6643
rect 2172 6477 2218 6534
rect 978 6431 2218 6477
rect 2266 8978 64773 9134
rect 2266 8933 3740 8978
rect 2266 8876 2491 8933
rect 978 5367 1068 6431
rect 1267 6339 1467 6350
rect 1267 6164 1278 6339
rect 1456 6258 1467 6339
rect 1456 6164 2013 6258
rect 1267 6065 2013 6164
rect 978 5321 1661 5367
rect 978 5264 1109 5321
rect 978 4060 1063 5264
rect 932 4003 1063 4060
rect 201 148 1063 4003
rect 1262 5160 1462 5162
rect 1262 5108 1275 5160
rect 1449 5108 1462 5160
rect 1262 5107 1462 5108
rect 1615 2687 1661 5321
rect 1813 4343 2013 6065
rect 1813 4215 1822 4343
rect 2002 4215 2013 4343
rect 1813 4201 2013 4215
rect 2094 2687 2184 6431
rect 2266 5860 2445 8876
rect 2957 8876 3003 8933
rect 2666 8856 2782 8857
rect 2666 8847 2678 8856
rect 2770 8847 2782 8856
rect 2666 8801 2677 8847
rect 2771 8801 2782 8847
rect 2589 8755 2635 8766
rect 2571 6103 2583 8230
rect 2589 5970 2635 5981
rect 2813 8755 2957 8766
rect 2859 5981 2957 8755
rect 2813 5970 2957 5981
rect 2666 5889 2677 5935
rect 2771 5889 2782 5935
rect 2666 5883 2678 5889
rect 2770 5883 2782 5889
rect 2666 5879 2782 5883
rect 2266 5803 2491 5860
rect 3469 8932 3740 8933
rect 64420 8932 64773 8978
rect 3469 8876 64773 8932
rect 3178 8856 3294 8857
rect 3178 8847 3190 8856
rect 3282 8847 3294 8856
rect 3178 8801 3189 8847
rect 3283 8801 3294 8847
rect 3083 8755 3147 8766
rect 3083 8754 3101 8755
rect 3083 5982 3095 8754
rect 3083 5981 3101 5982
rect 3083 5970 3147 5981
rect 3325 8755 3469 8766
rect 3371 5981 3469 8755
rect 3325 5970 3469 5981
rect 3178 5889 3189 5935
rect 3283 5889 3294 5935
rect 3178 5883 3190 5889
rect 3282 5883 3294 5889
rect 3178 5879 3294 5883
rect 2957 5803 3003 5860
rect 3515 8852 64773 8876
rect 3515 8840 34614 8852
rect 3515 8834 3870 8840
rect 23794 8834 34614 8840
rect 43980 8834 64773 8852
rect 3515 7122 3683 8834
rect 3850 8788 3861 8834
rect 23835 8788 24093 8834
rect 44067 8788 44325 8834
rect 64299 8788 64310 8834
rect 3729 8746 3815 8757
rect 3729 8739 3769 8746
rect 64345 8746 64431 8757
rect 3729 7309 3732 8739
rect 23870 8656 23881 8742
rect 24047 8656 24058 8742
rect 44102 8656 44113 8742
rect 44279 8656 44290 8742
rect 64391 8739 64431 8746
rect 3784 8641 3815 8652
rect 64345 8641 64375 8652
rect 24125 8616 33507 8628
rect 24125 8610 24133 8616
rect 44384 8616 64230 8628
rect 44384 8610 44392 8616
rect 3850 8564 3861 8610
rect 23835 8564 24093 8610
rect 44067 8564 44325 8610
rect 64299 8564 64310 8610
rect 64364 8533 64375 8641
rect 3784 8522 3815 8533
rect 64345 8522 64375 8533
rect 23870 8432 23881 8518
rect 24047 8432 24058 8518
rect 44102 8432 44113 8518
rect 44279 8432 44290 8518
rect 3784 8417 3815 8428
rect 64345 8417 64375 8428
rect 34614 8404 43980 8416
rect 3864 8392 23804 8404
rect 3864 8386 3872 8392
rect 23796 8386 23804 8392
rect 3850 8340 3861 8386
rect 23835 8340 24093 8386
rect 44067 8340 44325 8386
rect 64299 8340 64310 8386
rect 64364 8309 64375 8417
rect 3784 8298 3815 8309
rect 64345 8298 64375 8309
rect 23870 8208 23881 8294
rect 24047 8208 24058 8294
rect 44102 8208 44113 8294
rect 44279 8208 44290 8294
rect 3784 8193 3815 8204
rect 64345 8193 64375 8204
rect 24128 8168 33510 8180
rect 24128 8162 24136 8168
rect 44385 8168 64231 8180
rect 44385 8162 44392 8168
rect 3850 8116 3861 8162
rect 23835 8116 24093 8162
rect 44067 8116 44325 8162
rect 64299 8116 64310 8162
rect 64364 8085 64375 8193
rect 3784 8074 3815 8085
rect 64345 8074 64375 8085
rect 23870 7984 23881 8070
rect 24047 7984 24058 8070
rect 44102 7984 44113 8070
rect 44279 7984 44290 8070
rect 3784 7969 3815 7980
rect 64345 7969 64375 7980
rect 34611 7956 43977 7968
rect 3868 7944 23808 7956
rect 3868 7938 3876 7944
rect 23800 7938 23808 7944
rect 3850 7892 3861 7938
rect 23835 7892 24093 7938
rect 44067 7892 44325 7938
rect 64299 7892 64310 7938
rect 64364 7861 64375 7969
rect 3784 7850 3815 7861
rect 64345 7850 64375 7861
rect 23870 7760 23881 7846
rect 24047 7760 24058 7846
rect 44102 7760 44113 7846
rect 44279 7760 44290 7846
rect 3784 7745 3815 7756
rect 64345 7745 64375 7756
rect 24126 7720 33508 7732
rect 24126 7714 24134 7720
rect 44386 7720 64232 7732
rect 44386 7714 44392 7720
rect 3850 7668 3861 7714
rect 23835 7668 24093 7714
rect 44067 7668 44325 7714
rect 64299 7668 64310 7714
rect 64364 7637 64375 7745
rect 3784 7626 3815 7637
rect 64345 7626 64375 7637
rect 23870 7536 23881 7622
rect 24047 7536 24058 7622
rect 44102 7536 44113 7622
rect 44279 7536 44290 7622
rect 3784 7521 3815 7532
rect 64345 7521 64375 7532
rect 34607 7508 43973 7520
rect 3868 7496 23808 7508
rect 3868 7490 3876 7496
rect 23800 7490 23808 7496
rect 3850 7444 3861 7490
rect 23835 7444 24093 7490
rect 44067 7444 44325 7490
rect 64299 7444 64310 7490
rect 64364 7413 64375 7521
rect 3784 7402 3815 7413
rect 64345 7402 64375 7413
rect 23870 7312 23881 7398
rect 24047 7312 24058 7398
rect 44102 7312 44113 7398
rect 44279 7312 44290 7398
rect 3729 7308 3769 7309
rect 3729 7297 3815 7308
rect 64427 7309 64431 8739
rect 64391 7308 64431 7309
rect 64345 7297 64431 7308
rect 24128 7272 33510 7284
rect 24128 7266 24136 7272
rect 44381 7272 64227 7284
rect 44381 7266 44392 7272
rect 3850 7220 3861 7266
rect 23835 7220 24093 7266
rect 44067 7220 44325 7266
rect 64299 7220 64310 7266
rect 64477 7122 64773 8834
rect 3515 7076 3740 7122
rect 64420 7076 64773 7122
rect 3515 6722 3878 7076
rect 23802 6722 34608 7076
rect 43974 6722 64773 7076
rect 3515 6676 3740 6722
rect 64420 6676 64773 6722
rect 3515 6578 3878 6676
rect 23802 6578 34608 6676
rect 43974 6578 64773 6676
rect 3515 5860 3683 6578
rect 3850 6532 3861 6578
rect 23835 6532 24093 6578
rect 44067 6532 44325 6578
rect 64299 6532 64310 6578
rect 3469 5803 3683 5860
rect 2266 5757 3683 5803
rect 2266 5700 2357 5757
rect 1615 2641 2213 2687
rect 1615 2584 1661 2641
rect 1261 251 1275 303
rect 1449 251 1461 303
rect 201 91 1109 148
rect 2094 2584 2213 2641
rect 1815 2429 1827 2481
rect 2001 2429 2013 2481
rect 2094 2332 2167 2584
rect 1615 91 1661 148
rect 1816 257 1827 303
rect 2001 257 2012 303
rect 1816 91 2012 257
rect 2266 2684 2311 5700
rect 2823 5700 2869 5757
rect 2532 5671 2648 5681
rect 2532 5625 2543 5671
rect 2637 5625 2648 5671
rect 2550 5600 2621 5625
rect 2455 5579 2501 5590
rect 2405 4199 2455 4211
rect 2405 2800 2417 4199
rect 2469 2800 2501 2805
rect 2405 2794 2501 2800
rect 2550 5042 2557 5600
rect 2609 5042 2621 5600
rect 2550 2759 2621 5042
rect 2679 5579 2725 5590
rect 2731 3061 2743 5385
rect 2679 2794 2725 2805
rect 2532 2713 2543 2759
rect 2637 2713 2648 2759
rect 2532 2703 2648 2713
rect 2266 2627 2357 2684
rect 3335 5700 3683 5757
rect 3044 5671 3160 5681
rect 3044 5625 3055 5671
rect 3149 5625 3160 5671
rect 2967 5579 3013 5590
rect 2948 3056 2960 5380
rect 3078 2991 3125 5625
rect 2967 2794 3013 2805
rect 3061 2759 3073 2991
rect 3191 5579 3237 5590
rect 3243 3114 3255 5386
rect 3191 2794 3237 2805
rect 3044 2713 3055 2759
rect 3149 2713 3160 2759
rect 3044 2703 3056 2713
rect 3148 2703 3160 2713
rect 2823 2627 2869 2684
rect 3381 4866 3683 5700
rect 3729 6490 3815 6501
rect 3729 6489 3769 6490
rect 3729 5053 3732 6489
rect 64345 6490 64431 6501
rect 64391 6489 64431 6490
rect 23870 6400 23881 6486
rect 24047 6400 24058 6486
rect 44102 6400 44113 6486
rect 44279 6400 44290 6486
rect 3784 6385 3815 6396
rect 64345 6385 64375 6396
rect 24124 6360 33506 6372
rect 24124 6354 24132 6360
rect 44389 6360 64235 6372
rect 44389 6354 44392 6360
rect 3850 6308 3861 6354
rect 23835 6308 24093 6354
rect 44067 6308 44325 6354
rect 64299 6308 64310 6354
rect 64364 6277 64375 6385
rect 3784 6266 3815 6277
rect 64345 6266 64375 6277
rect 23870 6176 23881 6262
rect 24047 6176 24058 6262
rect 44102 6176 44113 6262
rect 44279 6176 44290 6262
rect 3784 6161 3815 6172
rect 64345 6161 64375 6172
rect 34613 6148 43979 6160
rect 3864 6136 23807 6148
rect 3864 6130 3872 6136
rect 23796 6130 23807 6136
rect 3850 6084 3861 6130
rect 23835 6084 24093 6130
rect 44067 6084 44325 6130
rect 64299 6084 64310 6130
rect 64364 6053 64375 6161
rect 3784 6042 3815 6053
rect 64345 6042 64375 6053
rect 23870 5952 23881 6038
rect 24047 5952 24058 6038
rect 44102 5952 44113 6038
rect 44279 5952 44290 6038
rect 3784 5937 3815 5948
rect 64345 5937 64375 5948
rect 24125 5912 33507 5924
rect 24125 5906 24133 5912
rect 44394 5912 64240 5924
rect 3850 5860 3861 5906
rect 23835 5860 24093 5906
rect 44067 5860 44325 5906
rect 64299 5860 64310 5906
rect 64364 5829 64375 5937
rect 3784 5818 3815 5829
rect 64345 5818 64375 5829
rect 23870 5728 23881 5814
rect 24047 5728 24058 5814
rect 44102 5728 44113 5814
rect 44279 5728 44290 5814
rect 3784 5713 3815 5724
rect 64345 5713 64375 5724
rect 34614 5700 43980 5712
rect 3863 5688 23810 5700
rect 3863 5682 3878 5688
rect 23802 5682 23810 5688
rect 3850 5636 3861 5682
rect 23835 5636 24093 5682
rect 44067 5636 44325 5682
rect 64299 5636 64310 5682
rect 64364 5605 64375 5713
rect 3784 5594 3815 5605
rect 64345 5594 64375 5605
rect 23870 5504 23881 5590
rect 24047 5504 24058 5590
rect 44102 5504 44113 5590
rect 44279 5504 44290 5590
rect 3784 5489 3815 5500
rect 64345 5489 64375 5500
rect 24123 5464 33505 5476
rect 24123 5458 24131 5464
rect 44396 5464 64242 5476
rect 3850 5412 3861 5458
rect 23835 5412 24093 5458
rect 44067 5412 44325 5458
rect 64299 5412 64310 5458
rect 64364 5381 64375 5489
rect 3784 5370 3815 5381
rect 64345 5370 64375 5381
rect 23870 5280 23881 5366
rect 24047 5280 24058 5366
rect 44102 5280 44113 5366
rect 44279 5280 44290 5366
rect 3784 5265 3815 5276
rect 64345 5265 64375 5276
rect 34612 5252 43978 5264
rect 3863 5240 23806 5252
rect 3863 5234 3871 5240
rect 23795 5234 23806 5240
rect 3850 5188 3861 5234
rect 23835 5188 24093 5234
rect 44067 5188 44325 5234
rect 64299 5188 64310 5234
rect 64364 5157 64375 5265
rect 3784 5146 3815 5157
rect 64345 5146 64375 5157
rect 23870 5056 23881 5142
rect 24047 5056 24058 5142
rect 44102 5056 44113 5142
rect 44279 5056 44290 5142
rect 3729 5052 3769 5053
rect 3729 5041 3815 5052
rect 64427 5053 64431 6489
rect 64391 5052 64431 5053
rect 64345 5041 64431 5052
rect 24118 5016 33507 5028
rect 24118 5010 24133 5016
rect 44387 5016 64233 5028
rect 3850 4964 3861 5010
rect 23835 4964 24093 5010
rect 44067 4964 44325 5010
rect 64299 4964 64310 5010
rect 64477 4866 64773 6578
rect 3381 4820 3740 4866
rect 64420 4820 64773 4866
rect 3381 4675 64773 4820
rect 3335 2627 3381 2684
rect 2266 2581 3381 2627
rect 3512 4628 4513 4629
rect 3512 4512 64645 4628
rect 3512 4466 3737 4512
rect 64417 4466 64645 4512
rect 3512 4387 64645 4466
rect 3512 4374 34630 4387
rect 3512 4368 3869 4374
rect 23791 4368 34630 4374
rect 43996 4368 64645 4387
rect 3512 2656 3680 4368
rect 3847 4322 3858 4368
rect 23832 4322 24090 4368
rect 44064 4322 44322 4368
rect 64296 4322 64307 4368
rect 3726 4280 3812 4291
rect 3726 4279 3766 4280
rect 64342 4280 64428 4291
rect 64388 4279 64428 4280
rect 23867 4190 23878 4276
rect 24044 4190 24055 4276
rect 44099 4190 44110 4276
rect 44276 4190 44287 4276
rect 3778 4175 3812 4186
rect 64342 4175 64376 4186
rect 24116 4150 33513 4162
rect 24116 4144 24139 4150
rect 44385 4150 64231 4162
rect 3847 4098 3858 4144
rect 23832 4098 24090 4144
rect 44064 4098 44322 4144
rect 64296 4098 64307 4144
rect 3778 4056 3812 4067
rect 64342 4056 64376 4067
rect 23867 3966 23878 4052
rect 24044 3966 24055 4052
rect 44099 3966 44110 4052
rect 44276 3966 44287 4052
rect 3778 3951 3812 3962
rect 64342 3951 64376 3962
rect 34632 3939 43998 3951
rect 3863 3926 23820 3938
rect 3863 3920 3875 3926
rect 23791 3920 23820 3926
rect 3847 3874 3858 3920
rect 23832 3874 24090 3920
rect 44064 3874 44322 3920
rect 64296 3874 64307 3920
rect 3778 3832 3812 3843
rect 64342 3832 64376 3843
rect 23867 3742 23878 3828
rect 24044 3742 24055 3828
rect 44099 3742 44110 3828
rect 44276 3742 44287 3828
rect 3778 3727 3812 3738
rect 64342 3727 64376 3738
rect 24115 3702 33512 3714
rect 24115 3696 24138 3702
rect 44389 3702 64235 3714
rect 3847 3650 3858 3696
rect 23832 3650 24090 3696
rect 44064 3650 44322 3696
rect 64296 3650 64307 3696
rect 3778 3608 3812 3619
rect 64342 3608 64376 3619
rect 23867 3518 23878 3604
rect 24044 3518 24055 3604
rect 44099 3518 44110 3604
rect 44276 3518 44287 3604
rect 3778 3503 3812 3514
rect 64342 3503 64376 3514
rect 34632 3491 43998 3503
rect 3865 3478 23822 3490
rect 3865 3472 3877 3478
rect 23791 3472 23822 3478
rect 3847 3426 3858 3472
rect 23832 3426 24090 3472
rect 44064 3426 44322 3472
rect 64296 3426 64307 3472
rect 3778 3384 3812 3395
rect 64342 3384 64376 3395
rect 23867 3294 23878 3380
rect 24044 3294 24055 3380
rect 44099 3294 44110 3380
rect 44276 3294 44287 3380
rect 3778 3279 3812 3290
rect 64342 3279 64376 3290
rect 24112 3254 33509 3266
rect 24112 3248 24135 3254
rect 44391 3254 64237 3266
rect 3847 3202 3858 3248
rect 23832 3202 24090 3248
rect 44064 3202 44322 3248
rect 64296 3202 64307 3248
rect 3778 3160 3812 3171
rect 64342 3160 64376 3171
rect 23867 3070 23878 3156
rect 24044 3070 24055 3156
rect 44099 3070 44110 3156
rect 44276 3070 44287 3156
rect 3778 3055 3812 3066
rect 64342 3055 64376 3066
rect 34631 3043 43997 3055
rect 3861 3030 23818 3042
rect 3861 3024 3873 3030
rect 23791 3024 23818 3030
rect 3847 2978 3858 3024
rect 23832 2978 24090 3024
rect 44064 2978 44322 3024
rect 64296 2978 64307 3024
rect 3778 2936 3812 2947
rect 64342 2936 64376 2947
rect 23867 2846 23878 2932
rect 24044 2846 24055 2932
rect 44099 2846 44110 2932
rect 44276 2846 44287 2932
rect 3726 2842 3766 2843
rect 3726 2831 3812 2842
rect 64388 2842 64428 2843
rect 64342 2831 64428 2842
rect 24113 2807 33510 2819
rect 24113 2800 24136 2807
rect 44386 2806 64232 2818
rect 3847 2754 3858 2800
rect 23832 2754 24090 2800
rect 44064 2754 44322 2800
rect 64296 2754 64307 2800
rect 64474 2656 64645 4368
rect 3512 2610 3737 2656
rect 64417 2610 64645 2656
rect 3512 2483 3867 2610
rect 2213 2437 3867 2483
rect 2213 2380 2512 2437
rect 2213 164 2466 2380
rect 2978 2380 3024 2437
rect 2687 2351 2803 2366
rect 2687 2305 2698 2351
rect 2792 2305 2803 2351
rect 2687 2270 2769 2305
rect 2610 2259 2769 2270
rect 2656 2258 2769 2259
rect 2667 1301 2769 2258
rect 2656 285 2769 1301
rect 2610 274 2769 285
rect 2834 2259 2978 2270
rect 2880 285 2978 2259
rect 2834 274 2978 285
rect 2687 239 2769 274
rect 2687 193 2698 239
rect 2792 193 2803 239
rect 2687 178 2803 193
rect 2213 148 2512 164
rect 2167 107 2512 148
rect 3490 2380 3867 2437
rect 3199 2351 3315 2366
rect 3199 2305 3210 2351
rect 3304 2305 3315 2351
rect 3024 2259 3168 2270
rect 3024 285 3122 2259
rect 3235 1392 3282 2305
rect 3219 1380 3282 1392
rect 3271 882 3282 1380
rect 3219 870 3282 882
rect 3024 274 3168 285
rect 3235 239 3282 870
rect 3346 2259 3392 2270
rect 3398 449 3410 2120
rect 3346 274 3392 285
rect 3199 193 3210 239
rect 3304 193 3315 239
rect 3199 178 3315 193
rect 2978 107 3024 164
rect 3536 2256 3867 2380
rect 23791 2256 34627 2610
rect 43993 2256 64645 2610
rect 3536 2210 3737 2256
rect 64417 2210 64645 2256
rect 3536 2112 3867 2210
rect 23791 2112 34627 2210
rect 43993 2131 64645 2210
rect 43994 2112 64645 2131
rect 3536 400 3680 2112
rect 3847 2066 3858 2112
rect 23832 2066 24090 2112
rect 44064 2066 44322 2112
rect 64296 2066 64307 2112
rect 3726 2024 3812 2035
rect 3726 2023 3766 2024
rect 64342 2024 64428 2035
rect 64388 2023 64428 2024
rect 23867 1934 23878 2020
rect 24044 1934 24055 2020
rect 44099 1934 44110 2020
rect 44276 1934 44287 2020
rect 3778 1919 3812 1930
rect 64342 1919 64376 1930
rect 24115 1894 33512 1906
rect 24115 1888 24138 1894
rect 44384 1894 64230 1906
rect 3847 1842 3858 1888
rect 23832 1842 24090 1888
rect 44064 1842 44322 1888
rect 64296 1842 64307 1888
rect 3778 1800 3812 1811
rect 64342 1800 64376 1811
rect 23867 1710 23878 1796
rect 24044 1710 24055 1796
rect 44099 1710 44110 1796
rect 44276 1710 44287 1796
rect 3778 1695 3812 1706
rect 64342 1695 64376 1706
rect 34633 1683 43999 1695
rect 3859 1670 23818 1682
rect 3859 1664 3871 1670
rect 23791 1664 23818 1670
rect 3847 1618 3858 1664
rect 23832 1618 24090 1664
rect 44064 1618 44322 1664
rect 64296 1618 64307 1664
rect 3778 1576 3812 1587
rect 64342 1576 64376 1587
rect 23867 1486 23878 1572
rect 24044 1486 24055 1572
rect 44099 1486 44110 1572
rect 44276 1486 44287 1572
rect 3778 1471 3812 1482
rect 64342 1471 64376 1482
rect 24116 1446 33513 1458
rect 24116 1440 24139 1446
rect 44385 1446 64231 1458
rect 3847 1394 3858 1440
rect 23832 1394 24090 1440
rect 44064 1394 44322 1440
rect 64296 1394 64307 1440
rect 3778 1352 3812 1363
rect 64342 1352 64376 1363
rect 23867 1262 23878 1348
rect 24044 1262 24055 1348
rect 44099 1262 44110 1348
rect 44276 1262 44287 1348
rect 3778 1247 3812 1258
rect 64342 1247 64376 1258
rect 34643 1235 44009 1247
rect 3858 1222 23818 1234
rect 3858 1216 3871 1222
rect 23791 1216 23818 1222
rect 3847 1170 3858 1216
rect 23832 1170 24090 1216
rect 44064 1170 44322 1216
rect 64296 1170 64307 1216
rect 3778 1128 3812 1139
rect 64342 1128 64376 1139
rect 23867 1038 23878 1124
rect 24044 1038 24055 1124
rect 44099 1038 44110 1124
rect 44276 1038 44287 1124
rect 3778 1023 3812 1034
rect 64342 1023 64376 1034
rect 24112 998 33509 1010
rect 24112 992 24135 998
rect 44390 998 64236 1010
rect 3847 946 3858 992
rect 23832 946 24090 992
rect 44064 946 44322 992
rect 64296 946 64307 992
rect 3778 904 3812 915
rect 64342 904 64376 915
rect 23867 814 23878 900
rect 24044 814 24055 900
rect 44099 814 44110 900
rect 44276 814 44287 900
rect 3778 799 3812 810
rect 64342 799 64376 810
rect 34626 787 43992 799
rect 3857 774 23806 786
rect 3857 768 3868 774
rect 23783 768 23806 774
rect 3847 722 3858 768
rect 23832 722 24090 768
rect 44064 722 44322 768
rect 64296 722 64307 768
rect 3778 680 3812 691
rect 64342 680 64376 691
rect 23867 590 23878 676
rect 24044 590 24055 676
rect 44099 590 44110 676
rect 44276 590 44287 676
rect 3726 586 3766 587
rect 3726 575 3812 586
rect 64388 586 64428 587
rect 64342 575 64428 586
rect 24132 550 33506 562
rect 44381 550 64227 562
rect 3847 498 3858 544
rect 23832 498 24090 544
rect 44064 498 44322 544
rect 64296 498 64307 544
rect 64474 400 64645 2112
rect 3536 354 3737 400
rect 64417 354 64645 400
rect 3536 164 64645 354
rect 3490 107 64645 164
rect 2167 91 64645 107
rect 201 16 64645 91
rect 0 1 64645 16
rect 64759 14 64773 4675
rect 64959 14 64971 12100
rect 64759 1 64971 14
rect 0 0 2265 1
rect 2466 0 64645 1
<< via1 >>
rect 15 16 201 12102
rect 592 11415 766 11423
rect 592 11371 766 11415
rect 1588 11415 1762 11423
rect 1588 11371 1762 11415
rect 2584 11415 2758 11423
rect 2584 11371 2758 11415
rect 3580 11415 3754 11423
rect 3580 11371 3754 11415
rect 4576 11415 4750 11423
rect 4576 11371 4750 11415
rect 5572 11415 5746 11423
rect 5572 11371 5746 11415
rect 6568 11415 6742 11423
rect 6568 11371 6742 11415
rect 7564 11415 7738 11423
rect 7564 11371 7738 11415
rect 8560 11415 8734 11423
rect 8560 11371 8734 11415
rect 9556 11415 9730 11423
rect 9556 11371 9730 11415
rect 10552 11415 10726 11423
rect 10552 11371 10726 11415
rect 11548 11415 11722 11423
rect 11548 11371 11722 11415
rect 11548 10443 11661 10449
rect 11548 10397 11661 10443
rect 601 10019 762 10022
rect 601 9845 638 10019
rect 638 9845 762 10019
rect 601 9842 762 9845
rect 11548 10019 11600 10020
rect 11548 9845 11594 10019
rect 11594 9845 11600 10019
rect 1272 9148 1462 9326
rect 592 8387 766 8393
rect 592 8341 766 8387
rect 584 5100 775 5180
rect 1280 8861 1454 8867
rect 1280 8815 1454 8861
rect 1280 6643 1454 6689
rect 1280 6630 1454 6643
rect 1823 8861 2014 8867
rect 1823 8815 1832 8861
rect 1832 8815 2006 8861
rect 2006 8815 2014 8861
rect 1278 6164 1456 6339
rect 1275 5155 1449 5160
rect 1275 5109 1449 5155
rect 1275 5108 1449 5109
rect 1822 4215 2002 4343
rect 2678 8847 2770 8856
rect 2678 8804 2770 8847
rect 2583 6103 2589 8230
rect 2589 6103 2635 8230
rect 2678 5889 2770 5935
rect 2678 5883 2770 5889
rect 3190 8847 3282 8856
rect 3190 8804 3282 8847
rect 3095 5982 3101 8754
rect 3101 5982 3147 8754
rect 3190 5889 3282 5935
rect 3190 5883 3282 5889
rect 3870 8834 23794 8840
rect 34614 8834 43980 8852
rect 3870 8788 23794 8834
rect 34614 8788 43980 8834
rect 3732 8652 3769 8739
rect 3769 8652 3784 8739
rect 23882 8656 23927 8742
rect 23927 8656 24001 8742
rect 24001 8656 24046 8742
rect 44114 8656 44159 8742
rect 44159 8656 44233 8742
rect 44233 8656 44278 8742
rect 3732 8522 3784 8652
rect 64375 8652 64391 8739
rect 64391 8652 64427 8739
rect 24133 8610 33507 8616
rect 44392 8610 64230 8616
rect 24133 8564 33507 8610
rect 44392 8564 64230 8610
rect 3732 8428 3769 8522
rect 3769 8428 3784 8522
rect 64375 8522 64427 8652
rect 23882 8432 23927 8518
rect 23927 8432 24001 8518
rect 24001 8432 24046 8518
rect 44114 8432 44159 8518
rect 44159 8432 44233 8518
rect 44233 8432 44278 8518
rect 3732 8298 3784 8428
rect 64375 8428 64391 8522
rect 64391 8428 64427 8522
rect 3872 8386 23796 8392
rect 34614 8386 43980 8404
rect 3872 8340 23796 8386
rect 34614 8340 43980 8386
rect 3732 8204 3769 8298
rect 3769 8204 3784 8298
rect 64375 8298 64427 8428
rect 23882 8208 23927 8294
rect 23927 8208 24001 8294
rect 24001 8208 24046 8294
rect 44114 8208 44159 8294
rect 44159 8208 44233 8294
rect 44233 8208 44278 8294
rect 3732 8074 3784 8204
rect 64375 8204 64391 8298
rect 64391 8204 64427 8298
rect 24136 8162 33510 8168
rect 44392 8162 64231 8168
rect 24136 8116 33510 8162
rect 44392 8116 64231 8162
rect 3732 7980 3769 8074
rect 3769 7980 3784 8074
rect 64375 8074 64427 8204
rect 23882 7984 23927 8070
rect 23927 7984 24001 8070
rect 24001 7984 24046 8070
rect 44114 7984 44159 8070
rect 44159 7984 44233 8070
rect 44233 7984 44278 8070
rect 3732 7850 3784 7980
rect 64375 7980 64391 8074
rect 64391 7980 64427 8074
rect 3876 7938 23800 7944
rect 34611 7938 43977 7956
rect 3876 7892 23800 7938
rect 34611 7892 43977 7938
rect 3732 7756 3769 7850
rect 3769 7756 3784 7850
rect 64375 7850 64427 7980
rect 23882 7760 23927 7846
rect 23927 7760 24001 7846
rect 24001 7760 24046 7846
rect 44114 7760 44159 7846
rect 44159 7760 44233 7846
rect 44233 7760 44278 7846
rect 3732 7626 3784 7756
rect 64375 7756 64391 7850
rect 64391 7756 64427 7850
rect 24134 7714 33508 7720
rect 44392 7714 64232 7720
rect 24134 7668 33508 7714
rect 44392 7668 64232 7714
rect 3732 7532 3769 7626
rect 3769 7532 3784 7626
rect 64375 7626 64427 7756
rect 23882 7536 23927 7622
rect 23927 7536 24001 7622
rect 24001 7536 24046 7622
rect 44114 7536 44159 7622
rect 44159 7536 44233 7622
rect 44233 7536 44278 7622
rect 3732 7402 3784 7532
rect 64375 7532 64391 7626
rect 64391 7532 64427 7626
rect 3876 7490 23800 7496
rect 34607 7490 43973 7508
rect 3876 7444 23800 7490
rect 34607 7444 43973 7490
rect 3732 7309 3769 7402
rect 3769 7309 3784 7402
rect 64375 7402 64427 7532
rect 23882 7312 23927 7398
rect 23927 7312 24001 7398
rect 24001 7312 24046 7398
rect 44114 7312 44159 7398
rect 44159 7312 44233 7398
rect 44233 7312 44278 7398
rect 64375 7309 64391 7402
rect 64391 7309 64427 7402
rect 24136 7266 33510 7272
rect 44392 7266 64227 7272
rect 24136 7220 33510 7266
rect 44392 7220 64227 7266
rect 3878 7076 23802 7115
rect 34608 7076 43974 7116
rect 3878 6722 23802 7076
rect 34608 6722 43974 7076
rect 3878 6676 23802 6722
rect 34608 6676 43974 6722
rect 3878 6578 23802 6676
rect 34608 6578 43974 6676
rect 3878 6532 23802 6578
rect 34608 6532 43974 6578
rect 1275 257 1449 303
rect 1275 251 1449 257
rect 1827 2475 2001 2481
rect 1827 2429 2001 2475
rect 2417 2805 2455 4199
rect 2455 2805 2469 4199
rect 2417 2800 2469 2805
rect 2557 5042 2609 5600
rect 2679 3061 2725 5385
rect 2725 3061 2731 5385
rect 2960 3056 2967 5380
rect 2967 3056 3012 5380
rect 3073 2759 3125 2991
rect 3191 3114 3237 5386
rect 3237 3114 3243 5386
rect 3056 2713 3148 2759
rect 3056 2703 3148 2713
rect 3732 6396 3769 6489
rect 3769 6396 3784 6489
rect 23882 6400 23927 6486
rect 23927 6400 24001 6486
rect 24001 6400 24046 6486
rect 44114 6400 44159 6486
rect 44159 6400 44233 6486
rect 44233 6400 44278 6486
rect 3732 6266 3784 6396
rect 64375 6396 64391 6489
rect 64391 6396 64427 6489
rect 24132 6354 33506 6360
rect 44392 6354 64235 6360
rect 24132 6308 33506 6354
rect 44392 6308 64235 6354
rect 3732 6172 3769 6266
rect 3769 6172 3784 6266
rect 64375 6266 64427 6396
rect 23882 6176 23927 6262
rect 23927 6176 24001 6262
rect 24001 6176 24046 6262
rect 44114 6176 44159 6262
rect 44159 6176 44233 6262
rect 44233 6176 44278 6262
rect 3732 6042 3784 6172
rect 64375 6172 64391 6266
rect 64391 6172 64427 6266
rect 3872 6130 23796 6136
rect 34613 6130 43979 6148
rect 3872 6084 23796 6130
rect 34613 6084 43979 6130
rect 3732 5948 3769 6042
rect 3769 5948 3784 6042
rect 64375 6042 64427 6172
rect 23882 5952 23927 6038
rect 23927 5952 24001 6038
rect 24001 5952 24046 6038
rect 44114 5952 44159 6038
rect 44159 5952 44233 6038
rect 44233 5952 44278 6038
rect 3732 5818 3784 5948
rect 64375 5948 64391 6042
rect 64391 5948 64427 6042
rect 24133 5906 33507 5912
rect 44394 5906 64240 5912
rect 24133 5860 33507 5906
rect 44394 5860 64240 5906
rect 3732 5724 3769 5818
rect 3769 5724 3784 5818
rect 64375 5818 64427 5948
rect 23882 5728 23927 5814
rect 23927 5728 24001 5814
rect 24001 5728 24046 5814
rect 44114 5728 44159 5814
rect 44159 5728 44233 5814
rect 44233 5728 44278 5814
rect 3732 5594 3784 5724
rect 64375 5724 64391 5818
rect 64391 5724 64427 5818
rect 3878 5682 23802 5688
rect 34614 5682 43980 5700
rect 3878 5636 23802 5682
rect 34614 5636 43980 5682
rect 3732 5500 3769 5594
rect 3769 5500 3784 5594
rect 64375 5594 64427 5724
rect 23882 5504 23927 5590
rect 23927 5504 24001 5590
rect 24001 5504 24046 5590
rect 44114 5504 44159 5590
rect 44159 5504 44233 5590
rect 44233 5504 44278 5590
rect 3732 5370 3784 5500
rect 64375 5500 64391 5594
rect 64391 5500 64427 5594
rect 24131 5458 33505 5464
rect 44396 5458 64242 5464
rect 24131 5412 33505 5458
rect 44396 5412 64242 5458
rect 3732 5276 3769 5370
rect 3769 5276 3784 5370
rect 64375 5370 64427 5500
rect 23882 5280 23927 5366
rect 23927 5280 24001 5366
rect 24001 5280 24046 5366
rect 44114 5280 44159 5366
rect 44159 5280 44233 5366
rect 44233 5280 44278 5366
rect 3732 5146 3784 5276
rect 64375 5276 64391 5370
rect 64391 5276 64427 5370
rect 3871 5234 23795 5240
rect 34612 5234 43978 5252
rect 3871 5188 23795 5234
rect 34612 5188 43978 5234
rect 3732 5053 3769 5146
rect 3769 5053 3784 5146
rect 64375 5146 64427 5276
rect 23882 5056 23927 5142
rect 23927 5056 24001 5142
rect 24001 5056 24046 5142
rect 44114 5056 44159 5142
rect 44159 5056 44233 5142
rect 44233 5056 44278 5142
rect 64375 5053 64391 5146
rect 64391 5053 64427 5146
rect 24133 5010 33507 5016
rect 44387 5010 64233 5016
rect 24133 4964 33507 5010
rect 44387 4964 64233 5010
rect 3869 4368 23791 4374
rect 34630 4368 43996 4387
rect 3869 4322 23791 4368
rect 34630 4322 43996 4368
rect 3726 4186 3766 4279
rect 3766 4186 3778 4279
rect 23879 4190 23924 4276
rect 23924 4190 23998 4276
rect 23998 4190 24043 4276
rect 44111 4190 44156 4276
rect 44156 4190 44230 4276
rect 44230 4190 44275 4276
rect 3726 4056 3778 4186
rect 64376 4186 64388 4279
rect 64388 4186 64428 4279
rect 24139 4144 33513 4150
rect 44385 4144 64231 4150
rect 24139 4098 33513 4144
rect 44385 4098 64231 4144
rect 3726 3962 3766 4056
rect 3766 3962 3778 4056
rect 64376 4056 64428 4186
rect 23879 3966 23924 4052
rect 23924 3966 23998 4052
rect 23998 3966 24043 4052
rect 44111 3966 44156 4052
rect 44156 3966 44230 4052
rect 44230 3966 44275 4052
rect 3726 3832 3778 3962
rect 64376 3962 64388 4056
rect 64388 3962 64428 4056
rect 3875 3920 23791 3926
rect 34632 3920 43998 3939
rect 3875 3874 23791 3920
rect 34632 3874 43998 3920
rect 3726 3738 3766 3832
rect 3766 3738 3778 3832
rect 64376 3832 64428 3962
rect 23879 3742 23924 3828
rect 23924 3742 23998 3828
rect 23998 3742 24043 3828
rect 44111 3742 44156 3828
rect 44156 3742 44230 3828
rect 44230 3742 44275 3828
rect 3726 3608 3778 3738
rect 64376 3738 64388 3832
rect 64388 3738 64428 3832
rect 24138 3696 33512 3702
rect 44389 3696 64235 3702
rect 24138 3650 33512 3696
rect 44389 3650 64235 3696
rect 3726 3514 3766 3608
rect 3766 3514 3778 3608
rect 64376 3608 64428 3738
rect 23879 3518 23924 3604
rect 23924 3518 23998 3604
rect 23998 3518 24043 3604
rect 44111 3518 44156 3604
rect 44156 3518 44230 3604
rect 44230 3518 44275 3604
rect 3726 3384 3778 3514
rect 64376 3514 64388 3608
rect 64388 3514 64428 3608
rect 3877 3472 23791 3478
rect 34632 3472 43998 3491
rect 3877 3426 23791 3472
rect 34632 3426 43998 3472
rect 3726 3290 3766 3384
rect 3766 3290 3778 3384
rect 64376 3384 64428 3514
rect 23879 3294 23924 3380
rect 23924 3294 23998 3380
rect 23998 3294 24043 3380
rect 44111 3294 44156 3380
rect 44156 3294 44230 3380
rect 44230 3294 44275 3380
rect 3726 3160 3778 3290
rect 64376 3290 64388 3384
rect 64388 3290 64428 3384
rect 24135 3248 33509 3254
rect 44391 3248 64237 3254
rect 24135 3202 33509 3248
rect 44391 3202 64237 3248
rect 3726 3066 3766 3160
rect 3766 3066 3778 3160
rect 64376 3160 64428 3290
rect 23879 3070 23924 3156
rect 23924 3070 23998 3156
rect 23998 3070 24043 3156
rect 44111 3070 44156 3156
rect 44156 3070 44230 3156
rect 44230 3070 44275 3156
rect 3726 2936 3778 3066
rect 64376 3066 64388 3160
rect 64388 3066 64428 3160
rect 3873 3024 23791 3030
rect 34631 3024 43997 3043
rect 3873 2978 23791 3024
rect 34631 2978 43997 3024
rect 3726 2843 3766 2936
rect 3766 2843 3778 2936
rect 64376 2936 64428 3066
rect 23879 2846 23924 2932
rect 23924 2846 23998 2932
rect 23998 2846 24043 2932
rect 44111 2846 44156 2932
rect 44156 2846 44230 2932
rect 44230 2846 44275 2932
rect 64376 2843 64388 2936
rect 64388 2843 64428 2936
rect 24136 2800 33510 2807
rect 44386 2800 64232 2806
rect 24136 2755 33510 2800
rect 44386 2754 64232 2800
rect 3867 2610 23791 2649
rect 34627 2610 43993 2650
rect 2615 1301 2656 2258
rect 2656 1301 2667 2258
rect 3219 882 3271 1380
rect 3346 449 3392 2120
rect 3392 449 3398 2120
rect 3867 2256 23791 2610
rect 34627 2256 43993 2610
rect 3867 2210 23791 2256
rect 34627 2210 43993 2256
rect 3867 2112 23791 2210
rect 34627 2131 43993 2210
rect 34627 2112 43994 2131
rect 3867 2066 23791 2112
rect 34627 2066 43994 2112
rect 3726 1930 3766 2023
rect 3766 1930 3778 2023
rect 23879 1934 23924 2020
rect 23924 1934 23998 2020
rect 23998 1934 24043 2020
rect 44111 1934 44156 2020
rect 44156 1934 44230 2020
rect 44230 1934 44275 2020
rect 3726 1800 3778 1930
rect 64376 1930 64388 2023
rect 64388 1930 64428 2023
rect 24138 1888 33512 1894
rect 44384 1888 64230 1894
rect 24138 1842 33512 1888
rect 44384 1842 64230 1888
rect 3726 1706 3766 1800
rect 3766 1706 3778 1800
rect 64376 1800 64428 1930
rect 23879 1710 23924 1796
rect 23924 1710 23998 1796
rect 23998 1710 24043 1796
rect 44111 1710 44156 1796
rect 44156 1710 44230 1796
rect 44230 1710 44275 1796
rect 3726 1576 3778 1706
rect 64376 1706 64388 1800
rect 64388 1706 64428 1800
rect 3871 1664 23791 1670
rect 34633 1664 43999 1683
rect 3871 1618 23791 1664
rect 34633 1618 43999 1664
rect 3726 1482 3766 1576
rect 3766 1482 3778 1576
rect 64376 1576 64428 1706
rect 23879 1486 23924 1572
rect 23924 1486 23998 1572
rect 23998 1486 24043 1572
rect 44111 1486 44156 1572
rect 44156 1486 44230 1572
rect 44230 1486 44275 1572
rect 3726 1352 3778 1482
rect 64376 1482 64388 1576
rect 64388 1482 64428 1576
rect 24139 1440 33513 1446
rect 44385 1440 64231 1446
rect 24139 1394 33513 1440
rect 44385 1394 64231 1440
rect 3726 1258 3766 1352
rect 3766 1258 3778 1352
rect 64376 1352 64428 1482
rect 23879 1262 23924 1348
rect 23924 1262 23998 1348
rect 23998 1262 24043 1348
rect 44111 1262 44156 1348
rect 44156 1262 44230 1348
rect 44230 1262 44275 1348
rect 3726 1128 3778 1258
rect 64376 1258 64388 1352
rect 64388 1258 64428 1352
rect 3871 1216 23791 1222
rect 34643 1216 44009 1235
rect 3871 1170 23791 1216
rect 34643 1170 44009 1216
rect 3726 1034 3766 1128
rect 3766 1034 3778 1128
rect 64376 1128 64428 1258
rect 23879 1038 23924 1124
rect 23924 1038 23998 1124
rect 23998 1038 24043 1124
rect 44111 1038 44156 1124
rect 44156 1038 44230 1124
rect 44230 1038 44275 1124
rect 3726 904 3778 1034
rect 64376 1034 64388 1128
rect 64388 1034 64428 1128
rect 24135 992 33509 998
rect 44390 992 64236 998
rect 24135 946 33509 992
rect 44390 946 64236 992
rect 3726 810 3766 904
rect 3766 810 3778 904
rect 64376 904 64428 1034
rect 23879 814 23924 900
rect 23924 814 23998 900
rect 23998 814 24043 900
rect 44111 814 44156 900
rect 44156 814 44230 900
rect 44230 814 44275 900
rect 3726 680 3778 810
rect 64376 810 64388 904
rect 64388 810 64428 904
rect 3868 768 23783 774
rect 34626 768 43992 787
rect 3868 722 23783 768
rect 34626 722 43992 768
rect 3726 587 3766 680
rect 3766 587 3778 680
rect 64376 680 64428 810
rect 23879 590 23924 676
rect 23924 590 23998 676
rect 23998 590 24043 676
rect 44111 590 44156 676
rect 44156 590 44230 676
rect 44230 590 44275 676
rect 64376 587 64388 680
rect 64388 587 64428 680
rect 24132 544 33506 550
rect 44381 544 64227 550
rect 24132 498 33506 544
rect 44381 498 64227 544
rect 64773 14 64959 12100
<< metal2 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 16 212 12102
rect 580 11423 778 12117
rect 580 11371 592 11423
rect 766 11371 778 11423
rect 580 11369 778 11371
rect 1576 11423 1774 12117
rect 1576 11371 1588 11423
rect 1762 11371 1774 11423
rect 1576 11369 1774 11371
rect 2572 11423 2770 12117
rect 2572 11371 2584 11423
rect 2758 11371 2770 11423
rect 2572 11369 2770 11371
rect 3568 11423 3766 12117
rect 3568 11371 3580 11423
rect 3754 11371 3766 11423
rect 3568 11369 3766 11371
rect 4564 11423 4762 12117
rect 4564 11371 4576 11423
rect 4750 11371 4762 11423
rect 4564 11369 4762 11371
rect 5560 11423 5758 12117
rect 5560 11371 5572 11423
rect 5746 11371 5758 11423
rect 5560 11369 5758 11371
rect 6556 11423 6754 12117
rect 6556 11371 6568 11423
rect 6742 11371 6754 11423
rect 6556 11369 6754 11371
rect 7552 11423 7750 12117
rect 7552 11371 7564 11423
rect 7738 11371 7750 11423
rect 7552 11369 7750 11371
rect 8548 11423 8746 12117
rect 8548 11371 8560 11423
rect 8734 11371 8746 11423
rect 8548 11369 8746 11371
rect 9544 11423 9742 12117
rect 9544 11371 9556 11423
rect 9730 11371 9742 11423
rect 9544 11369 9742 11371
rect 10540 11423 10738 12117
rect 10540 11371 10552 11423
rect 10726 11371 10738 11423
rect 10540 11369 10738 11371
rect 11536 11423 11734 12117
rect 51536 11510 51733 12118
rect 11536 11371 11548 11423
rect 11722 11371 11734 11423
rect 11536 11369 11734 11371
rect 51535 11369 51733 11510
rect 64759 12100 64971 12118
rect 51535 10998 51732 11369
rect 51535 10774 51536 10998
rect 51731 10774 51732 10998
rect 51535 10761 51732 10774
rect 11524 10449 11673 10453
rect 11524 10397 11548 10449
rect 11661 10397 11673 10449
rect 11524 10384 11673 10397
rect 578 10022 779 10051
rect 578 9842 601 10022
rect 762 9842 779 10022
rect 578 8393 779 9842
rect 11524 10020 11610 10384
rect 11524 9845 11548 10020
rect 11600 9845 11610 10020
rect 11524 9821 11610 9845
rect 1264 9326 1468 9338
rect 1264 9148 1272 9326
rect 1462 9148 1468 9326
rect 1264 8867 1468 9148
rect 3705 8947 64445 9070
rect 3705 8884 3786 8947
rect 1264 8815 1280 8867
rect 1454 8815 1468 8867
rect 1264 8810 1468 8815
rect 1808 8867 3786 8884
rect 1808 8815 1823 8867
rect 2014 8856 3786 8867
rect 2014 8815 2678 8856
rect 1808 8804 2678 8815
rect 2770 8804 3190 8856
rect 3282 8804 3786 8856
rect 1808 8799 3786 8804
rect 2665 8798 3786 8799
rect 578 8341 592 8393
rect 766 8341 779 8393
rect 578 8337 779 8341
rect 3066 8754 3149 8798
rect 2550 8230 2643 8240
rect 1267 6689 1467 6695
rect 1267 6630 1280 6689
rect 1454 6630 1467 6689
rect 1267 6339 1467 6630
rect 1267 6164 1278 6339
rect 1456 6164 1467 6339
rect 1267 6152 1467 6164
rect 2550 6103 2583 8230
rect 2635 6103 2643 8230
rect 2550 6094 2643 6103
rect 2550 5799 2620 6094
rect 3066 5982 3095 8754
rect 3147 5982 3149 8754
rect 2676 5939 2785 5947
rect 3066 5939 3149 5982
rect 3705 8739 3786 8798
rect 3705 7309 3732 8739
rect 3784 7309 3786 8739
rect 3705 6489 3786 7309
rect 3705 5939 3732 6489
rect 2676 5935 3732 5939
rect 2676 5883 2678 5935
rect 2770 5883 3190 5935
rect 3282 5883 3732 5935
rect 2676 5874 3732 5883
rect 2676 5871 2785 5874
rect 2550 5727 2745 5799
rect 2530 5600 2616 5612
rect 2530 5182 2557 5600
rect 572 5180 2557 5182
rect 572 5100 584 5180
rect 775 5160 2557 5180
rect 775 5108 1275 5160
rect 1449 5108 2557 5160
rect 775 5100 2557 5108
rect 572 5097 2557 5100
rect 2530 5042 2557 5097
rect 2609 5042 2616 5600
rect 2530 5030 2616 5042
rect 2672 5397 2745 5727
rect 2672 5385 3024 5397
rect 1814 4343 2615 4352
rect 1814 4215 1822 4343
rect 2002 4267 2615 4343
rect 2002 4215 2013 4267
rect 1814 2481 2013 4215
rect 1814 2429 1827 2481
rect 2001 2429 2013 2481
rect 1814 2427 2013 2429
rect 2391 4199 2474 4211
rect 2391 2800 2417 4199
rect 2469 2800 2474 4199
rect 2530 3420 2615 4267
rect 2530 2993 2616 3420
rect 2672 3061 2679 5385
rect 2731 5380 3024 5385
rect 2731 3061 2960 5380
rect 2672 3056 2960 3061
rect 3012 3056 3024 5380
rect 3183 5386 3258 5394
rect 3183 3114 3191 5386
rect 3243 3995 3258 5386
rect 3705 5053 3732 5874
rect 3784 5053 3786 6489
rect 3858 8840 23806 8865
rect 3858 8788 3870 8840
rect 23794 8788 23806 8840
rect 3858 8392 23806 8788
rect 3858 8340 3872 8392
rect 23796 8340 23806 8392
rect 3858 7944 23806 8340
rect 3858 7892 3876 7944
rect 23800 7892 23806 7944
rect 3858 7496 23806 7892
rect 3858 7444 3876 7496
rect 23800 7444 23806 7496
rect 3858 7115 23806 7444
rect 3858 6532 3878 7115
rect 23802 6532 23806 7115
rect 3858 6136 23806 6532
rect 3858 6084 3872 6136
rect 23796 6084 23806 6136
rect 3858 5688 23806 6084
rect 3858 5636 3878 5688
rect 23802 5636 23806 5688
rect 3858 5240 23806 5636
rect 3858 5188 3871 5240
rect 23795 5188 23806 5240
rect 3858 5164 23806 5188
rect 23870 8742 24058 8947
rect 23870 8656 23882 8742
rect 24046 8656 24058 8742
rect 34595 8852 43996 8874
rect 34595 8788 34614 8852
rect 43980 8788 43996 8852
rect 23870 8518 24058 8656
rect 23870 8432 23882 8518
rect 24046 8432 24058 8518
rect 23870 8294 24058 8432
rect 23870 8208 23882 8294
rect 24046 8208 24058 8294
rect 23870 8070 24058 8208
rect 23870 7984 23882 8070
rect 24046 7984 24058 8070
rect 23870 7846 24058 7984
rect 23870 7760 23882 7846
rect 24046 7760 24058 7846
rect 23870 7622 24058 7760
rect 23870 7536 23882 7622
rect 24046 7536 24058 7622
rect 23870 7398 24058 7536
rect 23870 7312 23882 7398
rect 24046 7312 24058 7398
rect 23870 6486 24058 7312
rect 23870 6400 23882 6486
rect 24046 6400 24058 6486
rect 23870 6262 24058 6400
rect 23870 6176 23882 6262
rect 24046 6176 24058 6262
rect 23870 6038 24058 6176
rect 23870 5952 23882 6038
rect 24046 5952 24058 6038
rect 23870 5814 24058 5952
rect 23870 5728 23882 5814
rect 24046 5728 24058 5814
rect 23870 5590 24058 5728
rect 23870 5504 23882 5590
rect 24046 5504 24058 5590
rect 23870 5366 24058 5504
rect 23870 5280 23882 5366
rect 24046 5280 24058 5366
rect 3705 5016 3786 5053
rect 23870 5142 24058 5280
rect 23870 5056 23882 5142
rect 24046 5056 24058 5142
rect 23870 5045 24058 5056
rect 24118 8616 33518 8679
rect 24118 8564 24133 8616
rect 33507 8564 33518 8616
rect 24118 8168 33518 8564
rect 24118 8116 24136 8168
rect 33510 8116 33518 8168
rect 24118 7720 33518 8116
rect 24118 7668 24134 7720
rect 33508 7668 33518 7720
rect 24118 7272 33518 7668
rect 24118 7220 24136 7272
rect 33510 7220 33518 7272
rect 24118 6360 33518 7220
rect 24118 6308 24132 6360
rect 33506 6308 33518 6360
rect 24118 5912 33518 6308
rect 24118 5860 24133 5912
rect 33507 5860 33518 5912
rect 24118 5464 33518 5860
rect 24118 5412 24131 5464
rect 33505 5412 33518 5464
rect 24118 5016 33518 5412
rect 34595 8404 43996 8788
rect 34595 8340 34614 8404
rect 43980 8340 43996 8404
rect 34595 7956 43996 8340
rect 34595 7892 34611 7956
rect 43977 7892 43996 7956
rect 34595 7508 43996 7892
rect 34595 7444 34607 7508
rect 43973 7444 43996 7508
rect 34595 7116 43996 7444
rect 34595 6532 34608 7116
rect 43974 6532 43996 7116
rect 34595 6148 43996 6532
rect 34595 6084 34613 6148
rect 43979 6084 43996 6148
rect 34595 5700 43996 6084
rect 34595 5636 34614 5700
rect 43980 5636 43996 5700
rect 34595 5252 43996 5636
rect 34595 5188 34612 5252
rect 43978 5188 43996 5252
rect 34595 5176 43996 5188
rect 44102 8742 44290 8947
rect 44102 8656 44114 8742
rect 44278 8656 44290 8742
rect 64364 8739 64445 8947
rect 44102 8518 44290 8656
rect 44102 8432 44114 8518
rect 44278 8432 44290 8518
rect 44102 8294 44290 8432
rect 44102 8208 44114 8294
rect 44278 8208 44290 8294
rect 44102 8070 44290 8208
rect 44102 7984 44114 8070
rect 44278 7984 44290 8070
rect 44102 7846 44290 7984
rect 44102 7760 44114 7846
rect 44278 7760 44290 7846
rect 44102 7622 44290 7760
rect 44102 7536 44114 7622
rect 44278 7536 44290 7622
rect 44102 7398 44290 7536
rect 44102 7312 44114 7398
rect 44278 7312 44290 7398
rect 44102 6486 44290 7312
rect 44102 6400 44114 6486
rect 44278 6400 44290 6486
rect 44102 6262 44290 6400
rect 44102 6176 44114 6262
rect 44278 6176 44290 6262
rect 44102 6038 44290 6176
rect 44102 5952 44114 6038
rect 44278 5952 44290 6038
rect 44102 5814 44290 5952
rect 44102 5728 44114 5814
rect 44278 5728 44290 5814
rect 44102 5590 44290 5728
rect 44102 5504 44114 5590
rect 44278 5504 44290 5590
rect 44102 5366 44290 5504
rect 44102 5280 44114 5366
rect 44278 5280 44290 5366
rect 44102 5142 44290 5280
rect 44102 5056 44114 5142
rect 44278 5056 44290 5142
rect 44102 5050 44290 5056
rect 44381 8616 64267 8679
rect 44381 8564 44392 8616
rect 64230 8564 64267 8616
rect 44381 8364 64267 8564
rect 44381 8168 51556 8364
rect 52428 8168 64267 8364
rect 44381 8116 44392 8168
rect 64231 8116 64267 8168
rect 44381 7720 51556 8116
rect 52428 7720 64267 8116
rect 44381 7668 44392 7720
rect 64232 7668 64267 7720
rect 44381 7464 51556 7668
rect 52428 7464 64267 7668
rect 44381 7272 64267 7464
rect 44381 7220 44392 7272
rect 64227 7220 64267 7272
rect 44381 6360 64267 7220
rect 44381 6308 44392 6360
rect 64235 6308 64267 6360
rect 44381 5912 64267 6308
rect 44381 5860 44394 5912
rect 64240 5860 64267 5912
rect 44381 5464 64267 5860
rect 44381 5412 44396 5464
rect 64242 5412 64267 5464
rect 24118 4964 24133 5016
rect 33507 4990 33518 5016
rect 44381 5016 64267 5412
rect 44381 4990 44387 5016
rect 33507 4964 44387 4990
rect 64233 4964 64267 5016
rect 64364 7309 64375 8739
rect 64427 7309 64445 8739
rect 64364 6489 64445 7309
rect 64364 5053 64375 6489
rect 64427 5053 64445 6489
rect 64364 5008 64445 5053
rect 24118 4482 64267 4964
rect 3851 4374 23793 4408
rect 3851 4322 3869 4374
rect 23791 4322 23793 4374
rect 3659 4279 3782 4305
rect 3659 3995 3726 4279
rect 3243 3437 3726 3995
rect 3243 3114 3258 3437
rect 3183 3106 3258 3114
rect 2672 3049 3024 3056
rect 2530 2991 3137 2993
rect 2530 2899 3073 2991
rect 2391 2392 2474 2800
rect 3043 2764 3073 2899
rect 3034 2759 3073 2764
rect 3125 2764 3137 2991
rect 3659 2843 3726 3437
rect 3778 2843 3782 4279
rect 3125 2759 3168 2764
rect 3034 2703 3056 2759
rect 3148 2703 3168 2759
rect 3034 2696 3168 2703
rect 2391 2309 2677 2392
rect 2594 2258 2677 2309
rect 2594 1301 2615 2258
rect 2667 1388 2677 2258
rect 3337 2120 3412 2128
rect 2667 1380 3281 1388
rect 2667 1301 3219 1380
rect 2594 1293 3219 1301
rect 3202 882 3219 1293
rect 3271 882 3281 1380
rect 3202 874 3281 882
rect 3337 449 3346 2120
rect 3398 2078 3412 2120
rect 3659 2078 3782 2843
rect 3398 2023 3782 2078
rect 3398 1520 3726 2023
rect 3398 449 3412 1520
rect 3337 441 3412 449
rect 3659 587 3726 1520
rect 3778 587 3782 2023
rect 3851 3926 23793 4322
rect 3851 3874 3875 3926
rect 23791 3874 23793 3926
rect 3851 3478 23793 3874
rect 3851 3426 3877 3478
rect 23791 3426 23793 3478
rect 3851 3030 23793 3426
rect 3851 2978 3873 3030
rect 23791 2978 23793 3030
rect 3851 2649 23793 2978
rect 3851 2066 3867 2649
rect 23791 2066 23793 2649
rect 3851 1670 23793 2066
rect 3851 1618 3871 1670
rect 23791 1618 23793 1670
rect 3851 1222 23793 1618
rect 3851 1170 3871 1222
rect 23791 1170 23793 1222
rect 3851 774 23793 1170
rect 3851 722 3868 774
rect 23783 722 23793 774
rect 3851 707 23793 722
rect 23867 4276 24055 4311
rect 23867 4190 23879 4276
rect 24043 4190 24055 4276
rect 23867 4052 24055 4190
rect 23867 3966 23879 4052
rect 24043 3966 24055 4052
rect 23867 3828 24055 3966
rect 23867 3742 23879 3828
rect 24043 3742 24055 3828
rect 23867 3604 24055 3742
rect 23867 3518 23879 3604
rect 24043 3518 24055 3604
rect 23867 3380 24055 3518
rect 23867 3294 23879 3380
rect 24043 3294 24055 3380
rect 23867 3156 24055 3294
rect 23867 3070 23879 3156
rect 24043 3070 24055 3156
rect 23867 2932 24055 3070
rect 23867 2846 23879 2932
rect 24043 2846 24055 2932
rect 23867 2020 24055 2846
rect 23867 1934 23879 2020
rect 24043 1934 24055 2020
rect 23867 1796 24055 1934
rect 23867 1710 23879 1796
rect 24043 1710 24055 1796
rect 23867 1572 24055 1710
rect 23867 1486 23879 1572
rect 24043 1486 24055 1572
rect 23867 1348 24055 1486
rect 23867 1262 23879 1348
rect 24043 1262 24055 1348
rect 23867 1124 24055 1262
rect 23867 1038 23879 1124
rect 24043 1038 24055 1124
rect 23867 900 24055 1038
rect 23867 814 23879 900
rect 24043 814 24055 900
rect 3659 423 3782 587
rect 23867 676 24055 814
rect 23867 590 23879 676
rect 24043 590 24055 676
rect 23867 423 24055 590
rect 24118 4150 33518 4482
rect 24118 4098 24139 4150
rect 33513 4098 33518 4150
rect 24118 3702 33518 4098
rect 24118 3650 24138 3702
rect 33512 3650 33518 3702
rect 24118 3254 33518 3650
rect 24118 3202 24135 3254
rect 33509 3202 33518 3254
rect 24118 2807 33518 3202
rect 24118 2755 24136 2807
rect 33510 2755 33518 2807
rect 24118 1894 33518 2755
rect 24118 1842 24138 1894
rect 33512 1842 33518 1894
rect 24118 1446 33518 1842
rect 24118 1394 24139 1446
rect 33513 1394 33518 1446
rect 24118 998 33518 1394
rect 24118 946 24135 998
rect 33509 946 33518 998
rect 24118 839 33518 946
rect 24118 550 24456 839
rect 24656 550 33518 839
rect 34619 4387 44020 4396
rect 34619 4322 34630 4387
rect 43996 4322 44020 4387
rect 34619 3939 44020 4322
rect 34619 3874 34632 3939
rect 43998 3874 44020 3939
rect 34619 3491 44020 3874
rect 34619 3426 34632 3491
rect 43998 3426 44020 3491
rect 34619 3043 44020 3426
rect 34619 2978 34631 3043
rect 43997 2978 44020 3043
rect 34619 2650 44020 2978
rect 34619 2066 34627 2650
rect 43993 2131 44020 2650
rect 43994 2066 44020 2131
rect 34619 1683 44020 2066
rect 34619 1618 34633 1683
rect 43999 1618 44020 1683
rect 34619 1235 44020 1618
rect 34619 1170 34643 1235
rect 44009 1170 44020 1235
rect 34619 787 44020 1170
rect 34619 722 34626 787
rect 43992 722 44020 787
rect 34619 700 44020 722
rect 44099 4276 44287 4310
rect 44099 4190 44111 4276
rect 44275 4190 44287 4276
rect 44099 4052 44287 4190
rect 44099 3966 44111 4052
rect 44275 3966 44287 4052
rect 44099 3828 44287 3966
rect 44099 3742 44111 3828
rect 44275 3742 44287 3828
rect 44099 3604 44287 3742
rect 44099 3518 44111 3604
rect 44275 3518 44287 3604
rect 44099 3380 44287 3518
rect 44099 3294 44111 3380
rect 44275 3294 44287 3380
rect 44099 3156 44287 3294
rect 44099 3070 44111 3156
rect 44275 3070 44287 3156
rect 44099 2932 44287 3070
rect 44099 2846 44111 2932
rect 44275 2846 44287 2932
rect 44099 2020 44287 2846
rect 44099 1934 44111 2020
rect 44275 1934 44287 2020
rect 44099 1796 44287 1934
rect 44099 1710 44111 1796
rect 44275 1710 44287 1796
rect 44099 1572 44287 1710
rect 44099 1486 44111 1572
rect 44275 1486 44287 1572
rect 44099 1348 44287 1486
rect 44099 1262 44111 1348
rect 44275 1262 44287 1348
rect 44099 1124 44287 1262
rect 44099 1038 44111 1124
rect 44275 1038 44287 1124
rect 44099 900 44287 1038
rect 44099 814 44111 900
rect 44275 814 44287 900
rect 24118 498 24132 550
rect 33506 498 33518 550
rect 24118 485 24456 498
rect 24656 485 33518 498
rect 24118 483 33518 485
rect 44099 676 44287 814
rect 44099 590 44111 676
rect 44275 590 44287 676
rect 44099 423 44287 590
rect 44360 4150 64267 4482
rect 44360 4098 44385 4150
rect 64231 4098 64267 4150
rect 44360 3702 64267 4098
rect 44360 3650 44389 3702
rect 64235 3650 64267 3702
rect 44360 3254 64267 3650
rect 44360 3202 44391 3254
rect 64237 3202 64267 3254
rect 44360 2806 64267 3202
rect 44360 2754 44386 2806
rect 64232 2754 64267 2806
rect 44360 1894 64267 2754
rect 44360 1842 44384 1894
rect 64230 1842 64267 1894
rect 44360 1446 64267 1842
rect 44360 1394 44385 1446
rect 64231 1394 64267 1446
rect 44360 998 64267 1394
rect 44360 946 44390 998
rect 64236 946 64267 998
rect 44360 550 64267 946
rect 44360 498 44381 550
rect 64227 498 64267 550
rect 44360 483 64267 498
rect 64369 4279 64450 4305
rect 64369 2843 64376 4279
rect 64428 2843 64450 4279
rect 64369 2023 64450 2843
rect 64369 587 64376 2023
rect 64428 587 64450 2023
rect 64369 423 64450 587
rect 1261 303 1462 309
rect 1261 251 1275 303
rect 1449 251 1462 303
rect 3659 300 64450 423
rect 1261 231 1462 251
rect 24450 231 24640 238
rect 1261 227 24640 231
rect 1261 113 24460 227
rect 24630 113 24640 227
rect 1261 108 24640 113
rect 24450 103 24640 108
rect 0 0 212 16
rect 64759 14 64773 12100
rect 64959 14 64971 12100
rect 64759 1 64971 14
<< via2 >>
rect 15 16 201 12102
rect 51536 10774 51731 10998
rect 51556 8168 52428 8364
rect 51556 8116 52428 8168
rect 51556 7720 52428 8116
rect 51556 7668 52428 7720
rect 51556 7464 52428 7668
rect 24456 550 24656 839
rect 24456 498 24656 550
rect 24456 485 24656 498
rect 24460 113 24630 227
rect 64773 14 64959 12100
<< metal3 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 16 212 12102
rect 64759 12100 64971 12118
rect 51535 10998 51732 11008
rect 51535 10774 51536 10998
rect 51731 10774 51732 10998
rect 51535 8385 51732 10774
rect 51535 8364 52452 8385
rect 51535 7464 51556 8364
rect 52428 7464 52452 8364
rect 51535 7435 52452 7464
rect 24456 839 24656 849
rect 24456 238 24656 485
rect 24450 227 24656 238
rect 24450 113 24460 227
rect 24630 113 24656 227
rect 24450 108 24656 113
rect 24450 103 24640 108
rect 0 0 212 16
rect 64759 14 64773 12100
rect 64959 14 64971 12100
rect 64759 1 64971 14
<< via3 >>
rect 15 16 201 12102
rect 64773 14 64959 12100
<< metal4 >>
rect 0 12102 212 12117
rect 0 16 15 12102
rect 201 16 212 12102
rect 0 0 212 16
rect 64759 12100 64971 12118
rect 64759 14 64773 12100
rect 64959 14 64971 12100
rect 64759 1 64971 14
<< labels >>
flabel metal2 51536 11369 51733 12118 0 FreeSans 200 0 0 0 OUT
port 1 nsew signal output
flabel metal2 11536 11369 11734 12117 0 FreeSans 200 0 0 0 D0
port 2 nsew signal input
flabel metal2 10540 11369 10738 12117 0 FreeSans 200 0 0 0 D1
port 3 nsew signal input
flabel metal2 9544 11369 9742 12117 0 FreeSans 200 0 0 0 D2
port 4 nsew signal input
flabel metal2 8548 11369 8746 12117 0 FreeSans 200 0 0 0 D3
port 5 nsew signal input
flabel metal2 7552 11369 7750 12117 0 FreeSans 200 0 0 0 D4
port 6 nsew signal input
flabel metal2 6556 11369 6754 12117 0 FreeSans 200 0 0 0 D5
port 7 nsew signal input
flabel metal2 5560 11369 5758 12117 0 FreeSans 200 0 0 0 D6
port 8 nsew signal input
flabel metal2 4564 11369 4762 12117 0 FreeSans 200 0 0 0 D7
port 9 nsew signal input
flabel metal2 3568 11369 3766 12117 0 FreeSans 200 0 0 0 D8
port 10 nsew signal input
flabel metal2 2572 11369 2770 12117 0 FreeSans 200 0 0 0 D9
port 11 nsew signal input
flabel metal2 1576 11369 1774 12117 0 FreeSans 200 0 0 0 D10
port 12 nsew signal input
flabel metal2 580 11369 778 12117 0 FreeSans 200 0 0 0 D11
port 13 nsew signal input
flabel metal4 64759 1 64971 12118 0 FreeSans 400 0 0 0 VDD
port 14 nsew power bidirectional
flabel metal4 0 0 212 12117 0 FreeSans 400 0 0 0 VSS
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 64971 12118
string MASKHINTS_DUALGATE 0 0 64971 12118
string MASKHINTS_V5_XTOR 0 0 64971 12118
<< end >>
