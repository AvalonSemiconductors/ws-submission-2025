`default_nettype none

module vga_demo(
	input clk,
	input rst_n,
	output [31:0] argb,
	output hsync,
	output vsync
);

wire display_on;
wire [9:0] hpos;
wire [9:0] vpos;

hvsync_generator_t hvsync_generator_t(
	.clk(clk),
	.reset(!rst_n),
	.hsync(hsync),
	.vsync(vsync),
	.display_on(display_on),
	.hpos(hpos),
	.vpos(vpos)
);

reg [9:0] frame;
reg last_frame;
reg dir;
always @(posedge clk) begin
	if(!rst_n) begin
		frame <= 0;
		last_frame <= 0;
		dir <= 0;
	end else begin
		last_frame <= vsync;
		if(vsync && !last_frame) begin
			frame <= frame + 1;
			if(frame[7:0] == 8'hFF) dir <= !dir;
		end
	end
end
  
wire [9:0] distance = vpos + hpos + frame;
  
wire bitmap;
bitmap_source bitmap_source(
	.column(hpos[6:0]),
	.row(vpos[6:0]),
	.pixel(bitmap)
);

wire active_area = display_on & !hpos[9] & (vpos >= 128 || hpos >= 128 || !bitmap);
wire [7:0] inv_frame = 255 - frame[7:0];
wire [15:0] test1 = hpos[8:1] * (dir != 0 ? {8'h00, inv_frame} : {8'h00, frame[7:0]});
assign argb = {8'hFF, test1[15:8], vpos[7:0], distance[8:1]} & {32{active_area}};


endmodule

/*
Video sync generator, used to drive a VGA monitor.
Timing from: https://en.wikipedia.org/wiki/Video_Graphics_Array
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
- From 8bitworkshop.com
*/

module hvsync_generator_t(clk, reset, hsync, vsync, display_on, hpos, vpos);

input clk;
input reset;
output reg hsync, vsync;
output display_on;
output reg [9:0] hpos;
output reg [9:0] vpos;

// declarations for TV-simulator sync parameters
// horizontal constants
parameter H_DISPLAY       = 640; // horizontal display width
parameter H_BACK          =  48; // horizontal left border (back porch)
parameter H_FRONT         =  16; // horizontal right border (front porch)
parameter H_SYNC          =  96; // horizontal sync width
// vertical constants
parameter V_DISPLAY       = 480; // vertical display height
parameter V_TOP           =  33; // vertical top border
parameter V_BOTTOM        =  10; // vertical bottom border
parameter V_SYNC          =   2; // vertical sync # lines
// derived constants
parameter H_SYNC_START    = H_DISPLAY + H_FRONT;
parameter H_SYNC_END      = H_DISPLAY + H_FRONT + H_SYNC - 1;
parameter H_MAX           = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
parameter V_SYNC_START    = V_DISPLAY + V_BOTTOM;
parameter V_SYNC_END      = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
parameter V_MAX           = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

wire hmaxxed = (hpos == H_MAX) || reset;	// set when hpos is maximum
wire vmaxxed = (vpos == V_MAX) || reset;	// set when vpos is maximum
  
// horizontal position counter
always @(posedge clk)
begin
	hsync <= (hpos>=H_SYNC_START && hpos<=H_SYNC_END);
	if(hmaxxed)
		hpos <= 0;
	else
		hpos <= hpos + 1;
end

// vertical position counter
always @(posedge clk)
begin
	vsync <= (vpos>=V_SYNC_START && vpos<=V_SYNC_END);
	if(hmaxxed)
		if (vmaxxed)
			vpos <= 0;
		else
			vpos <= vpos + 1;
end
  
// display_on is set when beam is in "safe" visible frame
assign display_on = (hpos<H_DISPLAY) && (vpos<V_DISPLAY);

endmodule

`default_nettype none

module bitmap_source(
input [6:0] column,
input [6:0] row,
output pixel
);

reg rom;
assign pixel = rom;
always @(*) begin
	case({column, row})
		default: rom = 1'bx;
		0: rom = 1'b0;
		1: rom = 1'b0;
		2: rom = 1'b0;
		3: rom = 1'b0;
		4: rom = 1'b0;
		5: rom = 1'b0;
		6: rom = 1'b0;
		7: rom = 1'b0;
		8: rom = 1'b0;
		9: rom = 1'b0;
		10: rom = 1'b0;
		11: rom = 1'b0;
		12: rom = 1'b0;
		13: rom = 1'b0;
		14: rom = 1'b0;
		15: rom = 1'b0;
		16: rom = 1'b0;
		17: rom = 1'b0;
		18: rom = 1'b0;
		19: rom = 1'b0;
		20: rom = 1'b0;
		21: rom = 1'b0;
		22: rom = 1'b0;
		23: rom = 1'b0;
		24: rom = 1'b0;
		25: rom = 1'b0;
		26: rom = 1'b0;
		27: rom = 1'b0;
		28: rom = 1'b0;
		29: rom = 1'b0;
		30: rom = 1'b0;
		31: rom = 1'b0;
		32: rom = 1'b0;
		33: rom = 1'b0;
		34: rom = 1'b0;
		35: rom = 1'b0;
		36: rom = 1'b0;
		37: rom = 1'b0;
		38: rom = 1'b0;
		39: rom = 1'b0;
		40: rom = 1'b0;
		41: rom = 1'b0;
		42: rom = 1'b0;
		43: rom = 1'b0;
		44: rom = 1'b0;
		45: rom = 1'b0;
		46: rom = 1'b0;
		47: rom = 1'b0;
		48: rom = 1'b0;
		49: rom = 1'b0;
		50: rom = 1'b0;
		51: rom = 1'b0;
		52: rom = 1'b0;
		53: rom = 1'b0;
		54: rom = 1'b0;
		55: rom = 1'b0;
		56: rom = 1'b0;
		57: rom = 1'b0;
		58: rom = 1'b0;
		59: rom = 1'b0;
		60: rom = 1'b0;
		61: rom = 1'b0;
		62: rom = 1'b0;
		63: rom = 1'b0;
		64: rom = 1'b0;
		65: rom = 1'b0;
		66: rom = 1'b0;
		67: rom = 1'b0;
		68: rom = 1'b0;
		69: rom = 1'b0;
		70: rom = 1'b0;
		71: rom = 1'b0;
		72: rom = 1'b0;
		73: rom = 1'b0;
		74: rom = 1'b0;
		75: rom = 1'b0;
		76: rom = 1'b0;
		77: rom = 1'b0;
		78: rom = 1'b0;
		79: rom = 1'b0;
		80: rom = 1'b0;
		81: rom = 1'b0;
		82: rom = 1'b0;
		83: rom = 1'b0;
		84: rom = 1'b0;
		85: rom = 1'b0;
		86: rom = 1'b0;
		87: rom = 1'b0;
		88: rom = 1'b0;
		89: rom = 1'b0;
		90: rom = 1'b0;
		91: rom = 1'b0;
		92: rom = 1'b0;
		93: rom = 1'b0;
		94: rom = 1'b0;
		95: rom = 1'b0;
		96: rom = 1'b0;
		97: rom = 1'b0;
		98: rom = 1'b0;
		99: rom = 1'b0;
		100: rom = 1'b0;
		101: rom = 1'b0;
		102: rom = 1'b0;
		103: rom = 1'b0;
		104: rom = 1'b0;
		105: rom = 1'b0;
		106: rom = 1'b0;
		107: rom = 1'b0;
		108: rom = 1'b0;
		109: rom = 1'b0;
		110: rom = 1'b0;
		111: rom = 1'b0;
		112: rom = 1'b0;
		113: rom = 1'b0;
		114: rom = 1'b0;
		115: rom = 1'b0;
		116: rom = 1'b0;
		117: rom = 1'b0;
		118: rom = 1'b0;
		119: rom = 1'b0;
		120: rom = 1'b0;
		121: rom = 1'b0;
		122: rom = 1'b0;
		123: rom = 1'b0;
		124: rom = 1'b0;
		125: rom = 1'b0;
		126: rom = 1'b0;
		127: rom = 1'b0;
		128: rom = 1'b0;
		129: rom = 1'b0;
		130: rom = 1'b0;
		131: rom = 1'b0;
		132: rom = 1'b0;
		133: rom = 1'b0;
		134: rom = 1'b0;
		135: rom = 1'b0;
		136: rom = 1'b0;
		137: rom = 1'b0;
		138: rom = 1'b0;
		139: rom = 1'b0;
		140: rom = 1'b0;
		141: rom = 1'b0;
		142: rom = 1'b0;
		143: rom = 1'b0;
		144: rom = 1'b0;
		145: rom = 1'b0;
		146: rom = 1'b0;
		147: rom = 1'b0;
		148: rom = 1'b0;
		149: rom = 1'b0;
		150: rom = 1'b0;
		151: rom = 1'b0;
		152: rom = 1'b0;
		153: rom = 1'b0;
		154: rom = 1'b0;
		155: rom = 1'b0;
		156: rom = 1'b0;
		157: rom = 1'b0;
		158: rom = 1'b0;
		159: rom = 1'b0;
		160: rom = 1'b0;
		161: rom = 1'b0;
		162: rom = 1'b0;
		163: rom = 1'b0;
		164: rom = 1'b0;
		165: rom = 1'b0;
		166: rom = 1'b0;
		167: rom = 1'b0;
		168: rom = 1'b0;
		169: rom = 1'b0;
		170: rom = 1'b0;
		171: rom = 1'b0;
		172: rom = 1'b0;
		173: rom = 1'b0;
		174: rom = 1'b0;
		175: rom = 1'b0;
		176: rom = 1'b0;
		177: rom = 1'b0;
		178: rom = 1'b0;
		179: rom = 1'b0;
		180: rom = 1'b0;
		181: rom = 1'b0;
		182: rom = 1'b0;
		183: rom = 1'b0;
		184: rom = 1'b0;
		185: rom = 1'b0;
		186: rom = 1'b0;
		187: rom = 1'b0;
		188: rom = 1'b0;
		189: rom = 1'b0;
		190: rom = 1'b0;
		191: rom = 1'b0;
		192: rom = 1'b0;
		193: rom = 1'b0;
		194: rom = 1'b0;
		195: rom = 1'b0;
		196: rom = 1'b0;
		197: rom = 1'b0;
		198: rom = 1'b0;
		199: rom = 1'b0;
		200: rom = 1'b0;
		201: rom = 1'b0;
		202: rom = 1'b0;
		203: rom = 1'b0;
		204: rom = 1'b0;
		205: rom = 1'b0;
		206: rom = 1'b0;
		207: rom = 1'b0;
		208: rom = 1'b0;
		209: rom = 1'b0;
		210: rom = 1'b0;
		211: rom = 1'b0;
		212: rom = 1'b0;
		213: rom = 1'b0;
		214: rom = 1'b0;
		215: rom = 1'b0;
		216: rom = 1'b0;
		217: rom = 1'b0;
		218: rom = 1'b0;
		219: rom = 1'b0;
		220: rom = 1'b0;
		221: rom = 1'b0;
		222: rom = 1'b0;
		223: rom = 1'b0;
		224: rom = 1'b0;
		225: rom = 1'b0;
		226: rom = 1'b0;
		227: rom = 1'b0;
		228: rom = 1'b0;
		229: rom = 1'b0;
		230: rom = 1'b0;
		231: rom = 1'b0;
		232: rom = 1'b0;
		233: rom = 1'b0;
		234: rom = 1'b0;
		235: rom = 1'b0;
		236: rom = 1'b0;
		237: rom = 1'b0;
		238: rom = 1'b0;
		239: rom = 1'b0;
		240: rom = 1'b0;
		241: rom = 1'b0;
		242: rom = 1'b0;
		243: rom = 1'b0;
		244: rom = 1'b0;
		245: rom = 1'b0;
		246: rom = 1'b0;
		247: rom = 1'b0;
		248: rom = 1'b0;
		249: rom = 1'b0;
		250: rom = 1'b0;
		251: rom = 1'b0;
		252: rom = 1'b0;
		253: rom = 1'b0;
		254: rom = 1'b0;
		255: rom = 1'b0;
		256: rom = 1'b0;
		257: rom = 1'b0;
		258: rom = 1'b0;
		259: rom = 1'b0;
		260: rom = 1'b0;
		261: rom = 1'b0;
		262: rom = 1'b0;
		263: rom = 1'b0;
		264: rom = 1'b0;
		265: rom = 1'b0;
		266: rom = 1'b0;
		267: rom = 1'b0;
		268: rom = 1'b0;
		269: rom = 1'b0;
		270: rom = 1'b0;
		271: rom = 1'b0;
		272: rom = 1'b0;
		273: rom = 1'b0;
		274: rom = 1'b0;
		275: rom = 1'b0;
		276: rom = 1'b0;
		277: rom = 1'b0;
		278: rom = 1'b0;
		279: rom = 1'b0;
		280: rom = 1'b0;
		281: rom = 1'b0;
		282: rom = 1'b0;
		283: rom = 1'b0;
		284: rom = 1'b0;
		285: rom = 1'b0;
		286: rom = 1'b0;
		287: rom = 1'b0;
		288: rom = 1'b0;
		289: rom = 1'b0;
		290: rom = 1'b0;
		291: rom = 1'b0;
		292: rom = 1'b0;
		293: rom = 1'b0;
		294: rom = 1'b0;
		295: rom = 1'b0;
		296: rom = 1'b0;
		297: rom = 1'b0;
		298: rom = 1'b0;
		299: rom = 1'b0;
		300: rom = 1'b0;
		301: rom = 1'b0;
		302: rom = 1'b0;
		303: rom = 1'b0;
		304: rom = 1'b0;
		305: rom = 1'b0;
		306: rom = 1'b0;
		307: rom = 1'b0;
		308: rom = 1'b0;
		309: rom = 1'b0;
		310: rom = 1'b0;
		311: rom = 1'b0;
		312: rom = 1'b0;
		313: rom = 1'b0;
		314: rom = 1'b0;
		315: rom = 1'b0;
		316: rom = 1'b0;
		317: rom = 1'b0;
		318: rom = 1'b0;
		319: rom = 1'b0;
		320: rom = 1'b0;
		321: rom = 1'b0;
		322: rom = 1'b0;
		323: rom = 1'b0;
		324: rom = 1'b0;
		325: rom = 1'b0;
		326: rom = 1'b0;
		327: rom = 1'b0;
		328: rom = 1'b0;
		329: rom = 1'b0;
		330: rom = 1'b0;
		331: rom = 1'b0;
		332: rom = 1'b0;
		333: rom = 1'b0;
		334: rom = 1'b0;
		335: rom = 1'b0;
		336: rom = 1'b0;
		337: rom = 1'b0;
		338: rom = 1'b0;
		339: rom = 1'b0;
		340: rom = 1'b0;
		341: rom = 1'b0;
		342: rom = 1'b0;
		343: rom = 1'b0;
		344: rom = 1'b0;
		345: rom = 1'b0;
		346: rom = 1'b0;
		347: rom = 1'b0;
		348: rom = 1'b0;
		349: rom = 1'b0;
		350: rom = 1'b0;
		351: rom = 1'b0;
		352: rom = 1'b0;
		353: rom = 1'b0;
		354: rom = 1'b0;
		355: rom = 1'b0;
		356: rom = 1'b0;
		357: rom = 1'b0;
		358: rom = 1'b0;
		359: rom = 1'b0;
		360: rom = 1'b0;
		361: rom = 1'b0;
		362: rom = 1'b0;
		363: rom = 1'b0;
		364: rom = 1'b0;
		365: rom = 1'b0;
		366: rom = 1'b0;
		367: rom = 1'b0;
		368: rom = 1'b0;
		369: rom = 1'b0;
		370: rom = 1'b0;
		371: rom = 1'b0;
		372: rom = 1'b0;
		373: rom = 1'b0;
		374: rom = 1'b0;
		375: rom = 1'b0;
		376: rom = 1'b0;
		377: rom = 1'b0;
		378: rom = 1'b0;
		379: rom = 1'b0;
		380: rom = 1'b0;
		381: rom = 1'b0;
		382: rom = 1'b0;
		383: rom = 1'b0;
		384: rom = 1'b0;
		385: rom = 1'b0;
		386: rom = 1'b0;
		387: rom = 1'b0;
		388: rom = 1'b0;
		389: rom = 1'b0;
		390: rom = 1'b0;
		391: rom = 1'b0;
		392: rom = 1'b0;
		393: rom = 1'b0;
		394: rom = 1'b0;
		395: rom = 1'b0;
		396: rom = 1'b0;
		397: rom = 1'b0;
		398: rom = 1'b0;
		399: rom = 1'b0;
		400: rom = 1'b0;
		401: rom = 1'b0;
		402: rom = 1'b0;
		403: rom = 1'b0;
		404: rom = 1'b0;
		405: rom = 1'b0;
		406: rom = 1'b0;
		407: rom = 1'b0;
		408: rom = 1'b0;
		409: rom = 1'b0;
		410: rom = 1'b0;
		411: rom = 1'b0;
		412: rom = 1'b0;
		413: rom = 1'b0;
		414: rom = 1'b0;
		415: rom = 1'b0;
		416: rom = 1'b0;
		417: rom = 1'b0;
		418: rom = 1'b0;
		419: rom = 1'b0;
		420: rom = 1'b0;
		421: rom = 1'b0;
		422: rom = 1'b0;
		423: rom = 1'b0;
		424: rom = 1'b0;
		425: rom = 1'b0;
		426: rom = 1'b0;
		427: rom = 1'b0;
		428: rom = 1'b0;
		429: rom = 1'b0;
		430: rom = 1'b0;
		431: rom = 1'b0;
		432: rom = 1'b0;
		433: rom = 1'b0;
		434: rom = 1'b0;
		435: rom = 1'b0;
		436: rom = 1'b0;
		437: rom = 1'b0;
		438: rom = 1'b0;
		439: rom = 1'b0;
		440: rom = 1'b0;
		441: rom = 1'b0;
		442: rom = 1'b0;
		443: rom = 1'b0;
		444: rom = 1'b0;
		445: rom = 1'b0;
		446: rom = 1'b0;
		447: rom = 1'b0;
		448: rom = 1'b0;
		449: rom = 1'b0;
		450: rom = 1'b0;
		451: rom = 1'b0;
		452: rom = 1'b0;
		453: rom = 1'b0;
		454: rom = 1'b0;
		455: rom = 1'b0;
		456: rom = 1'b0;
		457: rom = 1'b0;
		458: rom = 1'b0;
		459: rom = 1'b0;
		460: rom = 1'b0;
		461: rom = 1'b0;
		462: rom = 1'b0;
		463: rom = 1'b0;
		464: rom = 1'b0;
		465: rom = 1'b0;
		466: rom = 1'b0;
		467: rom = 1'b0;
		468: rom = 1'b0;
		469: rom = 1'b0;
		470: rom = 1'b0;
		471: rom = 1'b0;
		472: rom = 1'b0;
		473: rom = 1'b0;
		474: rom = 1'b0;
		475: rom = 1'b0;
		476: rom = 1'b0;
		477: rom = 1'b0;
		478: rom = 1'b0;
		479: rom = 1'b0;
		480: rom = 1'b0;
		481: rom = 1'b0;
		482: rom = 1'b0;
		483: rom = 1'b0;
		484: rom = 1'b0;
		485: rom = 1'b0;
		486: rom = 1'b0;
		487: rom = 1'b0;
		488: rom = 1'b0;
		489: rom = 1'b0;
		490: rom = 1'b0;
		491: rom = 1'b0;
		492: rom = 1'b0;
		493: rom = 1'b0;
		494: rom = 1'b0;
		495: rom = 1'b0;
		496: rom = 1'b0;
		497: rom = 1'b0;
		498: rom = 1'b0;
		499: rom = 1'b0;
		500: rom = 1'b0;
		501: rom = 1'b0;
		502: rom = 1'b0;
		503: rom = 1'b0;
		504: rom = 1'b0;
		505: rom = 1'b0;
		506: rom = 1'b0;
		507: rom = 1'b0;
		508: rom = 1'b0;
		509: rom = 1'b0;
		510: rom = 1'b0;
		511: rom = 1'b0;
		512: rom = 1'b0;
		513: rom = 1'b0;
		514: rom = 1'b0;
		515: rom = 1'b0;
		516: rom = 1'b0;
		517: rom = 1'b0;
		518: rom = 1'b0;
		519: rom = 1'b0;
		520: rom = 1'b0;
		521: rom = 1'b0;
		522: rom = 1'b0;
		523: rom = 1'b0;
		524: rom = 1'b0;
		525: rom = 1'b0;
		526: rom = 1'b0;
		527: rom = 1'b0;
		528: rom = 1'b0;
		529: rom = 1'b0;
		530: rom = 1'b0;
		531: rom = 1'b0;
		532: rom = 1'b0;
		533: rom = 1'b0;
		534: rom = 1'b0;
		535: rom = 1'b0;
		536: rom = 1'b0;
		537: rom = 1'b0;
		538: rom = 1'b0;
		539: rom = 1'b0;
		540: rom = 1'b0;
		541: rom = 1'b0;
		542: rom = 1'b0;
		543: rom = 1'b0;
		544: rom = 1'b0;
		545: rom = 1'b0;
		546: rom = 1'b0;
		547: rom = 1'b0;
		548: rom = 1'b0;
		549: rom = 1'b0;
		550: rom = 1'b0;
		551: rom = 1'b0;
		552: rom = 1'b0;
		553: rom = 1'b0;
		554: rom = 1'b0;
		555: rom = 1'b0;
		556: rom = 1'b0;
		557: rom = 1'b0;
		558: rom = 1'b0;
		559: rom = 1'b0;
		560: rom = 1'b0;
		561: rom = 1'b0;
		562: rom = 1'b0;
		563: rom = 1'b0;
		564: rom = 1'b0;
		565: rom = 1'b0;
		566: rom = 1'b0;
		567: rom = 1'b0;
		568: rom = 1'b0;
		569: rom = 1'b0;
		570: rom = 1'b0;
		571: rom = 1'b0;
		572: rom = 1'b0;
		573: rom = 1'b0;
		574: rom = 1'b0;
		575: rom = 1'b0;
		576: rom = 1'b1;
		577: rom = 1'b1;
		578: rom = 1'b1;
		579: rom = 1'b1;
		580: rom = 1'b1;
		581: rom = 1'b1;
		582: rom = 1'b1;
		583: rom = 1'b1;
		584: rom = 1'b1;
		585: rom = 1'b1;
		586: rom = 1'b1;
		587: rom = 1'b1;
		588: rom = 1'b1;
		589: rom = 1'b1;
		590: rom = 1'b1;
		591: rom = 1'b1;
		592: rom = 1'b1;
		593: rom = 1'b1;
		594: rom = 1'b0;
		595: rom = 1'b0;
		596: rom = 1'b0;
		597: rom = 1'b0;
		598: rom = 1'b0;
		599: rom = 1'b0;
		600: rom = 1'b0;
		601: rom = 1'b0;
		602: rom = 1'b0;
		603: rom = 1'b0;
		604: rom = 1'b0;
		605: rom = 1'b0;
		606: rom = 1'b0;
		607: rom = 1'b0;
		608: rom = 1'b0;
		609: rom = 1'b0;
		610: rom = 1'b0;
		611: rom = 1'b0;
		612: rom = 1'b0;
		613: rom = 1'b0;
		614: rom = 1'b0;
		615: rom = 1'b0;
		616: rom = 1'b0;
		617: rom = 1'b0;
		618: rom = 1'b0;
		619: rom = 1'b0;
		620: rom = 1'b0;
		621: rom = 1'b0;
		622: rom = 1'b0;
		623: rom = 1'b0;
		624: rom = 1'b0;
		625: rom = 1'b0;
		626: rom = 1'b0;
		627: rom = 1'b0;
		628: rom = 1'b0;
		629: rom = 1'b0;
		630: rom = 1'b0;
		631: rom = 1'b0;
		632: rom = 1'b0;
		633: rom = 1'b0;
		634: rom = 1'b0;
		635: rom = 1'b0;
		636: rom = 1'b0;
		637: rom = 1'b0;
		638: rom = 1'b0;
		639: rom = 1'b0;
		640: rom = 1'b0;
		641: rom = 1'b0;
		642: rom = 1'b0;
		643: rom = 1'b0;
		644: rom = 1'b0;
		645: rom = 1'b0;
		646: rom = 1'b0;
		647: rom = 1'b0;
		648: rom = 1'b0;
		649: rom = 1'b0;
		650: rom = 1'b0;
		651: rom = 1'b0;
		652: rom = 1'b0;
		653: rom = 1'b0;
		654: rom = 1'b0;
		655: rom = 1'b0;
		656: rom = 1'b0;
		657: rom = 1'b0;
		658: rom = 1'b0;
		659: rom = 1'b0;
		660: rom = 1'b0;
		661: rom = 1'b0;
		662: rom = 1'b0;
		663: rom = 1'b0;
		664: rom = 1'b0;
		665: rom = 1'b0;
		666: rom = 1'b0;
		667: rom = 1'b0;
		668: rom = 1'b0;
		669: rom = 1'b0;
		670: rom = 1'b0;
		671: rom = 1'b0;
		672: rom = 1'b0;
		673: rom = 1'b0;
		674: rom = 1'b0;
		675: rom = 1'b0;
		676: rom = 1'b0;
		677: rom = 1'b0;
		678: rom = 1'b0;
		679: rom = 1'b0;
		680: rom = 1'b0;
		681: rom = 1'b0;
		682: rom = 1'b0;
		683: rom = 1'b0;
		684: rom = 1'b0;
		685: rom = 1'b0;
		686: rom = 1'b0;
		687: rom = 1'b0;
		688: rom = 1'b0;
		689: rom = 1'b0;
		690: rom = 1'b0;
		691: rom = 1'b0;
		692: rom = 1'b0;
		693: rom = 1'b0;
		694: rom = 1'b0;
		695: rom = 1'b0;
		696: rom = 1'b0;
		697: rom = 1'b0;
		698: rom = 1'b0;
		699: rom = 1'b0;
		700: rom = 1'b1;
		701: rom = 1'b1;
		702: rom = 1'b1;
		703: rom = 1'b1;
		704: rom = 1'b1;
		705: rom = 1'b1;
		706: rom = 1'b1;
		707: rom = 1'b1;
		708: rom = 1'b1;
		709: rom = 1'b1;
		710: rom = 1'b1;
		711: rom = 1'b1;
		712: rom = 1'b1;
		713: rom = 1'b1;
		714: rom = 1'b1;
		715: rom = 1'b1;
		716: rom = 1'b1;
		717: rom = 1'b1;
		718: rom = 1'b1;
		719: rom = 1'b1;
		720: rom = 1'b1;
		721: rom = 1'b1;
		722: rom = 1'b0;
		723: rom = 1'b0;
		724: rom = 1'b0;
		725: rom = 1'b0;
		726: rom = 1'b0;
		727: rom = 1'b0;
		728: rom = 1'b0;
		729: rom = 1'b0;
		730: rom = 1'b0;
		731: rom = 1'b0;
		732: rom = 1'b0;
		733: rom = 1'b0;
		734: rom = 1'b0;
		735: rom = 1'b0;
		736: rom = 1'b0;
		737: rom = 1'b0;
		738: rom = 1'b0;
		739: rom = 1'b0;
		740: rom = 1'b0;
		741: rom = 1'b0;
		742: rom = 1'b0;
		743: rom = 1'b0;
		744: rom = 1'b0;
		745: rom = 1'b0;
		746: rom = 1'b0;
		747: rom = 1'b0;
		748: rom = 1'b0;
		749: rom = 1'b0;
		750: rom = 1'b0;
		751: rom = 1'b0;
		752: rom = 1'b0;
		753: rom = 1'b0;
		754: rom = 1'b0;
		755: rom = 1'b0;
		756: rom = 1'b0;
		757: rom = 1'b0;
		758: rom = 1'b0;
		759: rom = 1'b0;
		760: rom = 1'b0;
		761: rom = 1'b0;
		762: rom = 1'b0;
		763: rom = 1'b0;
		764: rom = 1'b0;
		765: rom = 1'b0;
		766: rom = 1'b0;
		767: rom = 1'b0;
		768: rom = 1'b0;
		769: rom = 1'b0;
		770: rom = 1'b0;
		771: rom = 1'b0;
		772: rom = 1'b0;
		773: rom = 1'b0;
		774: rom = 1'b0;
		775: rom = 1'b0;
		776: rom = 1'b0;
		777: rom = 1'b0;
		778: rom = 1'b0;
		779: rom = 1'b0;
		780: rom = 1'b0;
		781: rom = 1'b0;
		782: rom = 1'b0;
		783: rom = 1'b0;
		784: rom = 1'b0;
		785: rom = 1'b0;
		786: rom = 1'b0;
		787: rom = 1'b0;
		788: rom = 1'b0;
		789: rom = 1'b0;
		790: rom = 1'b0;
		791: rom = 1'b0;
		792: rom = 1'b0;
		793: rom = 1'b0;
		794: rom = 1'b0;
		795: rom = 1'b0;
		796: rom = 1'b0;
		797: rom = 1'b0;
		798: rom = 1'b0;
		799: rom = 1'b0;
		800: rom = 1'b0;
		801: rom = 1'b0;
		802: rom = 1'b0;
		803: rom = 1'b0;
		804: rom = 1'b0;
		805: rom = 1'b0;
		806: rom = 1'b0;
		807: rom = 1'b0;
		808: rom = 1'b0;
		809: rom = 1'b0;
		810: rom = 1'b0;
		811: rom = 1'b0;
		812: rom = 1'b0;
		813: rom = 1'b0;
		814: rom = 1'b0;
		815: rom = 1'b0;
		816: rom = 1'b0;
		817: rom = 1'b0;
		818: rom = 1'b0;
		819: rom = 1'b0;
		820: rom = 1'b0;
		821: rom = 1'b0;
		822: rom = 1'b0;
		823: rom = 1'b0;
		824: rom = 1'b0;
		825: rom = 1'b1;
		826: rom = 1'b1;
		827: rom = 1'b1;
		828: rom = 1'b1;
		829: rom = 1'b1;
		830: rom = 1'b1;
		831: rom = 1'b1;
		832: rom = 1'b1;
		833: rom = 1'b1;
		834: rom = 1'b1;
		835: rom = 1'b1;
		836: rom = 1'b1;
		837: rom = 1'b1;
		838: rom = 1'b1;
		839: rom = 1'b1;
		840: rom = 1'b1;
		841: rom = 1'b1;
		842: rom = 1'b1;
		843: rom = 1'b1;
		844: rom = 1'b1;
		845: rom = 1'b1;
		846: rom = 1'b1;
		847: rom = 1'b0;
		848: rom = 1'b0;
		849: rom = 1'b0;
		850: rom = 1'b0;
		851: rom = 1'b0;
		852: rom = 1'b0;
		853: rom = 1'b0;
		854: rom = 1'b0;
		855: rom = 1'b0;
		856: rom = 1'b0;
		857: rom = 1'b0;
		858: rom = 1'b0;
		859: rom = 1'b0;
		860: rom = 1'b0;
		861: rom = 1'b0;
		862: rom = 1'b0;
		863: rom = 1'b0;
		864: rom = 1'b0;
		865: rom = 1'b0;
		866: rom = 1'b0;
		867: rom = 1'b0;
		868: rom = 1'b0;
		869: rom = 1'b0;
		870: rom = 1'b0;
		871: rom = 1'b0;
		872: rom = 1'b0;
		873: rom = 1'b0;
		874: rom = 1'b0;
		875: rom = 1'b0;
		876: rom = 1'b0;
		877: rom = 1'b0;
		878: rom = 1'b0;
		879: rom = 1'b0;
		880: rom = 1'b0;
		881: rom = 1'b0;
		882: rom = 1'b0;
		883: rom = 1'b0;
		884: rom = 1'b0;
		885: rom = 1'b0;
		886: rom = 1'b0;
		887: rom = 1'b0;
		888: rom = 1'b0;
		889: rom = 1'b0;
		890: rom = 1'b0;
		891: rom = 1'b0;
		892: rom = 1'b0;
		893: rom = 1'b0;
		894: rom = 1'b0;
		895: rom = 1'b0;
		896: rom = 1'b0;
		897: rom = 1'b0;
		898: rom = 1'b0;
		899: rom = 1'b0;
		900: rom = 1'b0;
		901: rom = 1'b0;
		902: rom = 1'b0;
		903: rom = 1'b0;
		904: rom = 1'b0;
		905: rom = 1'b0;
		906: rom = 1'b0;
		907: rom = 1'b0;
		908: rom = 1'b0;
		909: rom = 1'b0;
		910: rom = 1'b0;
		911: rom = 1'b0;
		912: rom = 1'b0;
		913: rom = 1'b0;
		914: rom = 1'b0;
		915: rom = 1'b0;
		916: rom = 1'b0;
		917: rom = 1'b0;
		918: rom = 1'b0;
		919: rom = 1'b0;
		920: rom = 1'b0;
		921: rom = 1'b0;
		922: rom = 1'b0;
		923: rom = 1'b0;
		924: rom = 1'b0;
		925: rom = 1'b0;
		926: rom = 1'b0;
		927: rom = 1'b0;
		928: rom = 1'b0;
		929: rom = 1'b0;
		930: rom = 1'b0;
		931: rom = 1'b0;
		932: rom = 1'b0;
		933: rom = 1'b0;
		934: rom = 1'b0;
		935: rom = 1'b0;
		936: rom = 1'b0;
		937: rom = 1'b0;
		938: rom = 1'b0;
		939: rom = 1'b0;
		940: rom = 1'b0;
		941: rom = 1'b0;
		942: rom = 1'b0;
		943: rom = 1'b0;
		944: rom = 1'b0;
		945: rom = 1'b0;
		946: rom = 1'b0;
		947: rom = 1'b0;
		948: rom = 1'b0;
		949: rom = 1'b0;
		950: rom = 1'b0;
		951: rom = 1'b1;
		952: rom = 1'b1;
		953: rom = 1'b1;
		954: rom = 1'b1;
		955: rom = 1'b1;
		956: rom = 1'b1;
		957: rom = 1'b1;
		958: rom = 1'b1;
		959: rom = 1'b1;
		960: rom = 1'b1;
		961: rom = 1'b1;
		962: rom = 1'b1;
		963: rom = 1'b1;
		964: rom = 1'b1;
		965: rom = 1'b1;
		966: rom = 1'b1;
		967: rom = 1'b1;
		968: rom = 1'b1;
		969: rom = 1'b1;
		970: rom = 1'b1;
		971: rom = 1'b1;
		972: rom = 1'b1;
		973: rom = 1'b0;
		974: rom = 1'b0;
		975: rom = 1'b0;
		976: rom = 1'b0;
		977: rom = 1'b0;
		978: rom = 1'b0;
		979: rom = 1'b0;
		980: rom = 1'b0;
		981: rom = 1'b0;
		982: rom = 1'b0;
		983: rom = 1'b0;
		984: rom = 1'b0;
		985: rom = 1'b0;
		986: rom = 1'b0;
		987: rom = 1'b0;
		988: rom = 1'b0;
		989: rom = 1'b0;
		990: rom = 1'b0;
		991: rom = 1'b0;
		992: rom = 1'b0;
		993: rom = 1'b0;
		994: rom = 1'b0;
		995: rom = 1'b0;
		996: rom = 1'b0;
		997: rom = 1'b0;
		998: rom = 1'b0;
		999: rom = 1'b0;
		1000: rom = 1'b0;
		1001: rom = 1'b0;
		1002: rom = 1'b0;
		1003: rom = 1'b0;
		1004: rom = 1'b0;
		1005: rom = 1'b0;
		1006: rom = 1'b0;
		1007: rom = 1'b0;
		1008: rom = 1'b0;
		1009: rom = 1'b0;
		1010: rom = 1'b0;
		1011: rom = 1'b0;
		1012: rom = 1'b0;
		1013: rom = 1'b0;
		1014: rom = 1'b0;
		1015: rom = 1'b0;
		1016: rom = 1'b0;
		1017: rom = 1'b0;
		1018: rom = 1'b0;
		1019: rom = 1'b0;
		1020: rom = 1'b0;
		1021: rom = 1'b0;
		1022: rom = 1'b0;
		1023: rom = 1'b0;
		1024: rom = 1'b0;
		1025: rom = 1'b0;
		1026: rom = 1'b0;
		1027: rom = 1'b0;
		1028: rom = 1'b0;
		1029: rom = 1'b0;
		1030: rom = 1'b0;
		1031: rom = 1'b0;
		1032: rom = 1'b0;
		1033: rom = 1'b0;
		1034: rom = 1'b0;
		1035: rom = 1'b0;
		1036: rom = 1'b0;
		1037: rom = 1'b0;
		1038: rom = 1'b0;
		1039: rom = 1'b0;
		1040: rom = 1'b0;
		1041: rom = 1'b0;
		1042: rom = 1'b0;
		1043: rom = 1'b0;
		1044: rom = 1'b0;
		1045: rom = 1'b0;
		1046: rom = 1'b0;
		1047: rom = 1'b0;
		1048: rom = 1'b0;
		1049: rom = 1'b0;
		1050: rom = 1'b0;
		1051: rom = 1'b0;
		1052: rom = 1'b0;
		1053: rom = 1'b0;
		1054: rom = 1'b0;
		1055: rom = 1'b0;
		1056: rom = 1'b0;
		1057: rom = 1'b0;
		1058: rom = 1'b0;
		1059: rom = 1'b0;
		1060: rom = 1'b0;
		1061: rom = 1'b0;
		1062: rom = 1'b0;
		1063: rom = 1'b0;
		1064: rom = 1'b0;
		1065: rom = 1'b0;
		1066: rom = 1'b0;
		1067: rom = 1'b0;
		1068: rom = 1'b0;
		1069: rom = 1'b0;
		1070: rom = 1'b0;
		1071: rom = 1'b0;
		1072: rom = 1'b0;
		1073: rom = 1'b0;
		1074: rom = 1'b0;
		1075: rom = 1'b0;
		1076: rom = 1'b0;
		1077: rom = 1'b1;
		1078: rom = 1'b1;
		1079: rom = 1'b1;
		1080: rom = 1'b1;
		1081: rom = 1'b1;
		1082: rom = 1'b1;
		1083: rom = 1'b1;
		1084: rom = 1'b1;
		1085: rom = 1'b1;
		1086: rom = 1'b1;
		1087: rom = 1'b1;
		1088: rom = 1'b1;
		1089: rom = 1'b1;
		1090: rom = 1'b1;
		1091: rom = 1'b1;
		1092: rom = 1'b1;
		1093: rom = 1'b1;
		1094: rom = 1'b1;
		1095: rom = 1'b1;
		1096: rom = 1'b1;
		1097: rom = 1'b1;
		1098: rom = 1'b1;
		1099: rom = 1'b0;
		1100: rom = 1'b0;
		1101: rom = 1'b0;
		1102: rom = 1'b0;
		1103: rom = 1'b0;
		1104: rom = 1'b0;
		1105: rom = 1'b0;
		1106: rom = 1'b0;
		1107: rom = 1'b0;
		1108: rom = 1'b0;
		1109: rom = 1'b0;
		1110: rom = 1'b0;
		1111: rom = 1'b0;
		1112: rom = 1'b0;
		1113: rom = 1'b0;
		1114: rom = 1'b0;
		1115: rom = 1'b0;
		1116: rom = 1'b0;
		1117: rom = 1'b0;
		1118: rom = 1'b0;
		1119: rom = 1'b0;
		1120: rom = 1'b0;
		1121: rom = 1'b0;
		1122: rom = 1'b0;
		1123: rom = 1'b0;
		1124: rom = 1'b0;
		1125: rom = 1'b0;
		1126: rom = 1'b0;
		1127: rom = 1'b0;
		1128: rom = 1'b0;
		1129: rom = 1'b0;
		1130: rom = 1'b0;
		1131: rom = 1'b0;
		1132: rom = 1'b0;
		1133: rom = 1'b0;
		1134: rom = 1'b0;
		1135: rom = 1'b0;
		1136: rom = 1'b0;
		1137: rom = 1'b0;
		1138: rom = 1'b0;
		1139: rom = 1'b0;
		1140: rom = 1'b0;
		1141: rom = 1'b0;
		1142: rom = 1'b0;
		1143: rom = 1'b0;
		1144: rom = 1'b0;
		1145: rom = 1'b0;
		1146: rom = 1'b0;
		1147: rom = 1'b0;
		1148: rom = 1'b0;
		1149: rom = 1'b0;
		1150: rom = 1'b0;
		1151: rom = 1'b0;
		1152: rom = 1'b0;
		1153: rom = 1'b0;
		1154: rom = 1'b0;
		1155: rom = 1'b0;
		1156: rom = 1'b0;
		1157: rom = 1'b0;
		1158: rom = 1'b0;
		1159: rom = 1'b0;
		1160: rom = 1'b0;
		1161: rom = 1'b0;
		1162: rom = 1'b0;
		1163: rom = 1'b0;
		1164: rom = 1'b0;
		1165: rom = 1'b0;
		1166: rom = 1'b0;
		1167: rom = 1'b0;
		1168: rom = 1'b0;
		1169: rom = 1'b0;
		1170: rom = 1'b0;
		1171: rom = 1'b0;
		1172: rom = 1'b0;
		1173: rom = 1'b0;
		1174: rom = 1'b0;
		1175: rom = 1'b0;
		1176: rom = 1'b0;
		1177: rom = 1'b0;
		1178: rom = 1'b0;
		1179: rom = 1'b0;
		1180: rom = 1'b0;
		1181: rom = 1'b0;
		1182: rom = 1'b0;
		1183: rom = 1'b0;
		1184: rom = 1'b0;
		1185: rom = 1'b0;
		1186: rom = 1'b0;
		1187: rom = 1'b0;
		1188: rom = 1'b0;
		1189: rom = 1'b0;
		1190: rom = 1'b0;
		1191: rom = 1'b0;
		1192: rom = 1'b0;
		1193: rom = 1'b0;
		1194: rom = 1'b0;
		1195: rom = 1'b0;
		1196: rom = 1'b0;
		1197: rom = 1'b0;
		1198: rom = 1'b0;
		1199: rom = 1'b0;
		1200: rom = 1'b0;
		1201: rom = 1'b0;
		1202: rom = 1'b0;
		1203: rom = 1'b1;
		1204: rom = 1'b1;
		1205: rom = 1'b1;
		1206: rom = 1'b1;
		1207: rom = 1'b1;
		1208: rom = 1'b1;
		1209: rom = 1'b1;
		1210: rom = 1'b1;
		1211: rom = 1'b1;
		1212: rom = 1'b1;
		1213: rom = 1'b1;
		1214: rom = 1'b1;
		1215: rom = 1'b1;
		1216: rom = 1'b1;
		1217: rom = 1'b1;
		1218: rom = 1'b1;
		1219: rom = 1'b1;
		1220: rom = 1'b1;
		1221: rom = 1'b1;
		1222: rom = 1'b1;
		1223: rom = 1'b1;
		1224: rom = 1'b1;
		1225: rom = 1'b0;
		1226: rom = 1'b0;
		1227: rom = 1'b0;
		1228: rom = 1'b0;
		1229: rom = 1'b0;
		1230: rom = 1'b0;
		1231: rom = 1'b0;
		1232: rom = 1'b0;
		1233: rom = 1'b0;
		1234: rom = 1'b0;
		1235: rom = 1'b0;
		1236: rom = 1'b0;
		1237: rom = 1'b0;
		1238: rom = 1'b0;
		1239: rom = 1'b0;
		1240: rom = 1'b0;
		1241: rom = 1'b0;
		1242: rom = 1'b0;
		1243: rom = 1'b0;
		1244: rom = 1'b0;
		1245: rom = 1'b1;
		1246: rom = 1'b1;
		1247: rom = 1'b0;
		1248: rom = 1'b0;
		1249: rom = 1'b0;
		1250: rom = 1'b0;
		1251: rom = 1'b0;
		1252: rom = 1'b0;
		1253: rom = 1'b0;
		1254: rom = 1'b0;
		1255: rom = 1'b0;
		1256: rom = 1'b0;
		1257: rom = 1'b0;
		1258: rom = 1'b0;
		1259: rom = 1'b0;
		1260: rom = 1'b0;
		1261: rom = 1'b0;
		1262: rom = 1'b0;
		1263: rom = 1'b0;
		1264: rom = 1'b0;
		1265: rom = 1'b0;
		1266: rom = 1'b0;
		1267: rom = 1'b0;
		1268: rom = 1'b0;
		1269: rom = 1'b0;
		1270: rom = 1'b0;
		1271: rom = 1'b0;
		1272: rom = 1'b0;
		1273: rom = 1'b0;
		1274: rom = 1'b0;
		1275: rom = 1'b0;
		1276: rom = 1'b0;
		1277: rom = 1'b0;
		1278: rom = 1'b0;
		1279: rom = 1'b0;
		1280: rom = 1'b0;
		1281: rom = 1'b0;
		1282: rom = 1'b0;
		1283: rom = 1'b0;
		1284: rom = 1'b0;
		1285: rom = 1'b0;
		1286: rom = 1'b0;
		1287: rom = 1'b0;
		1288: rom = 1'b0;
		1289: rom = 1'b0;
		1290: rom = 1'b0;
		1291: rom = 1'b0;
		1292: rom = 1'b0;
		1293: rom = 1'b0;
		1294: rom = 1'b0;
		1295: rom = 1'b0;
		1296: rom = 1'b0;
		1297: rom = 1'b0;
		1298: rom = 1'b0;
		1299: rom = 1'b0;
		1300: rom = 1'b0;
		1301: rom = 1'b0;
		1302: rom = 1'b0;
		1303: rom = 1'b0;
		1304: rom = 1'b0;
		1305: rom = 1'b0;
		1306: rom = 1'b0;
		1307: rom = 1'b0;
		1308: rom = 1'b0;
		1309: rom = 1'b0;
		1310: rom = 1'b0;
		1311: rom = 1'b0;
		1312: rom = 1'b0;
		1313: rom = 1'b0;
		1314: rom = 1'b0;
		1315: rom = 1'b0;
		1316: rom = 1'b0;
		1317: rom = 1'b0;
		1318: rom = 1'b0;
		1319: rom = 1'b0;
		1320: rom = 1'b0;
		1321: rom = 1'b0;
		1322: rom = 1'b0;
		1323: rom = 1'b0;
		1324: rom = 1'b0;
		1325: rom = 1'b0;
		1326: rom = 1'b0;
		1327: rom = 1'b0;
		1328: rom = 1'b0;
		1329: rom = 1'b1;
		1330: rom = 1'b1;
		1331: rom = 1'b1;
		1332: rom = 1'b1;
		1333: rom = 1'b1;
		1334: rom = 1'b1;
		1335: rom = 1'b1;
		1336: rom = 1'b1;
		1337: rom = 1'b1;
		1338: rom = 1'b1;
		1339: rom = 1'b1;
		1340: rom = 1'b1;
		1341: rom = 1'b1;
		1342: rom = 1'b1;
		1343: rom = 1'b1;
		1344: rom = 1'b1;
		1345: rom = 1'b1;
		1346: rom = 1'b1;
		1347: rom = 1'b1;
		1348: rom = 1'b1;
		1349: rom = 1'b1;
		1350: rom = 1'b1;
		1351: rom = 1'b0;
		1352: rom = 1'b0;
		1353: rom = 1'b0;
		1354: rom = 1'b0;
		1355: rom = 1'b0;
		1356: rom = 1'b0;
		1357: rom = 1'b0;
		1358: rom = 1'b0;
		1359: rom = 1'b0;
		1360: rom = 1'b0;
		1361: rom = 1'b0;
		1362: rom = 1'b0;
		1363: rom = 1'b0;
		1364: rom = 1'b0;
		1365: rom = 1'b0;
		1366: rom = 1'b0;
		1367: rom = 1'b0;
		1368: rom = 1'b0;
		1369: rom = 1'b0;
		1370: rom = 1'b1;
		1371: rom = 1'b1;
		1372: rom = 1'b1;
		1373: rom = 1'b1;
		1374: rom = 1'b1;
		1375: rom = 1'b1;
		1376: rom = 1'b1;
		1377: rom = 1'b0;
		1378: rom = 1'b0;
		1379: rom = 1'b0;
		1380: rom = 1'b0;
		1381: rom = 1'b0;
		1382: rom = 1'b0;
		1383: rom = 1'b0;
		1384: rom = 1'b0;
		1385: rom = 1'b0;
		1386: rom = 1'b0;
		1387: rom = 1'b0;
		1388: rom = 1'b0;
		1389: rom = 1'b0;
		1390: rom = 1'b0;
		1391: rom = 1'b0;
		1392: rom = 1'b0;
		1393: rom = 1'b0;
		1394: rom = 1'b0;
		1395: rom = 1'b0;
		1396: rom = 1'b0;
		1397: rom = 1'b0;
		1398: rom = 1'b0;
		1399: rom = 1'b0;
		1400: rom = 1'b0;
		1401: rom = 1'b0;
		1402: rom = 1'b0;
		1403: rom = 1'b0;
		1404: rom = 1'b0;
		1405: rom = 1'b0;
		1406: rom = 1'b0;
		1407: rom = 1'b0;
		1408: rom = 1'b0;
		1409: rom = 1'b0;
		1410: rom = 1'b0;
		1411: rom = 1'b0;
		1412: rom = 1'b0;
		1413: rom = 1'b0;
		1414: rom = 1'b0;
		1415: rom = 1'b0;
		1416: rom = 1'b0;
		1417: rom = 1'b0;
		1418: rom = 1'b0;
		1419: rom = 1'b0;
		1420: rom = 1'b0;
		1421: rom = 1'b0;
		1422: rom = 1'b0;
		1423: rom = 1'b0;
		1424: rom = 1'b0;
		1425: rom = 1'b0;
		1426: rom = 1'b0;
		1427: rom = 1'b0;
		1428: rom = 1'b0;
		1429: rom = 1'b0;
		1430: rom = 1'b0;
		1431: rom = 1'b0;
		1432: rom = 1'b0;
		1433: rom = 1'b0;
		1434: rom = 1'b0;
		1435: rom = 1'b0;
		1436: rom = 1'b0;
		1437: rom = 1'b0;
		1438: rom = 1'b0;
		1439: rom = 1'b0;
		1440: rom = 1'b0;
		1441: rom = 1'b0;
		1442: rom = 1'b0;
		1443: rom = 1'b0;
		1444: rom = 1'b0;
		1445: rom = 1'b0;
		1446: rom = 1'b0;
		1447: rom = 1'b0;
		1448: rom = 1'b0;
		1449: rom = 1'b0;
		1450: rom = 1'b0;
		1451: rom = 1'b0;
		1452: rom = 1'b0;
		1453: rom = 1'b0;
		1454: rom = 1'b0;
		1455: rom = 1'b0;
		1456: rom = 1'b1;
		1457: rom = 1'b1;
		1458: rom = 1'b1;
		1459: rom = 1'b1;
		1460: rom = 1'b1;
		1461: rom = 1'b1;
		1462: rom = 1'b1;
		1463: rom = 1'b1;
		1464: rom = 1'b1;
		1465: rom = 1'b1;
		1466: rom = 1'b1;
		1467: rom = 1'b1;
		1468: rom = 1'b1;
		1469: rom = 1'b1;
		1470: rom = 1'b1;
		1471: rom = 1'b1;
		1472: rom = 1'b1;
		1473: rom = 1'b1;
		1474: rom = 1'b1;
		1475: rom = 1'b1;
		1476: rom = 1'b1;
		1477: rom = 1'b0;
		1478: rom = 1'b0;
		1479: rom = 1'b0;
		1480: rom = 1'b0;
		1481: rom = 1'b0;
		1482: rom = 1'b0;
		1483: rom = 1'b0;
		1484: rom = 1'b0;
		1485: rom = 1'b0;
		1486: rom = 1'b0;
		1487: rom = 1'b0;
		1488: rom = 1'b0;
		1489: rom = 1'b0;
		1490: rom = 1'b0;
		1491: rom = 1'b0;
		1492: rom = 1'b0;
		1493: rom = 1'b0;
		1494: rom = 1'b0;
		1495: rom = 1'b1;
		1496: rom = 1'b1;
		1497: rom = 1'b1;
		1498: rom = 1'b1;
		1499: rom = 1'b1;
		1500: rom = 1'b1;
		1501: rom = 1'b1;
		1502: rom = 1'b1;
		1503: rom = 1'b1;
		1504: rom = 1'b1;
		1505: rom = 1'b1;
		1506: rom = 1'b1;
		1507: rom = 1'b0;
		1508: rom = 1'b0;
		1509: rom = 1'b0;
		1510: rom = 1'b0;
		1511: rom = 1'b0;
		1512: rom = 1'b0;
		1513: rom = 1'b0;
		1514: rom = 1'b0;
		1515: rom = 1'b0;
		1516: rom = 1'b0;
		1517: rom = 1'b0;
		1518: rom = 1'b0;
		1519: rom = 1'b0;
		1520: rom = 1'b0;
		1521: rom = 1'b0;
		1522: rom = 1'b0;
		1523: rom = 1'b0;
		1524: rom = 1'b0;
		1525: rom = 1'b0;
		1526: rom = 1'b0;
		1527: rom = 1'b0;
		1528: rom = 1'b0;
		1529: rom = 1'b0;
		1530: rom = 1'b0;
		1531: rom = 1'b0;
		1532: rom = 1'b0;
		1533: rom = 1'b0;
		1534: rom = 1'b0;
		1535: rom = 1'b0;
		1536: rom = 1'b0;
		1537: rom = 1'b0;
		1538: rom = 1'b0;
		1539: rom = 1'b0;
		1540: rom = 1'b0;
		1541: rom = 1'b0;
		1542: rom = 1'b0;
		1543: rom = 1'b0;
		1544: rom = 1'b0;
		1545: rom = 1'b0;
		1546: rom = 1'b0;
		1547: rom = 1'b0;
		1548: rom = 1'b0;
		1549: rom = 1'b0;
		1550: rom = 1'b0;
		1551: rom = 1'b0;
		1552: rom = 1'b0;
		1553: rom = 1'b0;
		1554: rom = 1'b0;
		1555: rom = 1'b0;
		1556: rom = 1'b0;
		1557: rom = 1'b0;
		1558: rom = 1'b0;
		1559: rom = 1'b0;
		1560: rom = 1'b0;
		1561: rom = 1'b0;
		1562: rom = 1'b0;
		1563: rom = 1'b0;
		1564: rom = 1'b0;
		1565: rom = 1'b0;
		1566: rom = 1'b0;
		1567: rom = 1'b0;
		1568: rom = 1'b0;
		1569: rom = 1'b0;
		1570: rom = 1'b0;
		1571: rom = 1'b0;
		1572: rom = 1'b0;
		1573: rom = 1'b0;
		1574: rom = 1'b0;
		1575: rom = 1'b0;
		1576: rom = 1'b0;
		1577: rom = 1'b0;
		1578: rom = 1'b0;
		1579: rom = 1'b0;
		1580: rom = 1'b0;
		1581: rom = 1'b0;
		1582: rom = 1'b1;
		1583: rom = 1'b1;
		1584: rom = 1'b1;
		1585: rom = 1'b1;
		1586: rom = 1'b1;
		1587: rom = 1'b1;
		1588: rom = 1'b1;
		1589: rom = 1'b1;
		1590: rom = 1'b1;
		1591: rom = 1'b1;
		1592: rom = 1'b1;
		1593: rom = 1'b1;
		1594: rom = 1'b1;
		1595: rom = 1'b1;
		1596: rom = 1'b1;
		1597: rom = 1'b1;
		1598: rom = 1'b1;
		1599: rom = 1'b1;
		1600: rom = 1'b1;
		1601: rom = 1'b1;
		1602: rom = 1'b1;
		1603: rom = 1'b0;
		1604: rom = 1'b0;
		1605: rom = 1'b0;
		1606: rom = 1'b0;
		1607: rom = 1'b0;
		1608: rom = 1'b0;
		1609: rom = 1'b0;
		1610: rom = 1'b0;
		1611: rom = 1'b0;
		1612: rom = 1'b0;
		1613: rom = 1'b0;
		1614: rom = 1'b0;
		1615: rom = 1'b0;
		1616: rom = 1'b0;
		1617: rom = 1'b0;
		1618: rom = 1'b0;
		1619: rom = 1'b0;
		1620: rom = 1'b0;
		1621: rom = 1'b1;
		1622: rom = 1'b1;
		1623: rom = 1'b1;
		1624: rom = 1'b1;
		1625: rom = 1'b1;
		1626: rom = 1'b1;
		1627: rom = 1'b1;
		1628: rom = 1'b1;
		1629: rom = 1'b1;
		1630: rom = 1'b1;
		1631: rom = 1'b1;
		1632: rom = 1'b1;
		1633: rom = 1'b1;
		1634: rom = 1'b1;
		1635: rom = 1'b1;
		1636: rom = 1'b0;
		1637: rom = 1'b0;
		1638: rom = 1'b0;
		1639: rom = 1'b0;
		1640: rom = 1'b0;
		1641: rom = 1'b0;
		1642: rom = 1'b0;
		1643: rom = 1'b0;
		1644: rom = 1'b0;
		1645: rom = 1'b0;
		1646: rom = 1'b0;
		1647: rom = 1'b0;
		1648: rom = 1'b0;
		1649: rom = 1'b0;
		1650: rom = 1'b0;
		1651: rom = 1'b0;
		1652: rom = 1'b0;
		1653: rom = 1'b0;
		1654: rom = 1'b0;
		1655: rom = 1'b0;
		1656: rom = 1'b0;
		1657: rom = 1'b0;
		1658: rom = 1'b0;
		1659: rom = 1'b0;
		1660: rom = 1'b0;
		1661: rom = 1'b0;
		1662: rom = 1'b0;
		1663: rom = 1'b0;
		1664: rom = 1'b0;
		1665: rom = 1'b0;
		1666: rom = 1'b0;
		1667: rom = 1'b0;
		1668: rom = 1'b0;
		1669: rom = 1'b0;
		1670: rom = 1'b0;
		1671: rom = 1'b0;
		1672: rom = 1'b0;
		1673: rom = 1'b0;
		1674: rom = 1'b0;
		1675: rom = 1'b0;
		1676: rom = 1'b0;
		1677: rom = 1'b0;
		1678: rom = 1'b0;
		1679: rom = 1'b0;
		1680: rom = 1'b0;
		1681: rom = 1'b0;
		1682: rom = 1'b0;
		1683: rom = 1'b0;
		1684: rom = 1'b0;
		1685: rom = 1'b0;
		1686: rom = 1'b0;
		1687: rom = 1'b0;
		1688: rom = 1'b0;
		1689: rom = 1'b0;
		1690: rom = 1'b0;
		1691: rom = 1'b0;
		1692: rom = 1'b0;
		1693: rom = 1'b0;
		1694: rom = 1'b0;
		1695: rom = 1'b0;
		1696: rom = 1'b0;
		1697: rom = 1'b0;
		1698: rom = 1'b0;
		1699: rom = 1'b0;
		1700: rom = 1'b0;
		1701: rom = 1'b0;
		1702: rom = 1'b0;
		1703: rom = 1'b0;
		1704: rom = 1'b0;
		1705: rom = 1'b0;
		1706: rom = 1'b0;
		1707: rom = 1'b0;
		1708: rom = 1'b0;
		1709: rom = 1'b1;
		1710: rom = 1'b1;
		1711: rom = 1'b1;
		1712: rom = 1'b1;
		1713: rom = 1'b1;
		1714: rom = 1'b1;
		1715: rom = 1'b1;
		1716: rom = 1'b1;
		1717: rom = 1'b1;
		1718: rom = 1'b1;
		1719: rom = 1'b1;
		1720: rom = 1'b1;
		1721: rom = 1'b1;
		1722: rom = 1'b1;
		1723: rom = 1'b1;
		1724: rom = 1'b1;
		1725: rom = 1'b1;
		1726: rom = 1'b1;
		1727: rom = 1'b1;
		1728: rom = 1'b1;
		1729: rom = 1'b0;
		1730: rom = 1'b0;
		1731: rom = 1'b0;
		1732: rom = 1'b0;
		1733: rom = 1'b0;
		1734: rom = 1'b0;
		1735: rom = 1'b0;
		1736: rom = 1'b0;
		1737: rom = 1'b0;
		1738: rom = 1'b0;
		1739: rom = 1'b0;
		1740: rom = 1'b0;
		1741: rom = 1'b0;
		1742: rom = 1'b0;
		1743: rom = 1'b0;
		1744: rom = 1'b0;
		1745: rom = 1'b0;
		1746: rom = 1'b1;
		1747: rom = 1'b1;
		1748: rom = 1'b1;
		1749: rom = 1'b1;
		1750: rom = 1'b1;
		1751: rom = 1'b1;
		1752: rom = 1'b1;
		1753: rom = 1'b1;
		1754: rom = 1'b1;
		1755: rom = 1'b1;
		1756: rom = 1'b1;
		1757: rom = 1'b1;
		1758: rom = 1'b1;
		1759: rom = 1'b1;
		1760: rom = 1'b1;
		1761: rom = 1'b1;
		1762: rom = 1'b1;
		1763: rom = 1'b1;
		1764: rom = 1'b1;
		1765: rom = 1'b0;
		1766: rom = 1'b0;
		1767: rom = 1'b0;
		1768: rom = 1'b0;
		1769: rom = 1'b0;
		1770: rom = 1'b0;
		1771: rom = 1'b0;
		1772: rom = 1'b0;
		1773: rom = 1'b0;
		1774: rom = 1'b0;
		1775: rom = 1'b0;
		1776: rom = 1'b0;
		1777: rom = 1'b0;
		1778: rom = 1'b0;
		1779: rom = 1'b0;
		1780: rom = 1'b0;
		1781: rom = 1'b0;
		1782: rom = 1'b0;
		1783: rom = 1'b0;
		1784: rom = 1'b0;
		1785: rom = 1'b0;
		1786: rom = 1'b0;
		1787: rom = 1'b0;
		1788: rom = 1'b0;
		1789: rom = 1'b0;
		1790: rom = 1'b0;
		1791: rom = 1'b0;
		1792: rom = 1'b0;
		1793: rom = 1'b0;
		1794: rom = 1'b0;
		1795: rom = 1'b0;
		1796: rom = 1'b0;
		1797: rom = 1'b0;
		1798: rom = 1'b0;
		1799: rom = 1'b0;
		1800: rom = 1'b0;
		1801: rom = 1'b0;
		1802: rom = 1'b0;
		1803: rom = 1'b0;
		1804: rom = 1'b0;
		1805: rom = 1'b0;
		1806: rom = 1'b0;
		1807: rom = 1'b0;
		1808: rom = 1'b0;
		1809: rom = 1'b0;
		1810: rom = 1'b0;
		1811: rom = 1'b0;
		1812: rom = 1'b0;
		1813: rom = 1'b0;
		1814: rom = 1'b0;
		1815: rom = 1'b0;
		1816: rom = 1'b0;
		1817: rom = 1'b0;
		1818: rom = 1'b0;
		1819: rom = 1'b0;
		1820: rom = 1'b0;
		1821: rom = 1'b0;
		1822: rom = 1'b0;
		1823: rom = 1'b0;
		1824: rom = 1'b0;
		1825: rom = 1'b0;
		1826: rom = 1'b0;
		1827: rom = 1'b0;
		1828: rom = 1'b0;
		1829: rom = 1'b0;
		1830: rom = 1'b0;
		1831: rom = 1'b0;
		1832: rom = 1'b0;
		1833: rom = 1'b0;
		1834: rom = 1'b0;
		1835: rom = 1'b1;
		1836: rom = 1'b1;
		1837: rom = 1'b1;
		1838: rom = 1'b1;
		1839: rom = 1'b1;
		1840: rom = 1'b1;
		1841: rom = 1'b1;
		1842: rom = 1'b1;
		1843: rom = 1'b1;
		1844: rom = 1'b1;
		1845: rom = 1'b1;
		1846: rom = 1'b1;
		1847: rom = 1'b1;
		1848: rom = 1'b1;
		1849: rom = 1'b1;
		1850: rom = 1'b1;
		1851: rom = 1'b1;
		1852: rom = 1'b1;
		1853: rom = 1'b1;
		1854: rom = 1'b1;
		1855: rom = 1'b0;
		1856: rom = 1'b0;
		1857: rom = 1'b0;
		1858: rom = 1'b0;
		1859: rom = 1'b0;
		1860: rom = 1'b0;
		1861: rom = 1'b0;
		1862: rom = 1'b0;
		1863: rom = 1'b0;
		1864: rom = 1'b0;
		1865: rom = 1'b0;
		1866: rom = 1'b0;
		1867: rom = 1'b0;
		1868: rom = 1'b0;
		1869: rom = 1'b0;
		1870: rom = 1'b0;
		1871: rom = 1'b0;
		1872: rom = 1'b1;
		1873: rom = 1'b1;
		1874: rom = 1'b1;
		1875: rom = 1'b1;
		1876: rom = 1'b1;
		1877: rom = 1'b1;
		1878: rom = 1'b1;
		1879: rom = 1'b1;
		1880: rom = 1'b1;
		1881: rom = 1'b1;
		1882: rom = 1'b1;
		1883: rom = 1'b1;
		1884: rom = 1'b1;
		1885: rom = 1'b1;
		1886: rom = 1'b1;
		1887: rom = 1'b1;
		1888: rom = 1'b1;
		1889: rom = 1'b1;
		1890: rom = 1'b1;
		1891: rom = 1'b1;
		1892: rom = 1'b1;
		1893: rom = 1'b1;
		1894: rom = 1'b1;
		1895: rom = 1'b0;
		1896: rom = 1'b0;
		1897: rom = 1'b0;
		1898: rom = 1'b0;
		1899: rom = 1'b0;
		1900: rom = 1'b0;
		1901: rom = 1'b0;
		1902: rom = 1'b0;
		1903: rom = 1'b0;
		1904: rom = 1'b0;
		1905: rom = 1'b0;
		1906: rom = 1'b0;
		1907: rom = 1'b0;
		1908: rom = 1'b0;
		1909: rom = 1'b0;
		1910: rom = 1'b0;
		1911: rom = 1'b0;
		1912: rom = 1'b0;
		1913: rom = 1'b0;
		1914: rom = 1'b0;
		1915: rom = 1'b0;
		1916: rom = 1'b0;
		1917: rom = 1'b0;
		1918: rom = 1'b0;
		1919: rom = 1'b0;
		1920: rom = 1'b0;
		1921: rom = 1'b0;
		1922: rom = 1'b0;
		1923: rom = 1'b0;
		1924: rom = 1'b0;
		1925: rom = 1'b0;
		1926: rom = 1'b0;
		1927: rom = 1'b0;
		1928: rom = 1'b0;
		1929: rom = 1'b0;
		1930: rom = 1'b0;
		1931: rom = 1'b0;
		1932: rom = 1'b0;
		1933: rom = 1'b0;
		1934: rom = 1'b0;
		1935: rom = 1'b0;
		1936: rom = 1'b0;
		1937: rom = 1'b0;
		1938: rom = 1'b0;
		1939: rom = 1'b0;
		1940: rom = 1'b0;
		1941: rom = 1'b0;
		1942: rom = 1'b0;
		1943: rom = 1'b0;
		1944: rom = 1'b0;
		1945: rom = 1'b0;
		1946: rom = 1'b0;
		1947: rom = 1'b0;
		1948: rom = 1'b0;
		1949: rom = 1'b0;
		1950: rom = 1'b0;
		1951: rom = 1'b0;
		1952: rom = 1'b0;
		1953: rom = 1'b0;
		1954: rom = 1'b0;
		1955: rom = 1'b0;
		1956: rom = 1'b0;
		1957: rom = 1'b0;
		1958: rom = 1'b0;
		1959: rom = 1'b0;
		1960: rom = 1'b0;
		1961: rom = 1'b0;
		1962: rom = 1'b0;
		1963: rom = 1'b1;
		1964: rom = 1'b1;
		1965: rom = 1'b1;
		1966: rom = 1'b1;
		1967: rom = 1'b1;
		1968: rom = 1'b1;
		1969: rom = 1'b1;
		1970: rom = 1'b1;
		1971: rom = 1'b1;
		1972: rom = 1'b1;
		1973: rom = 1'b1;
		1974: rom = 1'b1;
		1975: rom = 1'b1;
		1976: rom = 1'b1;
		1977: rom = 1'b1;
		1978: rom = 1'b1;
		1979: rom = 1'b1;
		1980: rom = 1'b1;
		1981: rom = 1'b1;
		1982: rom = 1'b0;
		1983: rom = 1'b0;
		1984: rom = 1'b0;
		1985: rom = 1'b0;
		1986: rom = 1'b0;
		1987: rom = 1'b0;
		1988: rom = 1'b0;
		1989: rom = 1'b0;
		1990: rom = 1'b0;
		1991: rom = 1'b0;
		1992: rom = 1'b0;
		1993: rom = 1'b0;
		1994: rom = 1'b0;
		1995: rom = 1'b0;
		1996: rom = 1'b0;
		1997: rom = 1'b0;
		1998: rom = 1'b1;
		1999: rom = 1'b1;
		2000: rom = 1'b1;
		2001: rom = 1'b1;
		2002: rom = 1'b1;
		2003: rom = 1'b1;
		2004: rom = 1'b1;
		2005: rom = 1'b1;
		2006: rom = 1'b1;
		2007: rom = 1'b1;
		2008: rom = 1'b1;
		2009: rom = 1'b1;
		2010: rom = 1'b1;
		2011: rom = 1'b1;
		2012: rom = 1'b1;
		2013: rom = 1'b1;
		2014: rom = 1'b1;
		2015: rom = 1'b1;
		2016: rom = 1'b1;
		2017: rom = 1'b1;
		2018: rom = 1'b1;
		2019: rom = 1'b1;
		2020: rom = 1'b1;
		2021: rom = 1'b1;
		2022: rom = 1'b1;
		2023: rom = 1'b0;
		2024: rom = 1'b0;
		2025: rom = 1'b0;
		2026: rom = 1'b0;
		2027: rom = 1'b0;
		2028: rom = 1'b0;
		2029: rom = 1'b0;
		2030: rom = 1'b0;
		2031: rom = 1'b0;
		2032: rom = 1'b0;
		2033: rom = 1'b0;
		2034: rom = 1'b0;
		2035: rom = 1'b0;
		2036: rom = 1'b0;
		2037: rom = 1'b0;
		2038: rom = 1'b0;
		2039: rom = 1'b0;
		2040: rom = 1'b0;
		2041: rom = 1'b0;
		2042: rom = 1'b0;
		2043: rom = 1'b0;
		2044: rom = 1'b0;
		2045: rom = 1'b0;
		2046: rom = 1'b0;
		2047: rom = 1'b0;
		2048: rom = 1'b0;
		2049: rom = 1'b0;
		2050: rom = 1'b0;
		2051: rom = 1'b0;
		2052: rom = 1'b0;
		2053: rom = 1'b0;
		2054: rom = 1'b0;
		2055: rom = 1'b0;
		2056: rom = 1'b0;
		2057: rom = 1'b0;
		2058: rom = 1'b0;
		2059: rom = 1'b0;
		2060: rom = 1'b0;
		2061: rom = 1'b0;
		2062: rom = 1'b0;
		2063: rom = 1'b0;
		2064: rom = 1'b0;
		2065: rom = 1'b0;
		2066: rom = 1'b0;
		2067: rom = 1'b0;
		2068: rom = 1'b0;
		2069: rom = 1'b0;
		2070: rom = 1'b0;
		2071: rom = 1'b0;
		2072: rom = 1'b0;
		2073: rom = 1'b0;
		2074: rom = 1'b0;
		2075: rom = 1'b0;
		2076: rom = 1'b0;
		2077: rom = 1'b0;
		2078: rom = 1'b0;
		2079: rom = 1'b0;
		2080: rom = 1'b0;
		2081: rom = 1'b0;
		2082: rom = 1'b0;
		2083: rom = 1'b0;
		2084: rom = 1'b0;
		2085: rom = 1'b0;
		2086: rom = 1'b0;
		2087: rom = 1'b0;
		2088: rom = 1'b0;
		2089: rom = 1'b1;
		2090: rom = 1'b1;
		2091: rom = 1'b1;
		2092: rom = 1'b1;
		2093: rom = 1'b1;
		2094: rom = 1'b1;
		2095: rom = 1'b1;
		2096: rom = 1'b1;
		2097: rom = 1'b1;
		2098: rom = 1'b1;
		2099: rom = 1'b1;
		2100: rom = 1'b1;
		2101: rom = 1'b1;
		2102: rom = 1'b1;
		2103: rom = 1'b1;
		2104: rom = 1'b1;
		2105: rom = 1'b1;
		2106: rom = 1'b1;
		2107: rom = 1'b1;
		2108: rom = 1'b0;
		2109: rom = 1'b0;
		2110: rom = 1'b0;
		2111: rom = 1'b0;
		2112: rom = 1'b0;
		2113: rom = 1'b0;
		2114: rom = 1'b0;
		2115: rom = 1'b0;
		2116: rom = 1'b0;
		2117: rom = 1'b0;
		2118: rom = 1'b0;
		2119: rom = 1'b0;
		2120: rom = 1'b0;
		2121: rom = 1'b0;
		2122: rom = 1'b0;
		2123: rom = 1'b0;
		2124: rom = 1'b1;
		2125: rom = 1'b1;
		2126: rom = 1'b1;
		2127: rom = 1'b1;
		2128: rom = 1'b1;
		2129: rom = 1'b1;
		2130: rom = 1'b1;
		2131: rom = 1'b1;
		2132: rom = 1'b1;
		2133: rom = 1'b1;
		2134: rom = 1'b1;
		2135: rom = 1'b1;
		2136: rom = 1'b1;
		2137: rom = 1'b1;
		2138: rom = 1'b1;
		2139: rom = 1'b1;
		2140: rom = 1'b1;
		2141: rom = 1'b1;
		2142: rom = 1'b1;
		2143: rom = 1'b1;
		2144: rom = 1'b1;
		2145: rom = 1'b1;
		2146: rom = 1'b1;
		2147: rom = 1'b1;
		2148: rom = 1'b1;
		2149: rom = 1'b1;
		2150: rom = 1'b1;
		2151: rom = 1'b1;
		2152: rom = 1'b1;
		2153: rom = 1'b0;
		2154: rom = 1'b0;
		2155: rom = 1'b0;
		2156: rom = 1'b0;
		2157: rom = 1'b0;
		2158: rom = 1'b0;
		2159: rom = 1'b0;
		2160: rom = 1'b0;
		2161: rom = 1'b0;
		2162: rom = 1'b0;
		2163: rom = 1'b0;
		2164: rom = 1'b0;
		2165: rom = 1'b0;
		2166: rom = 1'b0;
		2167: rom = 1'b0;
		2168: rom = 1'b0;
		2169: rom = 1'b0;
		2170: rom = 1'b0;
		2171: rom = 1'b0;
		2172: rom = 1'b0;
		2173: rom = 1'b0;
		2174: rom = 1'b0;
		2175: rom = 1'b0;
		2176: rom = 1'b0;
		2177: rom = 1'b0;
		2178: rom = 1'b0;
		2179: rom = 1'b0;
		2180: rom = 1'b0;
		2181: rom = 1'b0;
		2182: rom = 1'b0;
		2183: rom = 1'b0;
		2184: rom = 1'b0;
		2185: rom = 1'b0;
		2186: rom = 1'b0;
		2187: rom = 1'b0;
		2188: rom = 1'b0;
		2189: rom = 1'b0;
		2190: rom = 1'b0;
		2191: rom = 1'b0;
		2192: rom = 1'b0;
		2193: rom = 1'b0;
		2194: rom = 1'b0;
		2195: rom = 1'b0;
		2196: rom = 1'b0;
		2197: rom = 1'b0;
		2198: rom = 1'b0;
		2199: rom = 1'b0;
		2200: rom = 1'b0;
		2201: rom = 1'b0;
		2202: rom = 1'b0;
		2203: rom = 1'b0;
		2204: rom = 1'b0;
		2205: rom = 1'b0;
		2206: rom = 1'b0;
		2207: rom = 1'b0;
		2208: rom = 1'b0;
		2209: rom = 1'b0;
		2210: rom = 1'b0;
		2211: rom = 1'b0;
		2212: rom = 1'b0;
		2213: rom = 1'b0;
		2214: rom = 1'b0;
		2215: rom = 1'b0;
		2216: rom = 1'b1;
		2217: rom = 1'b1;
		2218: rom = 1'b1;
		2219: rom = 1'b1;
		2220: rom = 1'b1;
		2221: rom = 1'b1;
		2222: rom = 1'b1;
		2223: rom = 1'b1;
		2224: rom = 1'b1;
		2225: rom = 1'b1;
		2226: rom = 1'b1;
		2227: rom = 1'b1;
		2228: rom = 1'b1;
		2229: rom = 1'b1;
		2230: rom = 1'b1;
		2231: rom = 1'b1;
		2232: rom = 1'b1;
		2233: rom = 1'b1;
		2234: rom = 1'b1;
		2235: rom = 1'b0;
		2236: rom = 1'b0;
		2237: rom = 1'b0;
		2238: rom = 1'b0;
		2239: rom = 1'b0;
		2240: rom = 1'b0;
		2241: rom = 1'b0;
		2242: rom = 1'b0;
		2243: rom = 1'b0;
		2244: rom = 1'b0;
		2245: rom = 1'b0;
		2246: rom = 1'b0;
		2247: rom = 1'b0;
		2248: rom = 1'b0;
		2249: rom = 1'b0;
		2250: rom = 1'b1;
		2251: rom = 1'b1;
		2252: rom = 1'b1;
		2253: rom = 1'b1;
		2254: rom = 1'b1;
		2255: rom = 1'b1;
		2256: rom = 1'b1;
		2257: rom = 1'b1;
		2258: rom = 1'b1;
		2259: rom = 1'b1;
		2260: rom = 1'b1;
		2261: rom = 1'b1;
		2262: rom = 1'b1;
		2263: rom = 1'b1;
		2264: rom = 1'b1;
		2265: rom = 1'b1;
		2266: rom = 1'b1;
		2267: rom = 1'b1;
		2268: rom = 1'b1;
		2269: rom = 1'b1;
		2270: rom = 1'b1;
		2271: rom = 1'b1;
		2272: rom = 1'b1;
		2273: rom = 1'b1;
		2274: rom = 1'b1;
		2275: rom = 1'b1;
		2276: rom = 1'b1;
		2277: rom = 1'b1;
		2278: rom = 1'b1;
		2279: rom = 1'b1;
		2280: rom = 1'b1;
		2281: rom = 1'b1;
		2282: rom = 1'b0;
		2283: rom = 1'b0;
		2284: rom = 1'b0;
		2285: rom = 1'b0;
		2286: rom = 1'b0;
		2287: rom = 1'b0;
		2288: rom = 1'b0;
		2289: rom = 1'b0;
		2290: rom = 1'b0;
		2291: rom = 1'b0;
		2292: rom = 1'b0;
		2293: rom = 1'b0;
		2294: rom = 1'b0;
		2295: rom = 1'b0;
		2296: rom = 1'b0;
		2297: rom = 1'b0;
		2298: rom = 1'b0;
		2299: rom = 1'b0;
		2300: rom = 1'b0;
		2301: rom = 1'b0;
		2302: rom = 1'b0;
		2303: rom = 1'b0;
		2304: rom = 1'b0;
		2305: rom = 1'b0;
		2306: rom = 1'b0;
		2307: rom = 1'b0;
		2308: rom = 1'b0;
		2309: rom = 1'b0;
		2310: rom = 1'b0;
		2311: rom = 1'b0;
		2312: rom = 1'b0;
		2313: rom = 1'b0;
		2314: rom = 1'b0;
		2315: rom = 1'b0;
		2316: rom = 1'b0;
		2317: rom = 1'b0;
		2318: rom = 1'b0;
		2319: rom = 1'b0;
		2320: rom = 1'b0;
		2321: rom = 1'b0;
		2322: rom = 1'b0;
		2323: rom = 1'b0;
		2324: rom = 1'b0;
		2325: rom = 1'b0;
		2326: rom = 1'b0;
		2327: rom = 1'b0;
		2328: rom = 1'b0;
		2329: rom = 1'b0;
		2330: rom = 1'b0;
		2331: rom = 1'b0;
		2332: rom = 1'b0;
		2333: rom = 1'b0;
		2334: rom = 1'b0;
		2335: rom = 1'b0;
		2336: rom = 1'b0;
		2337: rom = 1'b0;
		2338: rom = 1'b0;
		2339: rom = 1'b0;
		2340: rom = 1'b0;
		2341: rom = 1'b0;
		2342: rom = 1'b0;
		2343: rom = 1'b1;
		2344: rom = 1'b1;
		2345: rom = 1'b1;
		2346: rom = 1'b1;
		2347: rom = 1'b1;
		2348: rom = 1'b1;
		2349: rom = 1'b1;
		2350: rom = 1'b1;
		2351: rom = 1'b1;
		2352: rom = 1'b1;
		2353: rom = 1'b1;
		2354: rom = 1'b1;
		2355: rom = 1'b1;
		2356: rom = 1'b1;
		2357: rom = 1'b1;
		2358: rom = 1'b1;
		2359: rom = 1'b1;
		2360: rom = 1'b1;
		2361: rom = 1'b0;
		2362: rom = 1'b0;
		2363: rom = 1'b0;
		2364: rom = 1'b0;
		2365: rom = 1'b0;
		2366: rom = 1'b0;
		2367: rom = 1'b0;
		2368: rom = 1'b0;
		2369: rom = 1'b0;
		2370: rom = 1'b0;
		2371: rom = 1'b0;
		2372: rom = 1'b0;
		2373: rom = 1'b0;
		2374: rom = 1'b0;
		2375: rom = 1'b0;
		2376: rom = 1'b1;
		2377: rom = 1'b1;
		2378: rom = 1'b1;
		2379: rom = 1'b1;
		2380: rom = 1'b1;
		2381: rom = 1'b1;
		2382: rom = 1'b1;
		2383: rom = 1'b1;
		2384: rom = 1'b1;
		2385: rom = 1'b1;
		2386: rom = 1'b1;
		2387: rom = 1'b1;
		2388: rom = 1'b1;
		2389: rom = 1'b1;
		2390: rom = 1'b1;
		2391: rom = 1'b1;
		2392: rom = 1'b1;
		2393: rom = 1'b1;
		2394: rom = 1'b1;
		2395: rom = 1'b1;
		2396: rom = 1'b1;
		2397: rom = 1'b1;
		2398: rom = 1'b1;
		2399: rom = 1'b1;
		2400: rom = 1'b1;
		2401: rom = 1'b1;
		2402: rom = 1'b1;
		2403: rom = 1'b1;
		2404: rom = 1'b1;
		2405: rom = 1'b1;
		2406: rom = 1'b1;
		2407: rom = 1'b1;
		2408: rom = 1'b1;
		2409: rom = 1'b1;
		2410: rom = 1'b1;
		2411: rom = 1'b0;
		2412: rom = 1'b0;
		2413: rom = 1'b0;
		2414: rom = 1'b0;
		2415: rom = 1'b0;
		2416: rom = 1'b0;
		2417: rom = 1'b0;
		2418: rom = 1'b0;
		2419: rom = 1'b0;
		2420: rom = 1'b0;
		2421: rom = 1'b0;
		2422: rom = 1'b0;
		2423: rom = 1'b0;
		2424: rom = 1'b0;
		2425: rom = 1'b0;
		2426: rom = 1'b0;
		2427: rom = 1'b0;
		2428: rom = 1'b0;
		2429: rom = 1'b0;
		2430: rom = 1'b0;
		2431: rom = 1'b0;
		2432: rom = 1'b0;
		2433: rom = 1'b0;
		2434: rom = 1'b0;
		2435: rom = 1'b0;
		2436: rom = 1'b0;
		2437: rom = 1'b0;
		2438: rom = 1'b0;
		2439: rom = 1'b0;
		2440: rom = 1'b0;
		2441: rom = 1'b0;
		2442: rom = 1'b0;
		2443: rom = 1'b0;
		2444: rom = 1'b0;
		2445: rom = 1'b0;
		2446: rom = 1'b0;
		2447: rom = 1'b0;
		2448: rom = 1'b0;
		2449: rom = 1'b0;
		2450: rom = 1'b0;
		2451: rom = 1'b0;
		2452: rom = 1'b0;
		2453: rom = 1'b0;
		2454: rom = 1'b0;
		2455: rom = 1'b0;
		2456: rom = 1'b0;
		2457: rom = 1'b0;
		2458: rom = 1'b0;
		2459: rom = 1'b0;
		2460: rom = 1'b0;
		2461: rom = 1'b0;
		2462: rom = 1'b0;
		2463: rom = 1'b0;
		2464: rom = 1'b0;
		2465: rom = 1'b0;
		2466: rom = 1'b0;
		2467: rom = 1'b0;
		2468: rom = 1'b0;
		2469: rom = 1'b0;
		2470: rom = 1'b0;
		2471: rom = 1'b1;
		2472: rom = 1'b1;
		2473: rom = 1'b1;
		2474: rom = 1'b1;
		2475: rom = 1'b1;
		2476: rom = 1'b1;
		2477: rom = 1'b1;
		2478: rom = 1'b1;
		2479: rom = 1'b1;
		2480: rom = 1'b1;
		2481: rom = 1'b1;
		2482: rom = 1'b1;
		2483: rom = 1'b1;
		2484: rom = 1'b1;
		2485: rom = 1'b1;
		2486: rom = 1'b1;
		2487: rom = 1'b1;
		2488: rom = 1'b0;
		2489: rom = 1'b0;
		2490: rom = 1'b0;
		2491: rom = 1'b0;
		2492: rom = 1'b0;
		2493: rom = 1'b0;
		2494: rom = 1'b0;
		2495: rom = 1'b0;
		2496: rom = 1'b0;
		2497: rom = 1'b0;
		2498: rom = 1'b0;
		2499: rom = 1'b0;
		2500: rom = 1'b0;
		2501: rom = 1'b0;
		2502: rom = 1'b0;
		2503: rom = 1'b1;
		2504: rom = 1'b1;
		2505: rom = 1'b1;
		2506: rom = 1'b1;
		2507: rom = 1'b1;
		2508: rom = 1'b1;
		2509: rom = 1'b1;
		2510: rom = 1'b1;
		2511: rom = 1'b1;
		2512: rom = 1'b1;
		2513: rom = 1'b1;
		2514: rom = 1'b1;
		2515: rom = 1'b1;
		2516: rom = 1'b1;
		2517: rom = 1'b1;
		2518: rom = 1'b1;
		2519: rom = 1'b1;
		2520: rom = 1'b1;
		2521: rom = 1'b1;
		2522: rom = 1'b1;
		2523: rom = 1'b1;
		2524: rom = 1'b1;
		2525: rom = 1'b1;
		2526: rom = 1'b1;
		2527: rom = 1'b1;
		2528: rom = 1'b1;
		2529: rom = 1'b1;
		2530: rom = 1'b1;
		2531: rom = 1'b1;
		2532: rom = 1'b1;
		2533: rom = 1'b1;
		2534: rom = 1'b1;
		2535: rom = 1'b1;
		2536: rom = 1'b1;
		2537: rom = 1'b1;
		2538: rom = 1'b1;
		2539: rom = 1'b1;
		2540: rom = 1'b0;
		2541: rom = 1'b0;
		2542: rom = 1'b0;
		2543: rom = 1'b0;
		2544: rom = 1'b0;
		2545: rom = 1'b0;
		2546: rom = 1'b0;
		2547: rom = 1'b0;
		2548: rom = 1'b0;
		2549: rom = 1'b0;
		2550: rom = 1'b0;
		2551: rom = 1'b0;
		2552: rom = 1'b0;
		2553: rom = 1'b0;
		2554: rom = 1'b0;
		2555: rom = 1'b0;
		2556: rom = 1'b0;
		2557: rom = 1'b0;
		2558: rom = 1'b0;
		2559: rom = 1'b0;
		2560: rom = 1'b0;
		2561: rom = 1'b0;
		2562: rom = 1'b0;
		2563: rom = 1'b0;
		2564: rom = 1'b0;
		2565: rom = 1'b0;
		2566: rom = 1'b0;
		2567: rom = 1'b0;
		2568: rom = 1'b0;
		2569: rom = 1'b0;
		2570: rom = 1'b0;
		2571: rom = 1'b0;
		2572: rom = 1'b0;
		2573: rom = 1'b0;
		2574: rom = 1'b0;
		2575: rom = 1'b0;
		2576: rom = 1'b0;
		2577: rom = 1'b0;
		2578: rom = 1'b0;
		2579: rom = 1'b0;
		2580: rom = 1'b0;
		2581: rom = 1'b0;
		2582: rom = 1'b0;
		2583: rom = 1'b0;
		2584: rom = 1'b0;
		2585: rom = 1'b0;
		2586: rom = 1'b0;
		2587: rom = 1'b0;
		2588: rom = 1'b0;
		2589: rom = 1'b0;
		2590: rom = 1'b0;
		2591: rom = 1'b0;
		2592: rom = 1'b0;
		2593: rom = 1'b0;
		2594: rom = 1'b0;
		2595: rom = 1'b0;
		2596: rom = 1'b0;
		2597: rom = 1'b1;
		2598: rom = 1'b1;
		2599: rom = 1'b1;
		2600: rom = 1'b1;
		2601: rom = 1'b1;
		2602: rom = 1'b1;
		2603: rom = 1'b1;
		2604: rom = 1'b1;
		2605: rom = 1'b1;
		2606: rom = 1'b1;
		2607: rom = 1'b1;
		2608: rom = 1'b1;
		2609: rom = 1'b1;
		2610: rom = 1'b1;
		2611: rom = 1'b1;
		2612: rom = 1'b1;
		2613: rom = 1'b1;
		2614: rom = 1'b0;
		2615: rom = 1'b0;
		2616: rom = 1'b0;
		2617: rom = 1'b0;
		2618: rom = 1'b0;
		2619: rom = 1'b0;
		2620: rom = 1'b0;
		2621: rom = 1'b0;
		2622: rom = 1'b0;
		2623: rom = 1'b0;
		2624: rom = 1'b0;
		2625: rom = 1'b0;
		2626: rom = 1'b0;
		2627: rom = 1'b0;
		2628: rom = 1'b0;
		2629: rom = 1'b1;
		2630: rom = 1'b1;
		2631: rom = 1'b1;
		2632: rom = 1'b1;
		2633: rom = 1'b1;
		2634: rom = 1'b1;
		2635: rom = 1'b1;
		2636: rom = 1'b1;
		2637: rom = 1'b1;
		2638: rom = 1'b1;
		2639: rom = 1'b1;
		2640: rom = 1'b1;
		2641: rom = 1'b1;
		2642: rom = 1'b1;
		2643: rom = 1'b1;
		2644: rom = 1'b1;
		2645: rom = 1'b1;
		2646: rom = 1'b1;
		2647: rom = 1'b1;
		2648: rom = 1'b1;
		2649: rom = 1'b1;
		2650: rom = 1'b1;
		2651: rom = 1'b1;
		2652: rom = 1'b1;
		2653: rom = 1'b1;
		2654: rom = 1'b1;
		2655: rom = 1'b1;
		2656: rom = 1'b1;
		2657: rom = 1'b1;
		2658: rom = 1'b1;
		2659: rom = 1'b1;
		2660: rom = 1'b1;
		2661: rom = 1'b1;
		2662: rom = 1'b1;
		2663: rom = 1'b1;
		2664: rom = 1'b1;
		2665: rom = 1'b1;
		2666: rom = 1'b1;
		2667: rom = 1'b1;
		2668: rom = 1'b1;
		2669: rom = 1'b0;
		2670: rom = 1'b0;
		2671: rom = 1'b0;
		2672: rom = 1'b0;
		2673: rom = 1'b0;
		2674: rom = 1'b0;
		2675: rom = 1'b0;
		2676: rom = 1'b0;
		2677: rom = 1'b0;
		2678: rom = 1'b0;
		2679: rom = 1'b0;
		2680: rom = 1'b0;
		2681: rom = 1'b0;
		2682: rom = 1'b0;
		2683: rom = 1'b0;
		2684: rom = 1'b0;
		2685: rom = 1'b0;
		2686: rom = 1'b0;
		2687: rom = 1'b0;
		2688: rom = 1'b0;
		2689: rom = 1'b0;
		2690: rom = 1'b0;
		2691: rom = 1'b0;
		2692: rom = 1'b0;
		2693: rom = 1'b0;
		2694: rom = 1'b0;
		2695: rom = 1'b0;
		2696: rom = 1'b0;
		2697: rom = 1'b0;
		2698: rom = 1'b0;
		2699: rom = 1'b0;
		2700: rom = 1'b0;
		2701: rom = 1'b0;
		2702: rom = 1'b0;
		2703: rom = 1'b0;
		2704: rom = 1'b0;
		2705: rom = 1'b0;
		2706: rom = 1'b0;
		2707: rom = 1'b0;
		2708: rom = 1'b0;
		2709: rom = 1'b0;
		2710: rom = 1'b0;
		2711: rom = 1'b0;
		2712: rom = 1'b0;
		2713: rom = 1'b0;
		2714: rom = 1'b0;
		2715: rom = 1'b0;
		2716: rom = 1'b0;
		2717: rom = 1'b0;
		2718: rom = 1'b0;
		2719: rom = 1'b0;
		2720: rom = 1'b0;
		2721: rom = 1'b0;
		2722: rom = 1'b0;
		2723: rom = 1'b0;
		2724: rom = 1'b0;
		2725: rom = 1'b1;
		2726: rom = 1'b1;
		2727: rom = 1'b1;
		2728: rom = 1'b1;
		2729: rom = 1'b1;
		2730: rom = 1'b1;
		2731: rom = 1'b1;
		2732: rom = 1'b1;
		2733: rom = 1'b1;
		2734: rom = 1'b1;
		2735: rom = 1'b1;
		2736: rom = 1'b1;
		2737: rom = 1'b1;
		2738: rom = 1'b1;
		2739: rom = 1'b1;
		2740: rom = 1'b1;
		2741: rom = 1'b0;
		2742: rom = 1'b0;
		2743: rom = 1'b0;
		2744: rom = 1'b0;
		2745: rom = 1'b0;
		2746: rom = 1'b0;
		2747: rom = 1'b0;
		2748: rom = 1'b0;
		2749: rom = 1'b0;
		2750: rom = 1'b0;
		2751: rom = 1'b0;
		2752: rom = 1'b0;
		2753: rom = 1'b0;
		2754: rom = 1'b0;
		2755: rom = 1'b1;
		2756: rom = 1'b1;
		2757: rom = 1'b1;
		2758: rom = 1'b1;
		2759: rom = 1'b1;
		2760: rom = 1'b1;
		2761: rom = 1'b1;
		2762: rom = 1'b1;
		2763: rom = 1'b1;
		2764: rom = 1'b1;
		2765: rom = 1'b1;
		2766: rom = 1'b1;
		2767: rom = 1'b1;
		2768: rom = 1'b1;
		2769: rom = 1'b1;
		2770: rom = 1'b1;
		2771: rom = 1'b1;
		2772: rom = 1'b1;
		2773: rom = 1'b1;
		2774: rom = 1'b1;
		2775: rom = 1'b1;
		2776: rom = 1'b1;
		2777: rom = 1'b1;
		2778: rom = 1'b1;
		2779: rom = 1'b1;
		2780: rom = 1'b1;
		2781: rom = 1'b1;
		2782: rom = 1'b1;
		2783: rom = 1'b1;
		2784: rom = 1'b1;
		2785: rom = 1'b1;
		2786: rom = 1'b1;
		2787: rom = 1'b1;
		2788: rom = 1'b1;
		2789: rom = 1'b1;
		2790: rom = 1'b1;
		2791: rom = 1'b1;
		2792: rom = 1'b1;
		2793: rom = 1'b1;
		2794: rom = 1'b1;
		2795: rom = 1'b1;
		2796: rom = 1'b1;
		2797: rom = 1'b0;
		2798: rom = 1'b0;
		2799: rom = 1'b0;
		2800: rom = 1'b0;
		2801: rom = 1'b0;
		2802: rom = 1'b0;
		2803: rom = 1'b0;
		2804: rom = 1'b0;
		2805: rom = 1'b0;
		2806: rom = 1'b0;
		2807: rom = 1'b0;
		2808: rom = 1'b0;
		2809: rom = 1'b1;
		2810: rom = 1'b0;
		2811: rom = 1'b0;
		2812: rom = 1'b0;
		2813: rom = 1'b0;
		2814: rom = 1'b0;
		2815: rom = 1'b0;
		2816: rom = 1'b0;
		2817: rom = 1'b0;
		2818: rom = 1'b0;
		2819: rom = 1'b0;
		2820: rom = 1'b0;
		2821: rom = 1'b0;
		2822: rom = 1'b0;
		2823: rom = 1'b0;
		2824: rom = 1'b0;
		2825: rom = 1'b0;
		2826: rom = 1'b0;
		2827: rom = 1'b0;
		2828: rom = 1'b0;
		2829: rom = 1'b0;
		2830: rom = 1'b0;
		2831: rom = 1'b0;
		2832: rom = 1'b0;
		2833: rom = 1'b0;
		2834: rom = 1'b0;
		2835: rom = 1'b0;
		2836: rom = 1'b0;
		2837: rom = 1'b0;
		2838: rom = 1'b0;
		2839: rom = 1'b0;
		2840: rom = 1'b0;
		2841: rom = 1'b0;
		2842: rom = 1'b0;
		2843: rom = 1'b0;
		2844: rom = 1'b0;
		2845: rom = 1'b0;
		2846: rom = 1'b0;
		2847: rom = 1'b0;
		2848: rom = 1'b0;
		2849: rom = 1'b0;
		2850: rom = 1'b0;
		2851: rom = 1'b0;
		2852: rom = 1'b1;
		2853: rom = 1'b1;
		2854: rom = 1'b1;
		2855: rom = 1'b1;
		2856: rom = 1'b1;
		2857: rom = 1'b1;
		2858: rom = 1'b1;
		2859: rom = 1'b1;
		2860: rom = 1'b1;
		2861: rom = 1'b1;
		2862: rom = 1'b1;
		2863: rom = 1'b1;
		2864: rom = 1'b1;
		2865: rom = 1'b1;
		2866: rom = 1'b1;
		2867: rom = 1'b1;
		2868: rom = 1'b0;
		2869: rom = 1'b0;
		2870: rom = 1'b0;
		2871: rom = 1'b0;
		2872: rom = 1'b0;
		2873: rom = 1'b0;
		2874: rom = 1'b0;
		2875: rom = 1'b0;
		2876: rom = 1'b0;
		2877: rom = 1'b0;
		2878: rom = 1'b0;
		2879: rom = 1'b0;
		2880: rom = 1'b0;
		2881: rom = 1'b0;
		2882: rom = 1'b1;
		2883: rom = 1'b1;
		2884: rom = 1'b1;
		2885: rom = 1'b1;
		2886: rom = 1'b1;
		2887: rom = 1'b1;
		2888: rom = 1'b1;
		2889: rom = 1'b1;
		2890: rom = 1'b1;
		2891: rom = 1'b1;
		2892: rom = 1'b1;
		2893: rom = 1'b1;
		2894: rom = 1'b1;
		2895: rom = 1'b1;
		2896: rom = 1'b1;
		2897: rom = 1'b1;
		2898: rom = 1'b1;
		2899: rom = 1'b1;
		2900: rom = 1'b1;
		2901: rom = 1'b1;
		2902: rom = 1'b1;
		2903: rom = 1'b1;
		2904: rom = 1'b1;
		2905: rom = 1'b1;
		2906: rom = 1'b1;
		2907: rom = 1'b1;
		2908: rom = 1'b1;
		2909: rom = 1'b1;
		2910: rom = 1'b1;
		2911: rom = 1'b1;
		2912: rom = 1'b1;
		2913: rom = 1'b1;
		2914: rom = 1'b1;
		2915: rom = 1'b1;
		2916: rom = 1'b1;
		2917: rom = 1'b1;
		2918: rom = 1'b1;
		2919: rom = 1'b1;
		2920: rom = 1'b1;
		2921: rom = 1'b1;
		2922: rom = 1'b1;
		2923: rom = 1'b1;
		2924: rom = 1'b1;
		2925: rom = 1'b1;
		2926: rom = 1'b0;
		2927: rom = 1'b0;
		2928: rom = 1'b0;
		2929: rom = 1'b0;
		2930: rom = 1'b0;
		2931: rom = 1'b0;
		2932: rom = 1'b0;
		2933: rom = 1'b0;
		2934: rom = 1'b0;
		2935: rom = 1'b0;
		2936: rom = 1'b0;
		2937: rom = 1'b1;
		2938: rom = 1'b0;
		2939: rom = 1'b0;
		2940: rom = 1'b0;
		2941: rom = 1'b0;
		2942: rom = 1'b0;
		2943: rom = 1'b0;
		2944: rom = 1'b0;
		2945: rom = 1'b0;
		2946: rom = 1'b0;
		2947: rom = 1'b0;
		2948: rom = 1'b0;
		2949: rom = 1'b0;
		2950: rom = 1'b0;
		2951: rom = 1'b0;
		2952: rom = 1'b0;
		2953: rom = 1'b0;
		2954: rom = 1'b0;
		2955: rom = 1'b0;
		2956: rom = 1'b0;
		2957: rom = 1'b0;
		2958: rom = 1'b0;
		2959: rom = 1'b0;
		2960: rom = 1'b0;
		2961: rom = 1'b0;
		2962: rom = 1'b0;
		2963: rom = 1'b0;
		2964: rom = 1'b0;
		2965: rom = 1'b0;
		2966: rom = 1'b0;
		2967: rom = 1'b0;
		2968: rom = 1'b0;
		2969: rom = 1'b0;
		2970: rom = 1'b0;
		2971: rom = 1'b0;
		2972: rom = 1'b0;
		2973: rom = 1'b0;
		2974: rom = 1'b0;
		2975: rom = 1'b0;
		2976: rom = 1'b0;
		2977: rom = 1'b0;
		2978: rom = 1'b0;
		2979: rom = 1'b1;
		2980: rom = 1'b1;
		2981: rom = 1'b1;
		2982: rom = 1'b1;
		2983: rom = 1'b1;
		2984: rom = 1'b1;
		2985: rom = 1'b1;
		2986: rom = 1'b1;
		2987: rom = 1'b1;
		2988: rom = 1'b1;
		2989: rom = 1'b1;
		2990: rom = 1'b1;
		2991: rom = 1'b1;
		2992: rom = 1'b1;
		2993: rom = 1'b1;
		2994: rom = 1'b1;
		2995: rom = 1'b0;
		2996: rom = 1'b0;
		2997: rom = 1'b0;
		2998: rom = 1'b0;
		2999: rom = 1'b0;
		3000: rom = 1'b0;
		3001: rom = 1'b0;
		3002: rom = 1'b0;
		3003: rom = 1'b0;
		3004: rom = 1'b0;
		3005: rom = 1'b0;
		3006: rom = 1'b0;
		3007: rom = 1'b0;
		3008: rom = 1'b0;
		3009: rom = 1'b1;
		3010: rom = 1'b1;
		3011: rom = 1'b1;
		3012: rom = 1'b1;
		3013: rom = 1'b1;
		3014: rom = 1'b1;
		3015: rom = 1'b1;
		3016: rom = 1'b1;
		3017: rom = 1'b1;
		3018: rom = 1'b1;
		3019: rom = 1'b1;
		3020: rom = 1'b1;
		3021: rom = 1'b1;
		3022: rom = 1'b1;
		3023: rom = 1'b1;
		3024: rom = 1'b1;
		3025: rom = 1'b1;
		3026: rom = 1'b1;
		3027: rom = 1'b1;
		3028: rom = 1'b1;
		3029: rom = 1'b1;
		3030: rom = 1'b1;
		3031: rom = 1'b1;
		3032: rom = 1'b1;
		3033: rom = 1'b1;
		3034: rom = 1'b1;
		3035: rom = 1'b1;
		3036: rom = 1'b1;
		3037: rom = 1'b1;
		3038: rom = 1'b1;
		3039: rom = 1'b1;
		3040: rom = 1'b1;
		3041: rom = 1'b1;
		3042: rom = 1'b1;
		3043: rom = 1'b1;
		3044: rom = 1'b1;
		3045: rom = 1'b1;
		3046: rom = 1'b1;
		3047: rom = 1'b1;
		3048: rom = 1'b1;
		3049: rom = 1'b1;
		3050: rom = 1'b1;
		3051: rom = 1'b1;
		3052: rom = 1'b1;
		3053: rom = 1'b1;
		3054: rom = 1'b1;
		3055: rom = 1'b0;
		3056: rom = 1'b0;
		3057: rom = 1'b0;
		3058: rom = 1'b0;
		3059: rom = 1'b0;
		3060: rom = 1'b0;
		3061: rom = 1'b0;
		3062: rom = 1'b0;
		3063: rom = 1'b0;
		3064: rom = 1'b0;
		3065: rom = 1'b0;
		3066: rom = 1'b0;
		3067: rom = 1'b0;
		3068: rom = 1'b0;
		3069: rom = 1'b0;
		3070: rom = 1'b0;
		3071: rom = 1'b0;
		3072: rom = 1'b0;
		3073: rom = 1'b0;
		3074: rom = 1'b0;
		3075: rom = 1'b0;
		3076: rom = 1'b0;
		3077: rom = 1'b0;
		3078: rom = 1'b0;
		3079: rom = 1'b0;
		3080: rom = 1'b0;
		3081: rom = 1'b0;
		3082: rom = 1'b0;
		3083: rom = 1'b0;
		3084: rom = 1'b0;
		3085: rom = 1'b0;
		3086: rom = 1'b0;
		3087: rom = 1'b0;
		3088: rom = 1'b0;
		3089: rom = 1'b0;
		3090: rom = 1'b0;
		3091: rom = 1'b0;
		3092: rom = 1'b0;
		3093: rom = 1'b0;
		3094: rom = 1'b0;
		3095: rom = 1'b0;
		3096: rom = 1'b0;
		3097: rom = 1'b0;
		3098: rom = 1'b0;
		3099: rom = 1'b0;
		3100: rom = 1'b0;
		3101: rom = 1'b0;
		3102: rom = 1'b0;
		3103: rom = 1'b0;
		3104: rom = 1'b0;
		3105: rom = 1'b0;
		3106: rom = 1'b0;
		3107: rom = 1'b1;
		3108: rom = 1'b1;
		3109: rom = 1'b1;
		3110: rom = 1'b1;
		3111: rom = 1'b1;
		3112: rom = 1'b1;
		3113: rom = 1'b1;
		3114: rom = 1'b1;
		3115: rom = 1'b1;
		3116: rom = 1'b1;
		3117: rom = 1'b1;
		3118: rom = 1'b1;
		3119: rom = 1'b1;
		3120: rom = 1'b1;
		3121: rom = 1'b1;
		3122: rom = 1'b0;
		3123: rom = 1'b0;
		3124: rom = 1'b0;
		3125: rom = 1'b0;
		3126: rom = 1'b0;
		3127: rom = 1'b0;
		3128: rom = 1'b0;
		3129: rom = 1'b0;
		3130: rom = 1'b0;
		3131: rom = 1'b0;
		3132: rom = 1'b0;
		3133: rom = 1'b0;
		3134: rom = 1'b0;
		3135: rom = 1'b1;
		3136: rom = 1'b1;
		3137: rom = 1'b1;
		3138: rom = 1'b1;
		3139: rom = 1'b1;
		3140: rom = 1'b1;
		3141: rom = 1'b1;
		3142: rom = 1'b1;
		3143: rom = 1'b1;
		3144: rom = 1'b1;
		3145: rom = 1'b1;
		3146: rom = 1'b1;
		3147: rom = 1'b1;
		3148: rom = 1'b1;
		3149: rom = 1'b1;
		3150: rom = 1'b1;
		3151: rom = 1'b1;
		3152: rom = 1'b1;
		3153: rom = 1'b1;
		3154: rom = 1'b1;
		3155: rom = 1'b1;
		3156: rom = 1'b1;
		3157: rom = 1'b1;
		3158: rom = 1'b1;
		3159: rom = 1'b1;
		3160: rom = 1'b1;
		3161: rom = 1'b1;
		3162: rom = 1'b1;
		3163: rom = 1'b1;
		3164: rom = 1'b1;
		3165: rom = 1'b1;
		3166: rom = 1'b1;
		3167: rom = 1'b1;
		3168: rom = 1'b1;
		3169: rom = 1'b1;
		3170: rom = 1'b1;
		3171: rom = 1'b1;
		3172: rom = 1'b1;
		3173: rom = 1'b1;
		3174: rom = 1'b1;
		3175: rom = 1'b1;
		3176: rom = 1'b1;
		3177: rom = 1'b1;
		3178: rom = 1'b1;
		3179: rom = 1'b1;
		3180: rom = 1'b1;
		3181: rom = 1'b1;
		3182: rom = 1'b1;
		3183: rom = 1'b0;
		3184: rom = 1'b0;
		3185: rom = 1'b0;
		3186: rom = 1'b0;
		3187: rom = 1'b0;
		3188: rom = 1'b0;
		3189: rom = 1'b0;
		3190: rom = 1'b0;
		3191: rom = 1'b0;
		3192: rom = 1'b1;
		3193: rom = 1'b0;
		3194: rom = 1'b0;
		3195: rom = 1'b0;
		3196: rom = 1'b0;
		3197: rom = 1'b0;
		3198: rom = 1'b0;
		3199: rom = 1'b0;
		3200: rom = 1'b0;
		3201: rom = 1'b0;
		3202: rom = 1'b0;
		3203: rom = 1'b0;
		3204: rom = 1'b0;
		3205: rom = 1'b0;
		3206: rom = 1'b0;
		3207: rom = 1'b0;
		3208: rom = 1'b0;
		3209: rom = 1'b0;
		3210: rom = 1'b0;
		3211: rom = 1'b0;
		3212: rom = 1'b0;
		3213: rom = 1'b0;
		3214: rom = 1'b0;
		3215: rom = 1'b0;
		3216: rom = 1'b0;
		3217: rom = 1'b0;
		3218: rom = 1'b0;
		3219: rom = 1'b0;
		3220: rom = 1'b0;
		3221: rom = 1'b0;
		3222: rom = 1'b0;
		3223: rom = 1'b0;
		3224: rom = 1'b0;
		3225: rom = 1'b0;
		3226: rom = 1'b0;
		3227: rom = 1'b0;
		3228: rom = 1'b0;
		3229: rom = 1'b0;
		3230: rom = 1'b0;
		3231: rom = 1'b0;
		3232: rom = 1'b0;
		3233: rom = 1'b0;
		3234: rom = 1'b1;
		3235: rom = 1'b1;
		3236: rom = 1'b1;
		3237: rom = 1'b1;
		3238: rom = 1'b1;
		3239: rom = 1'b1;
		3240: rom = 1'b1;
		3241: rom = 1'b1;
		3242: rom = 1'b1;
		3243: rom = 1'b1;
		3244: rom = 1'b1;
		3245: rom = 1'b1;
		3246: rom = 1'b1;
		3247: rom = 1'b1;
		3248: rom = 1'b1;
		3249: rom = 1'b0;
		3250: rom = 1'b0;
		3251: rom = 1'b0;
		3252: rom = 1'b0;
		3253: rom = 1'b0;
		3254: rom = 1'b0;
		3255: rom = 1'b0;
		3256: rom = 1'b0;
		3257: rom = 1'b0;
		3258: rom = 1'b0;
		3259: rom = 1'b0;
		3260: rom = 1'b0;
		3261: rom = 1'b0;
		3262: rom = 1'b1;
		3263: rom = 1'b1;
		3264: rom = 1'b1;
		3265: rom = 1'b1;
		3266: rom = 1'b1;
		3267: rom = 1'b1;
		3268: rom = 1'b1;
		3269: rom = 1'b1;
		3270: rom = 1'b1;
		3271: rom = 1'b1;
		3272: rom = 1'b1;
		3273: rom = 1'b1;
		3274: rom = 1'b1;
		3275: rom = 1'b1;
		3276: rom = 1'b1;
		3277: rom = 1'b1;
		3278: rom = 1'b1;
		3279: rom = 1'b1;
		3280: rom = 1'b1;
		3281: rom = 1'b1;
		3282: rom = 1'b1;
		3283: rom = 1'b1;
		3284: rom = 1'b1;
		3285: rom = 1'b1;
		3286: rom = 1'b1;
		3287: rom = 1'b1;
		3288: rom = 1'b1;
		3289: rom = 1'b1;
		3290: rom = 1'b1;
		3291: rom = 1'b1;
		3292: rom = 1'b1;
		3293: rom = 1'b1;
		3294: rom = 1'b1;
		3295: rom = 1'b1;
		3296: rom = 1'b1;
		3297: rom = 1'b1;
		3298: rom = 1'b1;
		3299: rom = 1'b1;
		3300: rom = 1'b1;
		3301: rom = 1'b1;
		3302: rom = 1'b1;
		3303: rom = 1'b1;
		3304: rom = 1'b1;
		3305: rom = 1'b1;
		3306: rom = 1'b1;
		3307: rom = 1'b1;
		3308: rom = 1'b1;
		3309: rom = 1'b1;
		3310: rom = 1'b1;
		3311: rom = 1'b1;
		3312: rom = 1'b0;
		3313: rom = 1'b0;
		3314: rom = 1'b0;
		3315: rom = 1'b0;
		3316: rom = 1'b0;
		3317: rom = 1'b0;
		3318: rom = 1'b0;
		3319: rom = 1'b0;
		3320: rom = 1'b1;
		3321: rom = 1'b0;
		3322: rom = 1'b0;
		3323: rom = 1'b0;
		3324: rom = 1'b0;
		3325: rom = 1'b0;
		3326: rom = 1'b0;
		3327: rom = 1'b0;
		3328: rom = 1'b0;
		3329: rom = 1'b0;
		3330: rom = 1'b0;
		3331: rom = 1'b0;
		3332: rom = 1'b0;
		3333: rom = 1'b0;
		3334: rom = 1'b0;
		3335: rom = 1'b0;
		3336: rom = 1'b0;
		3337: rom = 1'b0;
		3338: rom = 1'b0;
		3339: rom = 1'b0;
		3340: rom = 1'b0;
		3341: rom = 1'b0;
		3342: rom = 1'b0;
		3343: rom = 1'b0;
		3344: rom = 1'b0;
		3345: rom = 1'b0;
		3346: rom = 1'b0;
		3347: rom = 1'b0;
		3348: rom = 1'b0;
		3349: rom = 1'b0;
		3350: rom = 1'b0;
		3351: rom = 1'b0;
		3352: rom = 1'b0;
		3353: rom = 1'b0;
		3354: rom = 1'b0;
		3355: rom = 1'b0;
		3356: rom = 1'b0;
		3357: rom = 1'b0;
		3358: rom = 1'b0;
		3359: rom = 1'b0;
		3360: rom = 1'b0;
		3361: rom = 1'b0;
		3362: rom = 1'b1;
		3363: rom = 1'b1;
		3364: rom = 1'b1;
		3365: rom = 1'b1;
		3366: rom = 1'b1;
		3367: rom = 1'b1;
		3368: rom = 1'b1;
		3369: rom = 1'b1;
		3370: rom = 1'b1;
		3371: rom = 1'b1;
		3372: rom = 1'b1;
		3373: rom = 1'b1;
		3374: rom = 1'b1;
		3375: rom = 1'b1;
		3376: rom = 1'b0;
		3377: rom = 1'b0;
		3378: rom = 1'b0;
		3379: rom = 1'b0;
		3380: rom = 1'b0;
		3381: rom = 1'b0;
		3382: rom = 1'b0;
		3383: rom = 1'b0;
		3384: rom = 1'b0;
		3385: rom = 1'b0;
		3386: rom = 1'b0;
		3387: rom = 1'b0;
		3388: rom = 1'b0;
		3389: rom = 1'b1;
		3390: rom = 1'b1;
		3391: rom = 1'b1;
		3392: rom = 1'b1;
		3393: rom = 1'b1;
		3394: rom = 1'b1;
		3395: rom = 1'b1;
		3396: rom = 1'b1;
		3397: rom = 1'b1;
		3398: rom = 1'b1;
		3399: rom = 1'b1;
		3400: rom = 1'b1;
		3401: rom = 1'b1;
		3402: rom = 1'b1;
		3403: rom = 1'b1;
		3404: rom = 1'b1;
		3405: rom = 1'b1;
		3406: rom = 1'b1;
		3407: rom = 1'b1;
		3408: rom = 1'b1;
		3409: rom = 1'b1;
		3410: rom = 1'b1;
		3411: rom = 1'b1;
		3412: rom = 1'b1;
		3413: rom = 1'b1;
		3414: rom = 1'b1;
		3415: rom = 1'b1;
		3416: rom = 1'b1;
		3417: rom = 1'b1;
		3418: rom = 1'b1;
		3419: rom = 1'b1;
		3420: rom = 1'b1;
		3421: rom = 1'b1;
		3422: rom = 1'b1;
		3423: rom = 1'b1;
		3424: rom = 1'b1;
		3425: rom = 1'b1;
		3426: rom = 1'b1;
		3427: rom = 1'b1;
		3428: rom = 1'b1;
		3429: rom = 1'b1;
		3430: rom = 1'b1;
		3431: rom = 1'b1;
		3432: rom = 1'b1;
		3433: rom = 1'b1;
		3434: rom = 1'b1;
		3435: rom = 1'b1;
		3436: rom = 1'b1;
		3437: rom = 1'b1;
		3438: rom = 1'b1;
		3439: rom = 1'b1;
		3440: rom = 1'b0;
		3441: rom = 1'b0;
		3442: rom = 1'b0;
		3443: rom = 1'b0;
		3444: rom = 1'b0;
		3445: rom = 1'b0;
		3446: rom = 1'b0;
		3447: rom = 1'b1;
		3448: rom = 1'b1;
		3449: rom = 1'b0;
		3450: rom = 1'b0;
		3451: rom = 1'b0;
		3452: rom = 1'b0;
		3453: rom = 1'b0;
		3454: rom = 1'b0;
		3455: rom = 1'b0;
		3456: rom = 1'b0;
		3457: rom = 1'b0;
		3458: rom = 1'b0;
		3459: rom = 1'b0;
		3460: rom = 1'b0;
		3461: rom = 1'b0;
		3462: rom = 1'b0;
		3463: rom = 1'b0;
		3464: rom = 1'b0;
		3465: rom = 1'b0;
		3466: rom = 1'b0;
		3467: rom = 1'b0;
		3468: rom = 1'b0;
		3469: rom = 1'b0;
		3470: rom = 1'b0;
		3471: rom = 1'b0;
		3472: rom = 1'b0;
		3473: rom = 1'b0;
		3474: rom = 1'b0;
		3475: rom = 1'b0;
		3476: rom = 1'b0;
		3477: rom = 1'b0;
		3478: rom = 1'b0;
		3479: rom = 1'b0;
		3480: rom = 1'b0;
		3481: rom = 1'b0;
		3482: rom = 1'b0;
		3483: rom = 1'b0;
		3484: rom = 1'b0;
		3485: rom = 1'b0;
		3486: rom = 1'b0;
		3487: rom = 1'b0;
		3488: rom = 1'b0;
		3489: rom = 1'b1;
		3490: rom = 1'b1;
		3491: rom = 1'b1;
		3492: rom = 1'b1;
		3493: rom = 1'b1;
		3494: rom = 1'b1;
		3495: rom = 1'b1;
		3496: rom = 1'b1;
		3497: rom = 1'b1;
		3498: rom = 1'b1;
		3499: rom = 1'b1;
		3500: rom = 1'b1;
		3501: rom = 1'b1;
		3502: rom = 1'b1;
		3503: rom = 1'b0;
		3504: rom = 1'b0;
		3505: rom = 1'b0;
		3506: rom = 1'b0;
		3507: rom = 1'b0;
		3508: rom = 1'b0;
		3509: rom = 1'b0;
		3510: rom = 1'b0;
		3511: rom = 1'b0;
		3512: rom = 1'b0;
		3513: rom = 1'b0;
		3514: rom = 1'b0;
		3515: rom = 1'b1;
		3516: rom = 1'b1;
		3517: rom = 1'b1;
		3518: rom = 1'b1;
		3519: rom = 1'b1;
		3520: rom = 1'b1;
		3521: rom = 1'b1;
		3522: rom = 1'b1;
		3523: rom = 1'b1;
		3524: rom = 1'b1;
		3525: rom = 1'b1;
		3526: rom = 1'b1;
		3527: rom = 1'b1;
		3528: rom = 1'b0;
		3529: rom = 1'b0;
		3530: rom = 1'b1;
		3531: rom = 1'b1;
		3532: rom = 1'b1;
		3533: rom = 1'b1;
		3534: rom = 1'b1;
		3535: rom = 1'b1;
		3536: rom = 1'b1;
		3537: rom = 1'b1;
		3538: rom = 1'b1;
		3539: rom = 1'b1;
		3540: rom = 1'b1;
		3541: rom = 1'b1;
		3542: rom = 1'b1;
		3543: rom = 1'b1;
		3544: rom = 1'b1;
		3545: rom = 1'b1;
		3546: rom = 1'b0;
		3547: rom = 1'b1;
		3548: rom = 1'b1;
		3549: rom = 1'b1;
		3550: rom = 1'b1;
		3551: rom = 1'b1;
		3552: rom = 1'b1;
		3553: rom = 1'b1;
		3554: rom = 1'b1;
		3555: rom = 1'b1;
		3556: rom = 1'b1;
		3557: rom = 1'b1;
		3558: rom = 1'b1;
		3559: rom = 1'b1;
		3560: rom = 1'b1;
		3561: rom = 1'b1;
		3562: rom = 1'b1;
		3563: rom = 1'b1;
		3564: rom = 1'b1;
		3565: rom = 1'b1;
		3566: rom = 1'b1;
		3567: rom = 1'b1;
		3568: rom = 1'b1;
		3569: rom = 1'b0;
		3570: rom = 1'b0;
		3571: rom = 1'b0;
		3572: rom = 1'b0;
		3573: rom = 1'b0;
		3574: rom = 1'b0;
		3575: rom = 1'b1;
		3576: rom = 1'b1;
		3577: rom = 1'b0;
		3578: rom = 1'b0;
		3579: rom = 1'b0;
		3580: rom = 1'b0;
		3581: rom = 1'b0;
		3582: rom = 1'b0;
		3583: rom = 1'b0;
		3584: rom = 1'b0;
		3585: rom = 1'b0;
		3586: rom = 1'b0;
		3587: rom = 1'b0;
		3588: rom = 1'b0;
		3589: rom = 1'b0;
		3590: rom = 1'b0;
		3591: rom = 1'b0;
		3592: rom = 1'b0;
		3593: rom = 1'b0;
		3594: rom = 1'b0;
		3595: rom = 1'b0;
		3596: rom = 1'b0;
		3597: rom = 1'b0;
		3598: rom = 1'b0;
		3599: rom = 1'b0;
		3600: rom = 1'b0;
		3601: rom = 1'b0;
		3602: rom = 1'b0;
		3603: rom = 1'b0;
		3604: rom = 1'b0;
		3605: rom = 1'b0;
		3606: rom = 1'b0;
		3607: rom = 1'b0;
		3608: rom = 1'b0;
		3609: rom = 1'b0;
		3610: rom = 1'b0;
		3611: rom = 1'b0;
		3612: rom = 1'b0;
		3613: rom = 1'b0;
		3614: rom = 1'b0;
		3615: rom = 1'b0;
		3616: rom = 1'b1;
		3617: rom = 1'b1;
		3618: rom = 1'b1;
		3619: rom = 1'b1;
		3620: rom = 1'b1;
		3621: rom = 1'b1;
		3622: rom = 1'b1;
		3623: rom = 1'b1;
		3624: rom = 1'b1;
		3625: rom = 1'b1;
		3626: rom = 1'b1;
		3627: rom = 1'b1;
		3628: rom = 1'b1;
		3629: rom = 1'b1;
		3630: rom = 1'b0;
		3631: rom = 1'b0;
		3632: rom = 1'b0;
		3633: rom = 1'b0;
		3634: rom = 1'b0;
		3635: rom = 1'b0;
		3636: rom = 1'b0;
		3637: rom = 1'b0;
		3638: rom = 1'b0;
		3639: rom = 1'b0;
		3640: rom = 1'b0;
		3641: rom = 1'b0;
		3642: rom = 1'b1;
		3643: rom = 1'b1;
		3644: rom = 1'b1;
		3645: rom = 1'b1;
		3646: rom = 1'b1;
		3647: rom = 1'b1;
		3648: rom = 1'b1;
		3649: rom = 1'b1;
		3650: rom = 1'b1;
		3651: rom = 1'b1;
		3652: rom = 1'b1;
		3653: rom = 1'b1;
		3654: rom = 1'b1;
		3655: rom = 1'b1;
		3656: rom = 1'b0;
		3657: rom = 1'b0;
		3658: rom = 1'b0;
		3659: rom = 1'b1;
		3660: rom = 1'b1;
		3661: rom = 1'b1;
		3662: rom = 1'b1;
		3663: rom = 1'b1;
		3664: rom = 1'b1;
		3665: rom = 1'b1;
		3666: rom = 1'b1;
		3667: rom = 1'b1;
		3668: rom = 1'b1;
		3669: rom = 1'b1;
		3670: rom = 1'b1;
		3671: rom = 1'b1;
		3672: rom = 1'b1;
		3673: rom = 1'b0;
		3674: rom = 1'b0;
		3675: rom = 1'b1;
		3676: rom = 1'b1;
		3677: rom = 1'b1;
		3678: rom = 1'b1;
		3679: rom = 1'b1;
		3680: rom = 1'b1;
		3681: rom = 1'b1;
		3682: rom = 1'b1;
		3683: rom = 1'b1;
		3684: rom = 1'b1;
		3685: rom = 1'b1;
		3686: rom = 1'b1;
		3687: rom = 1'b1;
		3688: rom = 1'b1;
		3689: rom = 1'b1;
		3690: rom = 1'b1;
		3691: rom = 1'b1;
		3692: rom = 1'b1;
		3693: rom = 1'b1;
		3694: rom = 1'b1;
		3695: rom = 1'b1;
		3696: rom = 1'b1;
		3697: rom = 1'b1;
		3698: rom = 1'b0;
		3699: rom = 1'b0;
		3700: rom = 1'b0;
		3701: rom = 1'b0;
		3702: rom = 1'b0;
		3703: rom = 1'b1;
		3704: rom = 1'b0;
		3705: rom = 1'b0;
		3706: rom = 1'b0;
		3707: rom = 1'b0;
		3708: rom = 1'b0;
		3709: rom = 1'b0;
		3710: rom = 1'b0;
		3711: rom = 1'b0;
		3712: rom = 1'b0;
		3713: rom = 1'b0;
		3714: rom = 1'b0;
		3715: rom = 1'b0;
		3716: rom = 1'b0;
		3717: rom = 1'b0;
		3718: rom = 1'b0;
		3719: rom = 1'b0;
		3720: rom = 1'b0;
		3721: rom = 1'b0;
		3722: rom = 1'b0;
		3723: rom = 1'b0;
		3724: rom = 1'b0;
		3725: rom = 1'b0;
		3726: rom = 1'b0;
		3727: rom = 1'b0;
		3728: rom = 1'b0;
		3729: rom = 1'b0;
		3730: rom = 1'b0;
		3731: rom = 1'b0;
		3732: rom = 1'b0;
		3733: rom = 1'b0;
		3734: rom = 1'b0;
		3735: rom = 1'b0;
		3736: rom = 1'b0;
		3737: rom = 1'b0;
		3738: rom = 1'b0;
		3739: rom = 1'b0;
		3740: rom = 1'b0;
		3741: rom = 1'b0;
		3742: rom = 1'b0;
		3743: rom = 1'b0;
		3744: rom = 1'b1;
		3745: rom = 1'b1;
		3746: rom = 1'b1;
		3747: rom = 1'b1;
		3748: rom = 1'b1;
		3749: rom = 1'b1;
		3750: rom = 1'b1;
		3751: rom = 1'b1;
		3752: rom = 1'b1;
		3753: rom = 1'b1;
		3754: rom = 1'b1;
		3755: rom = 1'b1;
		3756: rom = 1'b1;
		3757: rom = 1'b0;
		3758: rom = 1'b0;
		3759: rom = 1'b0;
		3760: rom = 1'b0;
		3761: rom = 1'b0;
		3762: rom = 1'b0;
		3763: rom = 1'b0;
		3764: rom = 1'b0;
		3765: rom = 1'b0;
		3766: rom = 1'b0;
		3767: rom = 1'b0;
		3768: rom = 1'b0;
		3769: rom = 1'b1;
		3770: rom = 1'b1;
		3771: rom = 1'b1;
		3772: rom = 1'b1;
		3773: rom = 1'b1;
		3774: rom = 1'b1;
		3775: rom = 1'b1;
		3776: rom = 1'b1;
		3777: rom = 1'b1;
		3778: rom = 1'b1;
		3779: rom = 1'b1;
		3780: rom = 1'b1;
		3781: rom = 1'b1;
		3782: rom = 1'b1;
		3783: rom = 1'b1;
		3784: rom = 1'b0;
		3785: rom = 1'b0;
		3786: rom = 1'b0;
		3787: rom = 1'b1;
		3788: rom = 1'b1;
		3789: rom = 1'b1;
		3790: rom = 1'b1;
		3791: rom = 1'b1;
		3792: rom = 1'b1;
		3793: rom = 1'b1;
		3794: rom = 1'b1;
		3795: rom = 1'b1;
		3796: rom = 1'b1;
		3797: rom = 1'b1;
		3798: rom = 1'b1;
		3799: rom = 1'b1;
		3800: rom = 1'b1;
		3801: rom = 1'b0;
		3802: rom = 1'b0;
		3803: rom = 1'b0;
		3804: rom = 1'b1;
		3805: rom = 1'b1;
		3806: rom = 1'b1;
		3807: rom = 1'b1;
		3808: rom = 1'b1;
		3809: rom = 1'b1;
		3810: rom = 1'b1;
		3811: rom = 1'b1;
		3812: rom = 1'b1;
		3813: rom = 1'b1;
		3814: rom = 1'b1;
		3815: rom = 1'b1;
		3816: rom = 1'b1;
		3817: rom = 1'b1;
		3818: rom = 1'b1;
		3819: rom = 1'b1;
		3820: rom = 1'b1;
		3821: rom = 1'b1;
		3822: rom = 1'b1;
		3823: rom = 1'b1;
		3824: rom = 1'b1;
		3825: rom = 1'b1;
		3826: rom = 1'b0;
		3827: rom = 1'b0;
		3828: rom = 1'b0;
		3829: rom = 1'b0;
		3830: rom = 1'b1;
		3831: rom = 1'b1;
		3832: rom = 1'b0;
		3833: rom = 1'b0;
		3834: rom = 1'b0;
		3835: rom = 1'b0;
		3836: rom = 1'b0;
		3837: rom = 1'b0;
		3838: rom = 1'b0;
		3839: rom = 1'b0;
		3840: rom = 1'b0;
		3841: rom = 1'b0;
		3842: rom = 1'b0;
		3843: rom = 1'b0;
		3844: rom = 1'b0;
		3845: rom = 1'b0;
		3846: rom = 1'b0;
		3847: rom = 1'b0;
		3848: rom = 1'b0;
		3849: rom = 1'b0;
		3850: rom = 1'b0;
		3851: rom = 1'b0;
		3852: rom = 1'b0;
		3853: rom = 1'b0;
		3854: rom = 1'b0;
		3855: rom = 1'b0;
		3856: rom = 1'b0;
		3857: rom = 1'b0;
		3858: rom = 1'b0;
		3859: rom = 1'b0;
		3860: rom = 1'b0;
		3861: rom = 1'b0;
		3862: rom = 1'b0;
		3863: rom = 1'b0;
		3864: rom = 1'b0;
		3865: rom = 1'b0;
		3866: rom = 1'b0;
		3867: rom = 1'b0;
		3868: rom = 1'b0;
		3869: rom = 1'b0;
		3870: rom = 1'b0;
		3871: rom = 1'b0;
		3872: rom = 1'b1;
		3873: rom = 1'b1;
		3874: rom = 1'b1;
		3875: rom = 1'b1;
		3876: rom = 1'b1;
		3877: rom = 1'b1;
		3878: rom = 1'b1;
		3879: rom = 1'b1;
		3880: rom = 1'b1;
		3881: rom = 1'b1;
		3882: rom = 1'b1;
		3883: rom = 1'b1;
		3884: rom = 1'b0;
		3885: rom = 1'b0;
		3886: rom = 1'b0;
		3887: rom = 1'b0;
		3888: rom = 1'b0;
		3889: rom = 1'b0;
		3890: rom = 1'b0;
		3891: rom = 1'b0;
		3892: rom = 1'b0;
		3893: rom = 1'b0;
		3894: rom = 1'b0;
		3895: rom = 1'b0;
		3896: rom = 1'b1;
		3897: rom = 1'b1;
		3898: rom = 1'b1;
		3899: rom = 1'b1;
		3900: rom = 1'b1;
		3901: rom = 1'b1;
		3902: rom = 1'b1;
		3903: rom = 1'b1;
		3904: rom = 1'b1;
		3905: rom = 1'b1;
		3906: rom = 1'b1;
		3907: rom = 1'b1;
		3908: rom = 1'b1;
		3909: rom = 1'b1;
		3910: rom = 1'b1;
		3911: rom = 1'b0;
		3912: rom = 1'b0;
		3913: rom = 1'b0;
		3914: rom = 1'b0;
		3915: rom = 1'b0;
		3916: rom = 1'b1;
		3917: rom = 1'b1;
		3918: rom = 1'b1;
		3919: rom = 1'b1;
		3920: rom = 1'b1;
		3921: rom = 1'b1;
		3922: rom = 1'b1;
		3923: rom = 1'b1;
		3924: rom = 1'b1;
		3925: rom = 1'b1;
		3926: rom = 1'b1;
		3927: rom = 1'b0;
		3928: rom = 1'b0;
		3929: rom = 1'b0;
		3930: rom = 1'b0;
		3931: rom = 1'b0;
		3932: rom = 1'b0;
		3933: rom = 1'b1;
		3934: rom = 1'b1;
		3935: rom = 1'b1;
		3936: rom = 1'b1;
		3937: rom = 1'b1;
		3938: rom = 1'b1;
		3939: rom = 1'b1;
		3940: rom = 1'b1;
		3941: rom = 1'b1;
		3942: rom = 1'b1;
		3943: rom = 1'b1;
		3944: rom = 1'b1;
		3945: rom = 1'b1;
		3946: rom = 1'b1;
		3947: rom = 1'b1;
		3948: rom = 1'b1;
		3949: rom = 1'b1;
		3950: rom = 1'b1;
		3951: rom = 1'b1;
		3952: rom = 1'b1;
		3953: rom = 1'b1;
		3954: rom = 1'b1;
		3955: rom = 1'b0;
		3956: rom = 1'b0;
		3957: rom = 1'b0;
		3958: rom = 1'b1;
		3959: rom = 1'b1;
		3960: rom = 1'b0;
		3961: rom = 1'b0;
		3962: rom = 1'b0;
		3963: rom = 1'b0;
		3964: rom = 1'b0;
		3965: rom = 1'b0;
		3966: rom = 1'b0;
		3967: rom = 1'b0;
		3968: rom = 1'b0;
		3969: rom = 1'b0;
		3970: rom = 1'b0;
		3971: rom = 1'b0;
		3972: rom = 1'b0;
		3973: rom = 1'b0;
		3974: rom = 1'b0;
		3975: rom = 1'b0;
		3976: rom = 1'b0;
		3977: rom = 1'b0;
		3978: rom = 1'b0;
		3979: rom = 1'b0;
		3980: rom = 1'b0;
		3981: rom = 1'b0;
		3982: rom = 1'b0;
		3983: rom = 1'b0;
		3984: rom = 1'b0;
		3985: rom = 1'b0;
		3986: rom = 1'b0;
		3987: rom = 1'b0;
		3988: rom = 1'b0;
		3989: rom = 1'b0;
		3990: rom = 1'b0;
		3991: rom = 1'b0;
		3992: rom = 1'b0;
		3993: rom = 1'b0;
		3994: rom = 1'b0;
		3995: rom = 1'b0;
		3996: rom = 1'b0;
		3997: rom = 1'b0;
		3998: rom = 1'b0;
		3999: rom = 1'b1;
		4000: rom = 1'b1;
		4001: rom = 1'b1;
		4002: rom = 1'b1;
		4003: rom = 1'b1;
		4004: rom = 1'b1;
		4005: rom = 1'b1;
		4006: rom = 1'b1;
		4007: rom = 1'b1;
		4008: rom = 1'b1;
		4009: rom = 1'b1;
		4010: rom = 1'b1;
		4011: rom = 1'b0;
		4012: rom = 1'b0;
		4013: rom = 1'b0;
		4014: rom = 1'b0;
		4015: rom = 1'b0;
		4016: rom = 1'b0;
		4017: rom = 1'b0;
		4018: rom = 1'b0;
		4019: rom = 1'b0;
		4020: rom = 1'b0;
		4021: rom = 1'b0;
		4022: rom = 1'b0;
		4023: rom = 1'b1;
		4024: rom = 1'b1;
		4025: rom = 1'b1;
		4026: rom = 1'b1;
		4027: rom = 1'b1;
		4028: rom = 1'b1;
		4029: rom = 1'b1;
		4030: rom = 1'b1;
		4031: rom = 1'b1;
		4032: rom = 1'b1;
		4033: rom = 1'b1;
		4034: rom = 1'b1;
		4035: rom = 1'b1;
		4036: rom = 1'b1;
		4037: rom = 1'b0;
		4038: rom = 1'b0;
		4039: rom = 1'b0;
		4040: rom = 1'b0;
		4041: rom = 1'b0;
		4042: rom = 1'b0;
		4043: rom = 1'b0;
		4044: rom = 1'b0;
		4045: rom = 1'b0;
		4046: rom = 1'b1;
		4047: rom = 1'b1;
		4048: rom = 1'b1;
		4049: rom = 1'b1;
		4050: rom = 1'b1;
		4051: rom = 1'b1;
		4052: rom = 1'b1;
		4053: rom = 1'b1;
		4054: rom = 1'b1;
		4055: rom = 1'b0;
		4056: rom = 1'b0;
		4057: rom = 1'b0;
		4058: rom = 1'b0;
		4059: rom = 1'b0;
		4060: rom = 1'b0;
		4061: rom = 1'b1;
		4062: rom = 1'b1;
		4063: rom = 1'b1;
		4064: rom = 1'b1;
		4065: rom = 1'b1;
		4066: rom = 1'b1;
		4067: rom = 1'b1;
		4068: rom = 1'b1;
		4069: rom = 1'b1;
		4070: rom = 1'b1;
		4071: rom = 1'b1;
		4072: rom = 1'b1;
		4073: rom = 1'b1;
		4074: rom = 1'b1;
		4075: rom = 1'b1;
		4076: rom = 1'b1;
		4077: rom = 1'b1;
		4078: rom = 1'b1;
		4079: rom = 1'b1;
		4080: rom = 1'b1;
		4081: rom = 1'b1;
		4082: rom = 1'b1;
		4083: rom = 1'b0;
		4084: rom = 1'b0;
		4085: rom = 1'b1;
		4086: rom = 1'b1;
		4087: rom = 1'b1;
		4088: rom = 1'b0;
		4089: rom = 1'b0;
		4090: rom = 1'b0;
		4091: rom = 1'b0;
		4092: rom = 1'b0;
		4093: rom = 1'b0;
		4094: rom = 1'b0;
		4095: rom = 1'b0;
		4096: rom = 1'b0;
		4097: rom = 1'b0;
		4098: rom = 1'b0;
		4099: rom = 1'b0;
		4100: rom = 1'b0;
		4101: rom = 1'b0;
		4102: rom = 1'b0;
		4103: rom = 1'b0;
		4104: rom = 1'b0;
		4105: rom = 1'b0;
		4106: rom = 1'b0;
		4107: rom = 1'b0;
		4108: rom = 1'b0;
		4109: rom = 1'b0;
		4110: rom = 1'b0;
		4111: rom = 1'b0;
		4112: rom = 1'b0;
		4113: rom = 1'b0;
		4114: rom = 1'b0;
		4115: rom = 1'b0;
		4116: rom = 1'b0;
		4117: rom = 1'b0;
		4118: rom = 1'b0;
		4119: rom = 1'b0;
		4120: rom = 1'b0;
		4121: rom = 1'b0;
		4122: rom = 1'b0;
		4123: rom = 1'b0;
		4124: rom = 1'b0;
		4125: rom = 1'b0;
		4126: rom = 1'b0;
		4127: rom = 1'b1;
		4128: rom = 1'b1;
		4129: rom = 1'b1;
		4130: rom = 1'b1;
		4131: rom = 1'b1;
		4132: rom = 1'b1;
		4133: rom = 1'b1;
		4134: rom = 1'b1;
		4135: rom = 1'b1;
		4136: rom = 1'b1;
		4137: rom = 1'b1;
		4138: rom = 1'b0;
		4139: rom = 1'b0;
		4140: rom = 1'b0;
		4141: rom = 1'b0;
		4142: rom = 1'b0;
		4143: rom = 1'b0;
		4144: rom = 1'b0;
		4145: rom = 1'b0;
		4146: rom = 1'b0;
		4147: rom = 1'b0;
		4148: rom = 1'b0;
		4149: rom = 1'b0;
		4150: rom = 1'b1;
		4151: rom = 1'b1;
		4152: rom = 1'b1;
		4153: rom = 1'b1;
		4154: rom = 1'b1;
		4155: rom = 1'b1;
		4156: rom = 1'b1;
		4157: rom = 1'b1;
		4158: rom = 1'b1;
		4159: rom = 1'b1;
		4160: rom = 1'b1;
		4161: rom = 1'b1;
		4162: rom = 1'b1;
		4163: rom = 1'b0;
		4164: rom = 1'b0;
		4165: rom = 1'b0;
		4166: rom = 1'b0;
		4167: rom = 1'b0;
		4168: rom = 1'b0;
		4169: rom = 1'b0;
		4170: rom = 1'b0;
		4171: rom = 1'b0;
		4172: rom = 1'b0;
		4173: rom = 1'b0;
		4174: rom = 1'b0;
		4175: rom = 1'b1;
		4176: rom = 1'b1;
		4177: rom = 1'b1;
		4178: rom = 1'b1;
		4179: rom = 1'b1;
		4180: rom = 1'b1;
		4181: rom = 1'b1;
		4182: rom = 1'b1;
		4183: rom = 1'b1;
		4184: rom = 1'b1;
		4185: rom = 1'b0;
		4186: rom = 1'b0;
		4187: rom = 1'b1;
		4188: rom = 1'b1;
		4189: rom = 1'b1;
		4190: rom = 1'b1;
		4191: rom = 1'b1;
		4192: rom = 1'b1;
		4193: rom = 1'b1;
		4194: rom = 1'b1;
		4195: rom = 1'b1;
		4196: rom = 1'b1;
		4197: rom = 1'b1;
		4198: rom = 1'b1;
		4199: rom = 1'b1;
		4200: rom = 1'b1;
		4201: rom = 1'b1;
		4202: rom = 1'b1;
		4203: rom = 1'b1;
		4204: rom = 1'b1;
		4205: rom = 1'b1;
		4206: rom = 1'b1;
		4207: rom = 1'b1;
		4208: rom = 1'b1;
		4209: rom = 1'b1;
		4210: rom = 1'b1;
		4211: rom = 1'b1;
		4212: rom = 1'b0;
		4213: rom = 1'b1;
		4214: rom = 1'b1;
		4215: rom = 1'b1;
		4216: rom = 1'b0;
		4217: rom = 1'b0;
		4218: rom = 1'b0;
		4219: rom = 1'b0;
		4220: rom = 1'b0;
		4221: rom = 1'b0;
		4222: rom = 1'b0;
		4223: rom = 1'b0;
		4224: rom = 1'b0;
		4225: rom = 1'b0;
		4226: rom = 1'b0;
		4227: rom = 1'b0;
		4228: rom = 1'b0;
		4229: rom = 1'b0;
		4230: rom = 1'b0;
		4231: rom = 1'b0;
		4232: rom = 1'b0;
		4233: rom = 1'b0;
		4234: rom = 1'b0;
		4235: rom = 1'b0;
		4236: rom = 1'b0;
		4237: rom = 1'b0;
		4238: rom = 1'b0;
		4239: rom = 1'b0;
		4240: rom = 1'b0;
		4241: rom = 1'b0;
		4242: rom = 1'b0;
		4243: rom = 1'b0;
		4244: rom = 1'b0;
		4245: rom = 1'b0;
		4246: rom = 1'b0;
		4247: rom = 1'b0;
		4248: rom = 1'b0;
		4249: rom = 1'b0;
		4250: rom = 1'b0;
		4251: rom = 1'b0;
		4252: rom = 1'b0;
		4253: rom = 1'b0;
		4254: rom = 1'b1;
		4255: rom = 1'b1;
		4256: rom = 1'b1;
		4257: rom = 1'b1;
		4258: rom = 1'b1;
		4259: rom = 1'b1;
		4260: rom = 1'b1;
		4261: rom = 1'b1;
		4262: rom = 1'b1;
		4263: rom = 1'b1;
		4264: rom = 1'b1;
		4265: rom = 1'b1;
		4266: rom = 1'b0;
		4267: rom = 1'b0;
		4268: rom = 1'b0;
		4269: rom = 1'b0;
		4270: rom = 1'b0;
		4271: rom = 1'b0;
		4272: rom = 1'b0;
		4273: rom = 1'b0;
		4274: rom = 1'b0;
		4275: rom = 1'b0;
		4276: rom = 1'b0;
		4277: rom = 1'b1;
		4278: rom = 1'b1;
		4279: rom = 1'b1;
		4280: rom = 1'b1;
		4281: rom = 1'b1;
		4282: rom = 1'b1;
		4283: rom = 1'b1;
		4284: rom = 1'b1;
		4285: rom = 1'b1;
		4286: rom = 1'b1;
		4287: rom = 1'b1;
		4288: rom = 1'b1;
		4289: rom = 1'b1;
		4290: rom = 1'b1;
		4291: rom = 1'b1;
		4292: rom = 1'b1;
		4293: rom = 1'b1;
		4294: rom = 1'b0;
		4295: rom = 1'b0;
		4296: rom = 1'b0;
		4297: rom = 1'b0;
		4298: rom = 1'b0;
		4299: rom = 1'b0;
		4300: rom = 1'b0;
		4301: rom = 1'b1;
		4302: rom = 1'b1;
		4303: rom = 1'b1;
		4304: rom = 1'b1;
		4305: rom = 1'b1;
		4306: rom = 1'b1;
		4307: rom = 1'b1;
		4308: rom = 1'b1;
		4309: rom = 1'b1;
		4310: rom = 1'b1;
		4311: rom = 1'b1;
		4312: rom = 1'b1;
		4313: rom = 1'b0;
		4314: rom = 1'b0;
		4315: rom = 1'b1;
		4316: rom = 1'b1;
		4317: rom = 1'b1;
		4318: rom = 1'b1;
		4319: rom = 1'b1;
		4320: rom = 1'b1;
		4321: rom = 1'b1;
		4322: rom = 1'b1;
		4323: rom = 1'b1;
		4324: rom = 1'b1;
		4325: rom = 1'b1;
		4326: rom = 1'b1;
		4327: rom = 1'b1;
		4328: rom = 1'b1;
		4329: rom = 1'b1;
		4330: rom = 1'b1;
		4331: rom = 1'b1;
		4332: rom = 1'b1;
		4333: rom = 1'b1;
		4334: rom = 1'b1;
		4335: rom = 1'b1;
		4336: rom = 1'b1;
		4337: rom = 1'b1;
		4338: rom = 1'b1;
		4339: rom = 1'b0;
		4340: rom = 1'b1;
		4341: rom = 1'b1;
		4342: rom = 1'b1;
		4343: rom = 1'b1;
		4344: rom = 1'b0;
		4345: rom = 1'b0;
		4346: rom = 1'b0;
		4347: rom = 1'b0;
		4348: rom = 1'b0;
		4349: rom = 1'b0;
		4350: rom = 1'b0;
		4351: rom = 1'b0;
		4352: rom = 1'b0;
		4353: rom = 1'b0;
		4354: rom = 1'b0;
		4355: rom = 1'b0;
		4356: rom = 1'b0;
		4357: rom = 1'b0;
		4358: rom = 1'b0;
		4359: rom = 1'b0;
		4360: rom = 1'b0;
		4361: rom = 1'b0;
		4362: rom = 1'b0;
		4363: rom = 1'b0;
		4364: rom = 1'b0;
		4365: rom = 1'b0;
		4366: rom = 1'b0;
		4367: rom = 1'b0;
		4368: rom = 1'b0;
		4369: rom = 1'b0;
		4370: rom = 1'b0;
		4371: rom = 1'b0;
		4372: rom = 1'b0;
		4373: rom = 1'b0;
		4374: rom = 1'b0;
		4375: rom = 1'b0;
		4376: rom = 1'b0;
		4377: rom = 1'b0;
		4378: rom = 1'b0;
		4379: rom = 1'b0;
		4380: rom = 1'b0;
		4381: rom = 1'b0;
		4382: rom = 1'b1;
		4383: rom = 1'b1;
		4384: rom = 1'b1;
		4385: rom = 1'b1;
		4386: rom = 1'b1;
		4387: rom = 1'b1;
		4388: rom = 1'b1;
		4389: rom = 1'b1;
		4390: rom = 1'b1;
		4391: rom = 1'b1;
		4392: rom = 1'b1;
		4393: rom = 1'b0;
		4394: rom = 1'b0;
		4395: rom = 1'b0;
		4396: rom = 1'b0;
		4397: rom = 1'b0;
		4398: rom = 1'b0;
		4399: rom = 1'b0;
		4400: rom = 1'b0;
		4401: rom = 1'b0;
		4402: rom = 1'b0;
		4403: rom = 1'b0;
		4404: rom = 1'b1;
		4405: rom = 1'b1;
		4406: rom = 1'b1;
		4407: rom = 1'b1;
		4408: rom = 1'b1;
		4409: rom = 1'b1;
		4410: rom = 1'b1;
		4411: rom = 1'b1;
		4412: rom = 1'b1;
		4413: rom = 1'b1;
		4414: rom = 1'b1;
		4415: rom = 1'b1;
		4416: rom = 1'b1;
		4417: rom = 1'b1;
		4418: rom = 1'b1;
		4419: rom = 1'b1;
		4420: rom = 1'b1;
		4421: rom = 1'b1;
		4422: rom = 1'b1;
		4423: rom = 1'b0;
		4424: rom = 1'b0;
		4425: rom = 1'b0;
		4426: rom = 1'b0;
		4427: rom = 1'b1;
		4428: rom = 1'b1;
		4429: rom = 1'b1;
		4430: rom = 1'b1;
		4431: rom = 1'b1;
		4432: rom = 1'b1;
		4433: rom = 1'b1;
		4434: rom = 1'b1;
		4435: rom = 1'b1;
		4436: rom = 1'b1;
		4437: rom = 1'b1;
		4438: rom = 1'b1;
		4439: rom = 1'b1;
		4440: rom = 1'b1;
		4441: rom = 1'b1;
		4442: rom = 1'b1;
		4443: rom = 1'b1;
		4444: rom = 1'b1;
		4445: rom = 1'b1;
		4446: rom = 1'b1;
		4447: rom = 1'b1;
		4448: rom = 1'b1;
		4449: rom = 1'b1;
		4450: rom = 1'b1;
		4451: rom = 1'b1;
		4452: rom = 1'b1;
		4453: rom = 1'b1;
		4454: rom = 1'b1;
		4455: rom = 1'b1;
		4456: rom = 1'b1;
		4457: rom = 1'b1;
		4458: rom = 1'b1;
		4459: rom = 1'b1;
		4460: rom = 1'b1;
		4461: rom = 1'b1;
		4462: rom = 1'b1;
		4463: rom = 1'b1;
		4464: rom = 1'b1;
		4465: rom = 1'b1;
		4466: rom = 1'b1;
		4467: rom = 1'b0;
		4468: rom = 1'b1;
		4469: rom = 1'b1;
		4470: rom = 1'b1;
		4471: rom = 1'b0;
		4472: rom = 1'b0;
		4473: rom = 1'b0;
		4474: rom = 1'b0;
		4475: rom = 1'b0;
		4476: rom = 1'b0;
		4477: rom = 1'b0;
		4478: rom = 1'b0;
		4479: rom = 1'b0;
		4480: rom = 1'b0;
		4481: rom = 1'b0;
		4482: rom = 1'b0;
		4483: rom = 1'b0;
		4484: rom = 1'b0;
		4485: rom = 1'b0;
		4486: rom = 1'b0;
		4487: rom = 1'b0;
		4488: rom = 1'b0;
		4489: rom = 1'b0;
		4490: rom = 1'b0;
		4491: rom = 1'b0;
		4492: rom = 1'b0;
		4493: rom = 1'b0;
		4494: rom = 1'b0;
		4495: rom = 1'b0;
		4496: rom = 1'b0;
		4497: rom = 1'b0;
		4498: rom = 1'b0;
		4499: rom = 1'b0;
		4500: rom = 1'b0;
		4501: rom = 1'b0;
		4502: rom = 1'b0;
		4503: rom = 1'b0;
		4504: rom = 1'b0;
		4505: rom = 1'b0;
		4506: rom = 1'b0;
		4507: rom = 1'b0;
		4508: rom = 1'b0;
		4509: rom = 1'b1;
		4510: rom = 1'b1;
		4511: rom = 1'b1;
		4512: rom = 1'b1;
		4513: rom = 1'b1;
		4514: rom = 1'b1;
		4515: rom = 1'b1;
		4516: rom = 1'b1;
		4517: rom = 1'b1;
		4518: rom = 1'b1;
		4519: rom = 1'b1;
		4520: rom = 1'b0;
		4521: rom = 1'b0;
		4522: rom = 1'b0;
		4523: rom = 1'b0;
		4524: rom = 1'b0;
		4525: rom = 1'b0;
		4526: rom = 1'b0;
		4527: rom = 1'b0;
		4528: rom = 1'b0;
		4529: rom = 1'b0;
		4530: rom = 1'b0;
		4531: rom = 1'b1;
		4532: rom = 1'b1;
		4533: rom = 1'b1;
		4534: rom = 1'b1;
		4535: rom = 1'b1;
		4536: rom = 1'b1;
		4537: rom = 1'b1;
		4538: rom = 1'b1;
		4539: rom = 1'b1;
		4540: rom = 1'b1;
		4541: rom = 1'b1;
		4542: rom = 1'b1;
		4543: rom = 1'b1;
		4544: rom = 1'b1;
		4545: rom = 1'b1;
		4546: rom = 1'b1;
		4547: rom = 1'b1;
		4548: rom = 1'b1;
		4549: rom = 1'b1;
		4550: rom = 1'b1;
		4551: rom = 1'b1;
		4552: rom = 1'b0;
		4553: rom = 1'b0;
		4554: rom = 1'b0;
		4555: rom = 1'b1;
		4556: rom = 1'b1;
		4557: rom = 1'b1;
		4558: rom = 1'b1;
		4559: rom = 1'b1;
		4560: rom = 1'b1;
		4561: rom = 1'b1;
		4562: rom = 1'b1;
		4563: rom = 1'b1;
		4564: rom = 1'b1;
		4565: rom = 1'b1;
		4566: rom = 1'b1;
		4567: rom = 1'b1;
		4568: rom = 1'b1;
		4569: rom = 1'b1;
		4570: rom = 1'b1;
		4571: rom = 1'b1;
		4572: rom = 1'b1;
		4573: rom = 1'b1;
		4574: rom = 1'b1;
		4575: rom = 1'b1;
		4576: rom = 1'b1;
		4577: rom = 1'b1;
		4578: rom = 1'b1;
		4579: rom = 1'b1;
		4580: rom = 1'b1;
		4581: rom = 1'b1;
		4582: rom = 1'b1;
		4583: rom = 1'b1;
		4584: rom = 1'b1;
		4585: rom = 1'b1;
		4586: rom = 1'b1;
		4587: rom = 1'b1;
		4588: rom = 1'b1;
		4589: rom = 1'b1;
		4590: rom = 1'b1;
		4591: rom = 1'b1;
		4592: rom = 1'b1;
		4593: rom = 1'b1;
		4594: rom = 1'b0;
		4595: rom = 1'b1;
		4596: rom = 1'b1;
		4597: rom = 1'b1;
		4598: rom = 1'b1;
		4599: rom = 1'b0;
		4600: rom = 1'b0;
		4601: rom = 1'b0;
		4602: rom = 1'b0;
		4603: rom = 1'b0;
		4604: rom = 1'b0;
		4605: rom = 1'b0;
		4606: rom = 1'b0;
		4607: rom = 1'b0;
		4608: rom = 1'b0;
		4609: rom = 1'b0;
		4610: rom = 1'b0;
		4611: rom = 1'b0;
		4612: rom = 1'b0;
		4613: rom = 1'b0;
		4614: rom = 1'b0;
		4615: rom = 1'b0;
		4616: rom = 1'b0;
		4617: rom = 1'b0;
		4618: rom = 1'b0;
		4619: rom = 1'b0;
		4620: rom = 1'b0;
		4621: rom = 1'b0;
		4622: rom = 1'b0;
		4623: rom = 1'b0;
		4624: rom = 1'b0;
		4625: rom = 1'b0;
		4626: rom = 1'b0;
		4627: rom = 1'b0;
		4628: rom = 1'b0;
		4629: rom = 1'b0;
		4630: rom = 1'b0;
		4631: rom = 1'b0;
		4632: rom = 1'b0;
		4633: rom = 1'b0;
		4634: rom = 1'b0;
		4635: rom = 1'b0;
		4636: rom = 1'b0;
		4637: rom = 1'b1;
		4638: rom = 1'b1;
		4639: rom = 1'b1;
		4640: rom = 1'b1;
		4641: rom = 1'b1;
		4642: rom = 1'b1;
		4643: rom = 1'b1;
		4644: rom = 1'b1;
		4645: rom = 1'b1;
		4646: rom = 1'b1;
		4647: rom = 1'b0;
		4648: rom = 1'b0;
		4649: rom = 1'b0;
		4650: rom = 1'b0;
		4651: rom = 1'b0;
		4652: rom = 1'b0;
		4653: rom = 1'b0;
		4654: rom = 1'b0;
		4655: rom = 1'b0;
		4656: rom = 1'b0;
		4657: rom = 1'b0;
		4658: rom = 1'b1;
		4659: rom = 1'b1;
		4660: rom = 1'b1;
		4661: rom = 1'b1;
		4662: rom = 1'b1;
		4663: rom = 1'b1;
		4664: rom = 1'b1;
		4665: rom = 1'b1;
		4666: rom = 1'b1;
		4667: rom = 1'b1;
		4668: rom = 1'b1;
		4669: rom = 1'b1;
		4670: rom = 1'b1;
		4671: rom = 1'b1;
		4672: rom = 1'b1;
		4673: rom = 1'b1;
		4674: rom = 1'b1;
		4675: rom = 1'b1;
		4676: rom = 1'b1;
		4677: rom = 1'b1;
		4678: rom = 1'b1;
		4679: rom = 1'b1;
		4680: rom = 1'b0;
		4681: rom = 1'b0;
		4682: rom = 1'b1;
		4683: rom = 1'b1;
		4684: rom = 1'b1;
		4685: rom = 1'b1;
		4686: rom = 1'b1;
		4687: rom = 1'b1;
		4688: rom = 1'b1;
		4689: rom = 1'b1;
		4690: rom = 1'b1;
		4691: rom = 1'b1;
		4692: rom = 1'b1;
		4693: rom = 1'b1;
		4694: rom = 1'b1;
		4695: rom = 1'b1;
		4696: rom = 1'b1;
		4697: rom = 1'b1;
		4698: rom = 1'b1;
		4699: rom = 1'b1;
		4700: rom = 1'b1;
		4701: rom = 1'b1;
		4702: rom = 1'b1;
		4703: rom = 1'b1;
		4704: rom = 1'b1;
		4705: rom = 1'b1;
		4706: rom = 1'b1;
		4707: rom = 1'b1;
		4708: rom = 1'b1;
		4709: rom = 1'b1;
		4710: rom = 1'b1;
		4711: rom = 1'b1;
		4712: rom = 1'b1;
		4713: rom = 1'b1;
		4714: rom = 1'b1;
		4715: rom = 1'b1;
		4716: rom = 1'b1;
		4717: rom = 1'b1;
		4718: rom = 1'b1;
		4719: rom = 1'b1;
		4720: rom = 1'b1;
		4721: rom = 1'b1;
		4722: rom = 1'b0;
		4723: rom = 1'b1;
		4724: rom = 1'b1;
		4725: rom = 1'b1;
		4726: rom = 1'b1;
		4727: rom = 1'b0;
		4728: rom = 1'b0;
		4729: rom = 1'b0;
		4730: rom = 1'b0;
		4731: rom = 1'b0;
		4732: rom = 1'b0;
		4733: rom = 1'b0;
		4734: rom = 1'b0;
		4735: rom = 1'b0;
		4736: rom = 1'b0;
		4737: rom = 1'b0;
		4738: rom = 1'b0;
		4739: rom = 1'b0;
		4740: rom = 1'b0;
		4741: rom = 1'b0;
		4742: rom = 1'b0;
		4743: rom = 1'b0;
		4744: rom = 1'b0;
		4745: rom = 1'b0;
		4746: rom = 1'b0;
		4747: rom = 1'b0;
		4748: rom = 1'b0;
		4749: rom = 1'b0;
		4750: rom = 1'b0;
		4751: rom = 1'b0;
		4752: rom = 1'b0;
		4753: rom = 1'b0;
		4754: rom = 1'b0;
		4755: rom = 1'b0;
		4756: rom = 1'b0;
		4757: rom = 1'b0;
		4758: rom = 1'b0;
		4759: rom = 1'b0;
		4760: rom = 1'b0;
		4761: rom = 1'b0;
		4762: rom = 1'b0;
		4763: rom = 1'b0;
		4764: rom = 1'b0;
		4765: rom = 1'b1;
		4766: rom = 1'b1;
		4767: rom = 1'b1;
		4768: rom = 1'b1;
		4769: rom = 1'b1;
		4770: rom = 1'b1;
		4771: rom = 1'b1;
		4772: rom = 1'b1;
		4773: rom = 1'b1;
		4774: rom = 1'b1;
		4775: rom = 1'b0;
		4776: rom = 1'b0;
		4777: rom = 1'b0;
		4778: rom = 1'b0;
		4779: rom = 1'b0;
		4780: rom = 1'b0;
		4781: rom = 1'b0;
		4782: rom = 1'b0;
		4783: rom = 1'b0;
		4784: rom = 1'b0;
		4785: rom = 1'b1;
		4786: rom = 1'b1;
		4787: rom = 1'b1;
		4788: rom = 1'b1;
		4789: rom = 1'b1;
		4790: rom = 1'b1;
		4791: rom = 1'b1;
		4792: rom = 1'b1;
		4793: rom = 1'b1;
		4794: rom = 1'b1;
		4795: rom = 1'b1;
		4796: rom = 1'b1;
		4797: rom = 1'b1;
		4798: rom = 1'b1;
		4799: rom = 1'b1;
		4800: rom = 1'b1;
		4801: rom = 1'b1;
		4802: rom = 1'b1;
		4803: rom = 1'b1;
		4804: rom = 1'b1;
		4805: rom = 1'b1;
		4806: rom = 1'b1;
		4807: rom = 1'b1;
		4808: rom = 1'b1;
		4809: rom = 1'b0;
		4810: rom = 1'b1;
		4811: rom = 1'b1;
		4812: rom = 1'b1;
		4813: rom = 1'b1;
		4814: rom = 1'b1;
		4815: rom = 1'b1;
		4816: rom = 1'b1;
		4817: rom = 1'b1;
		4818: rom = 1'b1;
		4819: rom = 1'b1;
		4820: rom = 1'b1;
		4821: rom = 1'b1;
		4822: rom = 1'b1;
		4823: rom = 1'b1;
		4824: rom = 1'b1;
		4825: rom = 1'b1;
		4826: rom = 1'b1;
		4827: rom = 1'b1;
		4828: rom = 1'b1;
		4829: rom = 1'b1;
		4830: rom = 1'b1;
		4831: rom = 1'b1;
		4832: rom = 1'b1;
		4833: rom = 1'b1;
		4834: rom = 1'b1;
		4835: rom = 1'b1;
		4836: rom = 1'b1;
		4837: rom = 1'b1;
		4838: rom = 1'b1;
		4839: rom = 1'b1;
		4840: rom = 1'b1;
		4841: rom = 1'b1;
		4842: rom = 1'b1;
		4843: rom = 1'b1;
		4844: rom = 1'b1;
		4845: rom = 1'b1;
		4846: rom = 1'b1;
		4847: rom = 1'b1;
		4848: rom = 1'b1;
		4849: rom = 1'b0;
		4850: rom = 1'b1;
		4851: rom = 1'b1;
		4852: rom = 1'b1;
		4853: rom = 1'b1;
		4854: rom = 1'b1;
		4855: rom = 1'b0;
		4856: rom = 1'b0;
		4857: rom = 1'b0;
		4858: rom = 1'b0;
		4859: rom = 1'b0;
		4860: rom = 1'b0;
		4861: rom = 1'b0;
		4862: rom = 1'b0;
		4863: rom = 1'b0;
		4864: rom = 1'b0;
		4865: rom = 1'b0;
		4866: rom = 1'b0;
		4867: rom = 1'b0;
		4868: rom = 1'b0;
		4869: rom = 1'b0;
		4870: rom = 1'b0;
		4871: rom = 1'b0;
		4872: rom = 1'b0;
		4873: rom = 1'b0;
		4874: rom = 1'b0;
		4875: rom = 1'b0;
		4876: rom = 1'b0;
		4877: rom = 1'b0;
		4878: rom = 1'b0;
		4879: rom = 1'b0;
		4880: rom = 1'b0;
		4881: rom = 1'b0;
		4882: rom = 1'b0;
		4883: rom = 1'b0;
		4884: rom = 1'b0;
		4885: rom = 1'b0;
		4886: rom = 1'b0;
		4887: rom = 1'b0;
		4888: rom = 1'b0;
		4889: rom = 1'b0;
		4890: rom = 1'b0;
		4891: rom = 1'b0;
		4892: rom = 1'b0;
		4893: rom = 1'b1;
		4894: rom = 1'b1;
		4895: rom = 1'b1;
		4896: rom = 1'b1;
		4897: rom = 1'b1;
		4898: rom = 1'b1;
		4899: rom = 1'b1;
		4900: rom = 1'b1;
		4901: rom = 1'b1;
		4902: rom = 1'b0;
		4903: rom = 1'b0;
		4904: rom = 1'b0;
		4905: rom = 1'b0;
		4906: rom = 1'b0;
		4907: rom = 1'b0;
		4908: rom = 1'b0;
		4909: rom = 1'b0;
		4910: rom = 1'b0;
		4911: rom = 1'b0;
		4912: rom = 1'b0;
		4913: rom = 1'b1;
		4914: rom = 1'b1;
		4915: rom = 1'b1;
		4916: rom = 1'b1;
		4917: rom = 1'b1;
		4918: rom = 1'b1;
		4919: rom = 1'b1;
		4920: rom = 1'b1;
		4921: rom = 1'b1;
		4922: rom = 1'b1;
		4923: rom = 1'b1;
		4924: rom = 1'b0;
		4925: rom = 1'b1;
		4926: rom = 1'b1;
		4927: rom = 1'b1;
		4928: rom = 1'b1;
		4929: rom = 1'b1;
		4930: rom = 1'b1;
		4931: rom = 1'b1;
		4932: rom = 1'b1;
		4933: rom = 1'b1;
		4934: rom = 1'b1;
		4935: rom = 1'b1;
		4936: rom = 1'b1;
		4937: rom = 1'b1;
		4938: rom = 1'b1;
		4939: rom = 1'b1;
		4940: rom = 1'b1;
		4941: rom = 1'b1;
		4942: rom = 1'b1;
		4943: rom = 1'b1;
		4944: rom = 1'b1;
		4945: rom = 1'b1;
		4946: rom = 1'b1;
		4947: rom = 1'b1;
		4948: rom = 1'b1;
		4949: rom = 1'b1;
		4950: rom = 1'b1;
		4951: rom = 1'b1;
		4952: rom = 1'b1;
		4953: rom = 1'b1;
		4954: rom = 1'b1;
		4955: rom = 1'b1;
		4956: rom = 1'b1;
		4957: rom = 1'b1;
		4958: rom = 1'b1;
		4959: rom = 1'b1;
		4960: rom = 1'b1;
		4961: rom = 1'b1;
		4962: rom = 1'b1;
		4963: rom = 1'b1;
		4964: rom = 1'b1;
		4965: rom = 1'b1;
		4966: rom = 1'b1;
		4967: rom = 1'b1;
		4968: rom = 1'b1;
		4969: rom = 1'b1;
		4970: rom = 1'b1;
		4971: rom = 1'b1;
		4972: rom = 1'b1;
		4973: rom = 1'b1;
		4974: rom = 1'b1;
		4975: rom = 1'b1;
		4976: rom = 1'b0;
		4977: rom = 1'b0;
		4978: rom = 1'b1;
		4979: rom = 1'b1;
		4980: rom = 1'b1;
		4981: rom = 1'b1;
		4982: rom = 1'b1;
		4983: rom = 1'b0;
		4984: rom = 1'b0;
		4985: rom = 1'b0;
		4986: rom = 1'b0;
		4987: rom = 1'b0;
		4988: rom = 1'b0;
		4989: rom = 1'b0;
		4990: rom = 1'b0;
		4991: rom = 1'b0;
		4992: rom = 1'b0;
		4993: rom = 1'b0;
		4994: rom = 1'b0;
		4995: rom = 1'b0;
		4996: rom = 1'b0;
		4997: rom = 1'b0;
		4998: rom = 1'b0;
		4999: rom = 1'b0;
		5000: rom = 1'b0;
		5001: rom = 1'b0;
		5002: rom = 1'b0;
		5003: rom = 1'b0;
		5004: rom = 1'b0;
		5005: rom = 1'b0;
		5006: rom = 1'b0;
		5007: rom = 1'b0;
		5008: rom = 1'b0;
		5009: rom = 1'b0;
		5010: rom = 1'b0;
		5011: rom = 1'b0;
		5012: rom = 1'b0;
		5013: rom = 1'b0;
		5014: rom = 1'b0;
		5015: rom = 1'b0;
		5016: rom = 1'b0;
		5017: rom = 1'b0;
		5018: rom = 1'b0;
		5019: rom = 1'b0;
		5020: rom = 1'b1;
		5021: rom = 1'b1;
		5022: rom = 1'b1;
		5023: rom = 1'b1;
		5024: rom = 1'b1;
		5025: rom = 1'b1;
		5026: rom = 1'b1;
		5027: rom = 1'b1;
		5028: rom = 1'b1;
		5029: rom = 1'b0;
		5030: rom = 1'b0;
		5031: rom = 1'b0;
		5032: rom = 1'b0;
		5033: rom = 1'b0;
		5034: rom = 1'b0;
		5035: rom = 1'b0;
		5036: rom = 1'b0;
		5037: rom = 1'b0;
		5038: rom = 1'b0;
		5039: rom = 1'b0;
		5040: rom = 1'b1;
		5041: rom = 1'b1;
		5042: rom = 1'b1;
		5043: rom = 1'b1;
		5044: rom = 1'b1;
		5045: rom = 1'b1;
		5046: rom = 1'b1;
		5047: rom = 1'b1;
		5048: rom = 1'b1;
		5049: rom = 1'b1;
		5050: rom = 1'b1;
		5051: rom = 1'b0;
		5052: rom = 1'b0;
		5053: rom = 1'b0;
		5054: rom = 1'b1;
		5055: rom = 1'b1;
		5056: rom = 1'b1;
		5057: rom = 1'b1;
		5058: rom = 1'b1;
		5059: rom = 1'b1;
		5060: rom = 1'b1;
		5061: rom = 1'b1;
		5062: rom = 1'b1;
		5063: rom = 1'b1;
		5064: rom = 1'b1;
		5065: rom = 1'b1;
		5066: rom = 1'b1;
		5067: rom = 1'b1;
		5068: rom = 1'b1;
		5069: rom = 1'b1;
		5070: rom = 1'b1;
		5071: rom = 1'b1;
		5072: rom = 1'b1;
		5073: rom = 1'b1;
		5074: rom = 1'b1;
		5075: rom = 1'b1;
		5076: rom = 1'b1;
		5077: rom = 1'b1;
		5078: rom = 1'b1;
		5079: rom = 1'b1;
		5080: rom = 1'b1;
		5081: rom = 1'b1;
		5082: rom = 1'b1;
		5083: rom = 1'b1;
		5084: rom = 1'b1;
		5085: rom = 1'b1;
		5086: rom = 1'b1;
		5087: rom = 1'b1;
		5088: rom = 1'b1;
		5089: rom = 1'b1;
		5090: rom = 1'b1;
		5091: rom = 1'b1;
		5092: rom = 1'b1;
		5093: rom = 1'b1;
		5094: rom = 1'b1;
		5095: rom = 1'b1;
		5096: rom = 1'b1;
		5097: rom = 1'b1;
		5098: rom = 1'b1;
		5099: rom = 1'b1;
		5100: rom = 1'b1;
		5101: rom = 1'b1;
		5102: rom = 1'b1;
		5103: rom = 1'b1;
		5104: rom = 1'b0;
		5105: rom = 1'b1;
		5106: rom = 1'b1;
		5107: rom = 1'b1;
		5108: rom = 1'b1;
		5109: rom = 1'b1;
		5110: rom = 1'b1;
		5111: rom = 1'b0;
		5112: rom = 1'b0;
		5113: rom = 1'b0;
		5114: rom = 1'b0;
		5115: rom = 1'b0;
		5116: rom = 1'b0;
		5117: rom = 1'b0;
		5118: rom = 1'b0;
		5119: rom = 1'b0;
		5120: rom = 1'b0;
		5121: rom = 1'b0;
		5122: rom = 1'b0;
		5123: rom = 1'b0;
		5124: rom = 1'b0;
		5125: rom = 1'b0;
		5126: rom = 1'b0;
		5127: rom = 1'b0;
		5128: rom = 1'b0;
		5129: rom = 1'b0;
		5130: rom = 1'b0;
		5131: rom = 1'b0;
		5132: rom = 1'b0;
		5133: rom = 1'b0;
		5134: rom = 1'b0;
		5135: rom = 1'b0;
		5136: rom = 1'b0;
		5137: rom = 1'b0;
		5138: rom = 1'b0;
		5139: rom = 1'b0;
		5140: rom = 1'b0;
		5141: rom = 1'b0;
		5142: rom = 1'b0;
		5143: rom = 1'b0;
		5144: rom = 1'b0;
		5145: rom = 1'b0;
		5146: rom = 1'b0;
		5147: rom = 1'b0;
		5148: rom = 1'b1;
		5149: rom = 1'b1;
		5150: rom = 1'b1;
		5151: rom = 1'b1;
		5152: rom = 1'b1;
		5153: rom = 1'b1;
		5154: rom = 1'b1;
		5155: rom = 1'b1;
		5156: rom = 1'b1;
		5157: rom = 1'b0;
		5158: rom = 1'b0;
		5159: rom = 1'b0;
		5160: rom = 1'b0;
		5161: rom = 1'b0;
		5162: rom = 1'b0;
		5163: rom = 1'b0;
		5164: rom = 1'b0;
		5165: rom = 1'b0;
		5166: rom = 1'b0;
		5167: rom = 1'b1;
		5168: rom = 1'b1;
		5169: rom = 1'b1;
		5170: rom = 1'b1;
		5171: rom = 1'b1;
		5172: rom = 1'b1;
		5173: rom = 1'b1;
		5174: rom = 1'b1;
		5175: rom = 1'b1;
		5176: rom = 1'b1;
		5177: rom = 1'b1;
		5178: rom = 1'b1;
		5179: rom = 1'b0;
		5180: rom = 1'b0;
		5181: rom = 1'b0;
		5182: rom = 1'b1;
		5183: rom = 1'b1;
		5184: rom = 1'b1;
		5185: rom = 1'b1;
		5186: rom = 1'b1;
		5187: rom = 1'b1;
		5188: rom = 1'b1;
		5189: rom = 1'b1;
		5190: rom = 1'b1;
		5191: rom = 1'b1;
		5192: rom = 1'b1;
		5193: rom = 1'b1;
		5194: rom = 1'b1;
		5195: rom = 1'b1;
		5196: rom = 1'b1;
		5197: rom = 1'b1;
		5198: rom = 1'b1;
		5199: rom = 1'b1;
		5200: rom = 1'b1;
		5201: rom = 1'b1;
		5202: rom = 1'b1;
		5203: rom = 1'b1;
		5204: rom = 1'b1;
		5205: rom = 1'b1;
		5206: rom = 1'b1;
		5207: rom = 1'b1;
		5208: rom = 1'b1;
		5209: rom = 1'b1;
		5210: rom = 1'b1;
		5211: rom = 1'b1;
		5212: rom = 1'b1;
		5213: rom = 1'b1;
		5214: rom = 1'b1;
		5215: rom = 1'b1;
		5216: rom = 1'b1;
		5217: rom = 1'b1;
		5218: rom = 1'b1;
		5219: rom = 1'b1;
		5220: rom = 1'b1;
		5221: rom = 1'b1;
		5222: rom = 1'b1;
		5223: rom = 1'b1;
		5224: rom = 1'b1;
		5225: rom = 1'b1;
		5226: rom = 1'b1;
		5227: rom = 1'b1;
		5228: rom = 1'b1;
		5229: rom = 1'b1;
		5230: rom = 1'b1;
		5231: rom = 1'b0;
		5232: rom = 1'b0;
		5233: rom = 1'b1;
		5234: rom = 1'b1;
		5235: rom = 1'b1;
		5236: rom = 1'b1;
		5237: rom = 1'b1;
		5238: rom = 1'b1;
		5239: rom = 1'b0;
		5240: rom = 1'b0;
		5241: rom = 1'b0;
		5242: rom = 1'b0;
		5243: rom = 1'b0;
		5244: rom = 1'b0;
		5245: rom = 1'b0;
		5246: rom = 1'b0;
		5247: rom = 1'b0;
		5248: rom = 1'b0;
		5249: rom = 1'b0;
		5250: rom = 1'b0;
		5251: rom = 1'b0;
		5252: rom = 1'b0;
		5253: rom = 1'b0;
		5254: rom = 1'b0;
		5255: rom = 1'b0;
		5256: rom = 1'b0;
		5257: rom = 1'b0;
		5258: rom = 1'b0;
		5259: rom = 1'b0;
		5260: rom = 1'b0;
		5261: rom = 1'b0;
		5262: rom = 1'b0;
		5263: rom = 1'b0;
		5264: rom = 1'b0;
		5265: rom = 1'b0;
		5266: rom = 1'b0;
		5267: rom = 1'b0;
		5268: rom = 1'b0;
		5269: rom = 1'b0;
		5270: rom = 1'b0;
		5271: rom = 1'b0;
		5272: rom = 1'b0;
		5273: rom = 1'b0;
		5274: rom = 1'b0;
		5275: rom = 1'b0;
		5276: rom = 1'b1;
		5277: rom = 1'b1;
		5278: rom = 1'b1;
		5279: rom = 1'b1;
		5280: rom = 1'b1;
		5281: rom = 1'b1;
		5282: rom = 1'b1;
		5283: rom = 1'b1;
		5284: rom = 1'b0;
		5285: rom = 1'b0;
		5286: rom = 1'b0;
		5287: rom = 1'b0;
		5288: rom = 1'b0;
		5289: rom = 1'b0;
		5290: rom = 1'b0;
		5291: rom = 1'b0;
		5292: rom = 1'b0;
		5293: rom = 1'b0;
		5294: rom = 1'b1;
		5295: rom = 1'b1;
		5296: rom = 1'b1;
		5297: rom = 1'b1;
		5298: rom = 1'b1;
		5299: rom = 1'b1;
		5300: rom = 1'b1;
		5301: rom = 1'b1;
		5302: rom = 1'b1;
		5303: rom = 1'b1;
		5304: rom = 1'b1;
		5305: rom = 1'b1;
		5306: rom = 1'b0;
		5307: rom = 1'b0;
		5308: rom = 1'b0;
		5309: rom = 1'b0;
		5310: rom = 1'b1;
		5311: rom = 1'b1;
		5312: rom = 1'b1;
		5313: rom = 1'b1;
		5314: rom = 1'b1;
		5315: rom = 1'b1;
		5316: rom = 1'b1;
		5317: rom = 1'b1;
		5318: rom = 1'b1;
		5319: rom = 1'b1;
		5320: rom = 1'b1;
		5321: rom = 1'b1;
		5322: rom = 1'b1;
		5323: rom = 1'b1;
		5324: rom = 1'b1;
		5325: rom = 1'b1;
		5326: rom = 1'b1;
		5327: rom = 1'b1;
		5328: rom = 1'b1;
		5329: rom = 1'b1;
		5330: rom = 1'b1;
		5331: rom = 1'b1;
		5332: rom = 1'b1;
		5333: rom = 1'b1;
		5334: rom = 1'b1;
		5335: rom = 1'b1;
		5336: rom = 1'b1;
		5337: rom = 1'b1;
		5338: rom = 1'b1;
		5339: rom = 1'b1;
		5340: rom = 1'b1;
		5341: rom = 1'b1;
		5342: rom = 1'b1;
		5343: rom = 1'b1;
		5344: rom = 1'b1;
		5345: rom = 1'b1;
		5346: rom = 1'b1;
		5347: rom = 1'b1;
		5348: rom = 1'b1;
		5349: rom = 1'b1;
		5350: rom = 1'b1;
		5351: rom = 1'b1;
		5352: rom = 1'b1;
		5353: rom = 1'b1;
		5354: rom = 1'b1;
		5355: rom = 1'b1;
		5356: rom = 1'b1;
		5357: rom = 1'b1;
		5358: rom = 1'b1;
		5359: rom = 1'b0;
		5360: rom = 1'b1;
		5361: rom = 1'b1;
		5362: rom = 1'b1;
		5363: rom = 1'b1;
		5364: rom = 1'b1;
		5365: rom = 1'b1;
		5366: rom = 1'b1;
		5367: rom = 1'b0;
		5368: rom = 1'b0;
		5369: rom = 1'b0;
		5370: rom = 1'b0;
		5371: rom = 1'b0;
		5372: rom = 1'b0;
		5373: rom = 1'b0;
		5374: rom = 1'b0;
		5375: rom = 1'b0;
		5376: rom = 1'b0;
		5377: rom = 1'b0;
		5378: rom = 1'b0;
		5379: rom = 1'b0;
		5380: rom = 1'b0;
		5381: rom = 1'b0;
		5382: rom = 1'b0;
		5383: rom = 1'b0;
		5384: rom = 1'b0;
		5385: rom = 1'b0;
		5386: rom = 1'b0;
		5387: rom = 1'b0;
		5388: rom = 1'b0;
		5389: rom = 1'b0;
		5390: rom = 1'b0;
		5391: rom = 1'b0;
		5392: rom = 1'b0;
		5393: rom = 1'b0;
		5394: rom = 1'b0;
		5395: rom = 1'b0;
		5396: rom = 1'b0;
		5397: rom = 1'b0;
		5398: rom = 1'b0;
		5399: rom = 1'b0;
		5400: rom = 1'b0;
		5401: rom = 1'b0;
		5402: rom = 1'b0;
		5403: rom = 1'b0;
		5404: rom = 1'b1;
		5405: rom = 1'b1;
		5406: rom = 1'b1;
		5407: rom = 1'b1;
		5408: rom = 1'b1;
		5409: rom = 1'b1;
		5410: rom = 1'b1;
		5411: rom = 1'b1;
		5412: rom = 1'b0;
		5413: rom = 1'b0;
		5414: rom = 1'b0;
		5415: rom = 1'b0;
		5416: rom = 1'b0;
		5417: rom = 1'b0;
		5418: rom = 1'b0;
		5419: rom = 1'b0;
		5420: rom = 1'b0;
		5421: rom = 1'b0;
		5422: rom = 1'b1;
		5423: rom = 1'b1;
		5424: rom = 1'b1;
		5425: rom = 1'b1;
		5426: rom = 1'b1;
		5427: rom = 1'b1;
		5428: rom = 1'b1;
		5429: rom = 1'b1;
		5430: rom = 1'b1;
		5431: rom = 1'b1;
		5432: rom = 1'b1;
		5433: rom = 1'b1;
		5434: rom = 1'b0;
		5435: rom = 1'b0;
		5436: rom = 1'b0;
		5437: rom = 1'b0;
		5438: rom = 1'b0;
		5439: rom = 1'b1;
		5440: rom = 1'b1;
		5441: rom = 1'b1;
		5442: rom = 1'b1;
		5443: rom = 1'b1;
		5444: rom = 1'b1;
		5445: rom = 1'b1;
		5446: rom = 1'b1;
		5447: rom = 1'b1;
		5448: rom = 1'b1;
		5449: rom = 1'b1;
		5450: rom = 1'b1;
		5451: rom = 1'b1;
		5452: rom = 1'b1;
		5453: rom = 1'b1;
		5454: rom = 1'b1;
		5455: rom = 1'b1;
		5456: rom = 1'b1;
		5457: rom = 1'b1;
		5458: rom = 1'b1;
		5459: rom = 1'b1;
		5460: rom = 1'b0;
		5461: rom = 1'b1;
		5462: rom = 1'b1;
		5463: rom = 1'b1;
		5464: rom = 1'b1;
		5465: rom = 1'b1;
		5466: rom = 1'b1;
		5467: rom = 1'b1;
		5468: rom = 1'b1;
		5469: rom = 1'b1;
		5470: rom = 1'b1;
		5471: rom = 1'b1;
		5472: rom = 1'b1;
		5473: rom = 1'b1;
		5474: rom = 1'b1;
		5475: rom = 1'b1;
		5476: rom = 1'b1;
		5477: rom = 1'b1;
		5478: rom = 1'b1;
		5479: rom = 1'b1;
		5480: rom = 1'b1;
		5481: rom = 1'b1;
		5482: rom = 1'b1;
		5483: rom = 1'b1;
		5484: rom = 1'b1;
		5485: rom = 1'b1;
		5486: rom = 1'b0;
		5487: rom = 1'b0;
		5488: rom = 1'b1;
		5489: rom = 1'b1;
		5490: rom = 1'b1;
		5491: rom = 1'b1;
		5492: rom = 1'b1;
		5493: rom = 1'b1;
		5494: rom = 1'b1;
		5495: rom = 1'b0;
		5496: rom = 1'b0;
		5497: rom = 1'b0;
		5498: rom = 1'b0;
		5499: rom = 1'b0;
		5500: rom = 1'b0;
		5501: rom = 1'b0;
		5502: rom = 1'b0;
		5503: rom = 1'b0;
		5504: rom = 1'b0;
		5505: rom = 1'b0;
		5506: rom = 1'b0;
		5507: rom = 1'b0;
		5508: rom = 1'b0;
		5509: rom = 1'b0;
		5510: rom = 1'b0;
		5511: rom = 1'b0;
		5512: rom = 1'b0;
		5513: rom = 1'b0;
		5514: rom = 1'b0;
		5515: rom = 1'b0;
		5516: rom = 1'b0;
		5517: rom = 1'b0;
		5518: rom = 1'b0;
		5519: rom = 1'b0;
		5520: rom = 1'b0;
		5521: rom = 1'b0;
		5522: rom = 1'b0;
		5523: rom = 1'b0;
		5524: rom = 1'b0;
		5525: rom = 1'b0;
		5526: rom = 1'b0;
		5527: rom = 1'b0;
		5528: rom = 1'b0;
		5529: rom = 1'b0;
		5530: rom = 1'b0;
		5531: rom = 1'b0;
		5532: rom = 1'b1;
		5533: rom = 1'b1;
		5534: rom = 1'b1;
		5535: rom = 1'b1;
		5536: rom = 1'b1;
		5537: rom = 1'b1;
		5538: rom = 1'b1;
		5539: rom = 1'b0;
		5540: rom = 1'b0;
		5541: rom = 1'b0;
		5542: rom = 1'b0;
		5543: rom = 1'b0;
		5544: rom = 1'b0;
		5545: rom = 1'b0;
		5546: rom = 1'b0;
		5547: rom = 1'b0;
		5548: rom = 1'b0;
		5549: rom = 1'b1;
		5550: rom = 1'b1;
		5551: rom = 1'b1;
		5552: rom = 1'b1;
		5553: rom = 1'b1;
		5554: rom = 1'b1;
		5555: rom = 1'b1;
		5556: rom = 1'b1;
		5557: rom = 1'b1;
		5558: rom = 1'b1;
		5559: rom = 1'b1;
		5560: rom = 1'b0;
		5561: rom = 1'b0;
		5562: rom = 1'b0;
		5563: rom = 1'b0;
		5564: rom = 1'b0;
		5565: rom = 1'b0;
		5566: rom = 1'b0;
		5567: rom = 1'b1;
		5568: rom = 1'b1;
		5569: rom = 1'b1;
		5570: rom = 1'b1;
		5571: rom = 1'b1;
		5572: rom = 1'b1;
		5573: rom = 1'b1;
		5574: rom = 1'b1;
		5575: rom = 1'b1;
		5576: rom = 1'b1;
		5577: rom = 1'b1;
		5578: rom = 1'b1;
		5579: rom = 1'b1;
		5580: rom = 1'b1;
		5581: rom = 1'b1;
		5582: rom = 1'b1;
		5583: rom = 1'b1;
		5584: rom = 1'b1;
		5585: rom = 1'b1;
		5586: rom = 1'b1;
		5587: rom = 1'b1;
		5588: rom = 1'b0;
		5589: rom = 1'b1;
		5590: rom = 1'b1;
		5591: rom = 1'b1;
		5592: rom = 1'b1;
		5593: rom = 1'b1;
		5594: rom = 1'b1;
		5595: rom = 1'b1;
		5596: rom = 1'b1;
		5597: rom = 1'b1;
		5598: rom = 1'b1;
		5599: rom = 1'b1;
		5600: rom = 1'b1;
		5601: rom = 1'b1;
		5602: rom = 1'b1;
		5603: rom = 1'b1;
		5604: rom = 1'b1;
		5605: rom = 1'b1;
		5606: rom = 1'b1;
		5607: rom = 1'b1;
		5608: rom = 1'b1;
		5609: rom = 1'b1;
		5610: rom = 1'b1;
		5611: rom = 1'b1;
		5612: rom = 1'b1;
		5613: rom = 1'b1;
		5614: rom = 1'b0;
		5615: rom = 1'b1;
		5616: rom = 1'b1;
		5617: rom = 1'b1;
		5618: rom = 1'b1;
		5619: rom = 1'b1;
		5620: rom = 1'b1;
		5621: rom = 1'b1;
		5622: rom = 1'b1;
		5623: rom = 1'b0;
		5624: rom = 1'b0;
		5625: rom = 1'b0;
		5626: rom = 1'b0;
		5627: rom = 1'b0;
		5628: rom = 1'b0;
		5629: rom = 1'b0;
		5630: rom = 1'b0;
		5631: rom = 1'b0;
		5632: rom = 1'b0;
		5633: rom = 1'b0;
		5634: rom = 1'b0;
		5635: rom = 1'b0;
		5636: rom = 1'b0;
		5637: rom = 1'b0;
		5638: rom = 1'b0;
		5639: rom = 1'b0;
		5640: rom = 1'b0;
		5641: rom = 1'b0;
		5642: rom = 1'b0;
		5643: rom = 1'b0;
		5644: rom = 1'b0;
		5645: rom = 1'b0;
		5646: rom = 1'b0;
		5647: rom = 1'b0;
		5648: rom = 1'b0;
		5649: rom = 1'b0;
		5650: rom = 1'b0;
		5651: rom = 1'b0;
		5652: rom = 1'b0;
		5653: rom = 1'b0;
		5654: rom = 1'b0;
		5655: rom = 1'b0;
		5656: rom = 1'b0;
		5657: rom = 1'b0;
		5658: rom = 1'b0;
		5659: rom = 1'b0;
		5660: rom = 1'b1;
		5661: rom = 1'b1;
		5662: rom = 1'b1;
		5663: rom = 1'b1;
		5664: rom = 1'b1;
		5665: rom = 1'b1;
		5666: rom = 1'b1;
		5667: rom = 1'b0;
		5668: rom = 1'b0;
		5669: rom = 1'b0;
		5670: rom = 1'b0;
		5671: rom = 1'b0;
		5672: rom = 1'b0;
		5673: rom = 1'b0;
		5674: rom = 1'b0;
		5675: rom = 1'b0;
		5676: rom = 1'b1;
		5677: rom = 1'b1;
		5678: rom = 1'b1;
		5679: rom = 1'b1;
		5680: rom = 1'b1;
		5681: rom = 1'b1;
		5682: rom = 1'b1;
		5683: rom = 1'b1;
		5684: rom = 1'b1;
		5685: rom = 1'b1;
		5686: rom = 1'b0;
		5687: rom = 1'b0;
		5688: rom = 1'b0;
		5689: rom = 1'b0;
		5690: rom = 1'b0;
		5691: rom = 1'b0;
		5692: rom = 1'b0;
		5693: rom = 1'b0;
		5694: rom = 1'b0;
		5695: rom = 1'b0;
		5696: rom = 1'b0;
		5697: rom = 1'b1;
		5698: rom = 1'b1;
		5699: rom = 1'b1;
		5700: rom = 1'b1;
		5701: rom = 1'b1;
		5702: rom = 1'b1;
		5703: rom = 1'b1;
		5704: rom = 1'b1;
		5705: rom = 1'b1;
		5706: rom = 1'b1;
		5707: rom = 1'b1;
		5708: rom = 1'b1;
		5709: rom = 1'b1;
		5710: rom = 1'b1;
		5711: rom = 1'b1;
		5712: rom = 1'b1;
		5713: rom = 1'b1;
		5714: rom = 1'b1;
		5715: rom = 1'b0;
		5716: rom = 1'b0;
		5717: rom = 1'b0;
		5718: rom = 1'b1;
		5719: rom = 1'b1;
		5720: rom = 1'b1;
		5721: rom = 1'b1;
		5722: rom = 1'b1;
		5723: rom = 1'b1;
		5724: rom = 1'b1;
		5725: rom = 1'b1;
		5726: rom = 1'b1;
		5727: rom = 1'b1;
		5728: rom = 1'b1;
		5729: rom = 1'b1;
		5730: rom = 1'b1;
		5731: rom = 1'b1;
		5732: rom = 1'b1;
		5733: rom = 1'b1;
		5734: rom = 1'b1;
		5735: rom = 1'b1;
		5736: rom = 1'b1;
		5737: rom = 1'b1;
		5738: rom = 1'b1;
		5739: rom = 1'b1;
		5740: rom = 1'b1;
		5741: rom = 1'b0;
		5742: rom = 1'b1;
		5743: rom = 1'b1;
		5744: rom = 1'b1;
		5745: rom = 1'b1;
		5746: rom = 1'b1;
		5747: rom = 1'b1;
		5748: rom = 1'b1;
		5749: rom = 1'b1;
		5750: rom = 1'b1;
		5751: rom = 1'b0;
		5752: rom = 1'b0;
		5753: rom = 1'b0;
		5754: rom = 1'b0;
		5755: rom = 1'b0;
		5756: rom = 1'b0;
		5757: rom = 1'b0;
		5758: rom = 1'b0;
		5759: rom = 1'b0;
		5760: rom = 1'b0;
		5761: rom = 1'b0;
		5762: rom = 1'b0;
		5763: rom = 1'b0;
		5764: rom = 1'b0;
		5765: rom = 1'b0;
		5766: rom = 1'b0;
		5767: rom = 1'b0;
		5768: rom = 1'b0;
		5769: rom = 1'b0;
		5770: rom = 1'b0;
		5771: rom = 1'b0;
		5772: rom = 1'b0;
		5773: rom = 1'b0;
		5774: rom = 1'b0;
		5775: rom = 1'b0;
		5776: rom = 1'b0;
		5777: rom = 1'b0;
		5778: rom = 1'b0;
		5779: rom = 1'b0;
		5780: rom = 1'b0;
		5781: rom = 1'b0;
		5782: rom = 1'b0;
		5783: rom = 1'b0;
		5784: rom = 1'b0;
		5785: rom = 1'b0;
		5786: rom = 1'b0;
		5787: rom = 1'b1;
		5788: rom = 1'b1;
		5789: rom = 1'b1;
		5790: rom = 1'b1;
		5791: rom = 1'b1;
		5792: rom = 1'b1;
		5793: rom = 1'b1;
		5794: rom = 1'b1;
		5795: rom = 1'b0;
		5796: rom = 1'b0;
		5797: rom = 1'b0;
		5798: rom = 1'b0;
		5799: rom = 1'b0;
		5800: rom = 1'b0;
		5801: rom = 1'b0;
		5802: rom = 1'b0;
		5803: rom = 1'b0;
		5804: rom = 1'b1;
		5805: rom = 1'b1;
		5806: rom = 1'b1;
		5807: rom = 1'b1;
		5808: rom = 1'b1;
		5809: rom = 1'b1;
		5810: rom = 1'b1;
		5811: rom = 1'b1;
		5812: rom = 1'b0;
		5813: rom = 1'b0;
		5814: rom = 1'b0;
		5815: rom = 1'b0;
		5816: rom = 1'b0;
		5817: rom = 1'b0;
		5818: rom = 1'b0;
		5819: rom = 1'b0;
		5820: rom = 1'b0;
		5821: rom = 1'b0;
		5822: rom = 1'b0;
		5823: rom = 1'b0;
		5824: rom = 1'b0;
		5825: rom = 1'b0;
		5826: rom = 1'b1;
		5827: rom = 1'b1;
		5828: rom = 1'b1;
		5829: rom = 1'b1;
		5830: rom = 1'b1;
		5831: rom = 1'b1;
		5832: rom = 1'b1;
		5833: rom = 1'b1;
		5834: rom = 1'b1;
		5835: rom = 1'b1;
		5836: rom = 1'b1;
		5837: rom = 1'b1;
		5838: rom = 1'b1;
		5839: rom = 1'b1;
		5840: rom = 1'b1;
		5841: rom = 1'b0;
		5842: rom = 1'b0;
		5843: rom = 1'b0;
		5844: rom = 1'b0;
		5845: rom = 1'b0;
		5846: rom = 1'b0;
		5847: rom = 1'b0;
		5848: rom = 1'b1;
		5849: rom = 1'b1;
		5850: rom = 1'b1;
		5851: rom = 1'b1;
		5852: rom = 1'b1;
		5853: rom = 1'b1;
		5854: rom = 1'b1;
		5855: rom = 1'b1;
		5856: rom = 1'b1;
		5857: rom = 1'b1;
		5858: rom = 1'b1;
		5859: rom = 1'b1;
		5860: rom = 1'b1;
		5861: rom = 1'b1;
		5862: rom = 1'b1;
		5863: rom = 1'b1;
		5864: rom = 1'b1;
		5865: rom = 1'b1;
		5866: rom = 1'b1;
		5867: rom = 1'b1;
		5868: rom = 1'b0;
		5869: rom = 1'b0;
		5870: rom = 1'b1;
		5871: rom = 1'b1;
		5872: rom = 1'b1;
		5873: rom = 1'b1;
		5874: rom = 1'b1;
		5875: rom = 1'b1;
		5876: rom = 1'b1;
		5877: rom = 1'b1;
		5878: rom = 1'b1;
		5879: rom = 1'b0;
		5880: rom = 1'b0;
		5881: rom = 1'b0;
		5882: rom = 1'b0;
		5883: rom = 1'b0;
		5884: rom = 1'b0;
		5885: rom = 1'b0;
		5886: rom = 1'b0;
		5887: rom = 1'b0;
		5888: rom = 1'b0;
		5889: rom = 1'b0;
		5890: rom = 1'b0;
		5891: rom = 1'b0;
		5892: rom = 1'b0;
		5893: rom = 1'b0;
		5894: rom = 1'b0;
		5895: rom = 1'b0;
		5896: rom = 1'b0;
		5897: rom = 1'b0;
		5898: rom = 1'b0;
		5899: rom = 1'b0;
		5900: rom = 1'b0;
		5901: rom = 1'b0;
		5902: rom = 1'b0;
		5903: rom = 1'b0;
		5904: rom = 1'b0;
		5905: rom = 1'b0;
		5906: rom = 1'b0;
		5907: rom = 1'b0;
		5908: rom = 1'b0;
		5909: rom = 1'b0;
		5910: rom = 1'b0;
		5911: rom = 1'b0;
		5912: rom = 1'b0;
		5913: rom = 1'b0;
		5914: rom = 1'b0;
		5915: rom = 1'b1;
		5916: rom = 1'b1;
		5917: rom = 1'b1;
		5918: rom = 1'b1;
		5919: rom = 1'b1;
		5920: rom = 1'b1;
		5921: rom = 1'b1;
		5922: rom = 1'b0;
		5923: rom = 1'b0;
		5924: rom = 1'b0;
		5925: rom = 1'b0;
		5926: rom = 1'b0;
		5927: rom = 1'b0;
		5928: rom = 1'b0;
		5929: rom = 1'b0;
		5930: rom = 1'b0;
		5931: rom = 1'b1;
		5932: rom = 1'b1;
		5933: rom = 1'b1;
		5934: rom = 1'b1;
		5935: rom = 1'b1;
		5936: rom = 1'b1;
		5937: rom = 1'b1;
		5938: rom = 1'b1;
		5939: rom = 1'b1;
		5940: rom = 1'b1;
		5941: rom = 1'b0;
		5942: rom = 1'b0;
		5943: rom = 1'b0;
		5944: rom = 1'b0;
		5945: rom = 1'b0;
		5946: rom = 1'b0;
		5947: rom = 1'b0;
		5948: rom = 1'b0;
		5949: rom = 1'b0;
		5950: rom = 1'b0;
		5951: rom = 1'b0;
		5952: rom = 1'b0;
		5953: rom = 1'b0;
		5954: rom = 1'b0;
		5955: rom = 1'b0;
		5956: rom = 1'b1;
		5957: rom = 1'b1;
		5958: rom = 1'b1;
		5959: rom = 1'b1;
		5960: rom = 1'b1;
		5961: rom = 1'b1;
		5962: rom = 1'b1;
		5963: rom = 1'b1;
		5964: rom = 1'b1;
		5965: rom = 1'b1;
		5966: rom = 1'b1;
		5967: rom = 1'b1;
		5968: rom = 1'b1;
		5969: rom = 1'b1;
		5970: rom = 1'b0;
		5971: rom = 1'b0;
		5972: rom = 1'b0;
		5973: rom = 1'b0;
		5974: rom = 1'b0;
		5975: rom = 1'b1;
		5976: rom = 1'b1;
		5977: rom = 1'b1;
		5978: rom = 1'b1;
		5979: rom = 1'b1;
		5980: rom = 1'b1;
		5981: rom = 1'b1;
		5982: rom = 1'b1;
		5983: rom = 1'b1;
		5984: rom = 1'b1;
		5985: rom = 1'b1;
		5986: rom = 1'b1;
		5987: rom = 1'b1;
		5988: rom = 1'b1;
		5989: rom = 1'b1;
		5990: rom = 1'b1;
		5991: rom = 1'b1;
		5992: rom = 1'b1;
		5993: rom = 1'b1;
		5994: rom = 1'b1;
		5995: rom = 1'b0;
		5996: rom = 1'b0;
		5997: rom = 1'b1;
		5998: rom = 1'b1;
		5999: rom = 1'b1;
		6000: rom = 1'b1;
		6001: rom = 1'b1;
		6002: rom = 1'b1;
		6003: rom = 1'b1;
		6004: rom = 1'b1;
		6005: rom = 1'b1;
		6006: rom = 1'b1;
		6007: rom = 1'b0;
		6008: rom = 1'b0;
		6009: rom = 1'b0;
		6010: rom = 1'b0;
		6011: rom = 1'b0;
		6012: rom = 1'b0;
		6013: rom = 1'b0;
		6014: rom = 1'b0;
		6015: rom = 1'b0;
		6016: rom = 1'b0;
		6017: rom = 1'b0;
		6018: rom = 1'b0;
		6019: rom = 1'b0;
		6020: rom = 1'b0;
		6021: rom = 1'b0;
		6022: rom = 1'b0;
		6023: rom = 1'b0;
		6024: rom = 1'b0;
		6025: rom = 1'b0;
		6026: rom = 1'b0;
		6027: rom = 1'b0;
		6028: rom = 1'b0;
		6029: rom = 1'b0;
		6030: rom = 1'b0;
		6031: rom = 1'b0;
		6032: rom = 1'b0;
		6033: rom = 1'b0;
		6034: rom = 1'b0;
		6035: rom = 1'b0;
		6036: rom = 1'b0;
		6037: rom = 1'b0;
		6038: rom = 1'b0;
		6039: rom = 1'b0;
		6040: rom = 1'b0;
		6041: rom = 1'b0;
		6042: rom = 1'b0;
		6043: rom = 1'b1;
		6044: rom = 1'b1;
		6045: rom = 1'b1;
		6046: rom = 1'b1;
		6047: rom = 1'b1;
		6048: rom = 1'b1;
		6049: rom = 1'b1;
		6050: rom = 1'b0;
		6051: rom = 1'b0;
		6052: rom = 1'b0;
		6053: rom = 1'b0;
		6054: rom = 1'b0;
		6055: rom = 1'b0;
		6056: rom = 1'b0;
		6057: rom = 1'b0;
		6058: rom = 1'b1;
		6059: rom = 1'b1;
		6060: rom = 1'b1;
		6061: rom = 1'b1;
		6062: rom = 1'b1;
		6063: rom = 1'b1;
		6064: rom = 1'b1;
		6065: rom = 1'b1;
		6066: rom = 1'b1;
		6067: rom = 1'b1;
		6068: rom = 1'b1;
		6069: rom = 1'b1;
		6070: rom = 1'b0;
		6071: rom = 1'b0;
		6072: rom = 1'b0;
		6073: rom = 1'b0;
		6074: rom = 1'b0;
		6075: rom = 1'b0;
		6076: rom = 1'b0;
		6077: rom = 1'b0;
		6078: rom = 1'b0;
		6079: rom = 1'b0;
		6080: rom = 1'b0;
		6081: rom = 1'b0;
		6082: rom = 1'b0;
		6083: rom = 1'b1;
		6084: rom = 1'b1;
		6085: rom = 1'b1;
		6086: rom = 1'b1;
		6087: rom = 1'b1;
		6088: rom = 1'b1;
		6089: rom = 1'b1;
		6090: rom = 1'b1;
		6091: rom = 1'b1;
		6092: rom = 1'b1;
		6093: rom = 1'b1;
		6094: rom = 1'b1;
		6095: rom = 1'b1;
		6096: rom = 1'b1;
		6097: rom = 1'b1;
		6098: rom = 1'b1;
		6099: rom = 1'b1;
		6100: rom = 1'b0;
		6101: rom = 1'b1;
		6102: rom = 1'b1;
		6103: rom = 1'b1;
		6104: rom = 1'b1;
		6105: rom = 1'b1;
		6106: rom = 1'b1;
		6107: rom = 1'b1;
		6108: rom = 1'b1;
		6109: rom = 1'b1;
		6110: rom = 1'b1;
		6111: rom = 1'b1;
		6112: rom = 1'b1;
		6113: rom = 1'b1;
		6114: rom = 1'b1;
		6115: rom = 1'b1;
		6116: rom = 1'b1;
		6117: rom = 1'b1;
		6118: rom = 1'b1;
		6119: rom = 1'b1;
		6120: rom = 1'b1;
		6121: rom = 1'b1;
		6122: rom = 1'b0;
		6123: rom = 1'b1;
		6124: rom = 1'b0;
		6125: rom = 1'b1;
		6126: rom = 1'b1;
		6127: rom = 1'b1;
		6128: rom = 1'b1;
		6129: rom = 1'b1;
		6130: rom = 1'b1;
		6131: rom = 1'b1;
		6132: rom = 1'b1;
		6133: rom = 1'b1;
		6134: rom = 1'b1;
		6135: rom = 1'b0;
		6136: rom = 1'b0;
		6137: rom = 1'b0;
		6138: rom = 1'b0;
		6139: rom = 1'b0;
		6140: rom = 1'b0;
		6141: rom = 1'b0;
		6142: rom = 1'b0;
		6143: rom = 1'b0;
		6144: rom = 1'b0;
		6145: rom = 1'b0;
		6146: rom = 1'b0;
		6147: rom = 1'b0;
		6148: rom = 1'b0;
		6149: rom = 1'b0;
		6150: rom = 1'b0;
		6151: rom = 1'b0;
		6152: rom = 1'b0;
		6153: rom = 1'b0;
		6154: rom = 1'b0;
		6155: rom = 1'b0;
		6156: rom = 1'b0;
		6157: rom = 1'b0;
		6158: rom = 1'b0;
		6159: rom = 1'b0;
		6160: rom = 1'b0;
		6161: rom = 1'b0;
		6162: rom = 1'b0;
		6163: rom = 1'b0;
		6164: rom = 1'b0;
		6165: rom = 1'b0;
		6166: rom = 1'b0;
		6167: rom = 1'b0;
		6168: rom = 1'b0;
		6169: rom = 1'b0;
		6170: rom = 1'b0;
		6171: rom = 1'b1;
		6172: rom = 1'b1;
		6173: rom = 1'b1;
		6174: rom = 1'b1;
		6175: rom = 1'b1;
		6176: rom = 1'b1;
		6177: rom = 1'b0;
		6178: rom = 1'b0;
		6179: rom = 1'b0;
		6180: rom = 1'b0;
		6181: rom = 1'b0;
		6182: rom = 1'b0;
		6183: rom = 1'b0;
		6184: rom = 1'b0;
		6185: rom = 1'b0;
		6186: rom = 1'b1;
		6187: rom = 1'b1;
		6188: rom = 1'b1;
		6189: rom = 1'b1;
		6190: rom = 1'b1;
		6191: rom = 1'b1;
		6192: rom = 1'b1;
		6193: rom = 1'b1;
		6194: rom = 1'b1;
		6195: rom = 1'b1;
		6196: rom = 1'b1;
		6197: rom = 1'b1;
		6198: rom = 1'b1;
		6199: rom = 1'b1;
		6200: rom = 1'b0;
		6201: rom = 1'b0;
		6202: rom = 1'b0;
		6203: rom = 1'b0;
		6204: rom = 1'b0;
		6205: rom = 1'b0;
		6206: rom = 1'b0;
		6207: rom = 1'b0;
		6208: rom = 1'b0;
		6209: rom = 1'b1;
		6210: rom = 1'b1;
		6211: rom = 1'b1;
		6212: rom = 1'b1;
		6213: rom = 1'b1;
		6214: rom = 1'b1;
		6215: rom = 1'b1;
		6216: rom = 1'b1;
		6217: rom = 1'b1;
		6218: rom = 1'b1;
		6219: rom = 1'b1;
		6220: rom = 1'b1;
		6221: rom = 1'b1;
		6222: rom = 1'b1;
		6223: rom = 1'b1;
		6224: rom = 1'b1;
		6225: rom = 1'b1;
		6226: rom = 1'b1;
		6227: rom = 1'b1;
		6228: rom = 1'b0;
		6229: rom = 1'b1;
		6230: rom = 1'b1;
		6231: rom = 1'b1;
		6232: rom = 1'b1;
		6233: rom = 1'b1;
		6234: rom = 1'b1;
		6235: rom = 1'b1;
		6236: rom = 1'b1;
		6237: rom = 1'b1;
		6238: rom = 1'b1;
		6239: rom = 1'b1;
		6240: rom = 1'b1;
		6241: rom = 1'b1;
		6242: rom = 1'b1;
		6243: rom = 1'b1;
		6244: rom = 1'b1;
		6245: rom = 1'b1;
		6246: rom = 1'b1;
		6247: rom = 1'b1;
		6248: rom = 1'b1;
		6249: rom = 1'b0;
		6250: rom = 1'b1;
		6251: rom = 1'b0;
		6252: rom = 1'b1;
		6253: rom = 1'b1;
		6254: rom = 1'b1;
		6255: rom = 1'b1;
		6256: rom = 1'b1;
		6257: rom = 1'b1;
		6258: rom = 1'b1;
		6259: rom = 1'b1;
		6260: rom = 1'b1;
		6261: rom = 1'b1;
		6262: rom = 1'b1;
		6263: rom = 1'b0;
		6264: rom = 1'b0;
		6265: rom = 1'b0;
		6266: rom = 1'b0;
		6267: rom = 1'b0;
		6268: rom = 1'b0;
		6269: rom = 1'b0;
		6270: rom = 1'b0;
		6271: rom = 1'b0;
		6272: rom = 1'b0;
		6273: rom = 1'b0;
		6274: rom = 1'b0;
		6275: rom = 1'b0;
		6276: rom = 1'b0;
		6277: rom = 1'b0;
		6278: rom = 1'b0;
		6279: rom = 1'b0;
		6280: rom = 1'b0;
		6281: rom = 1'b0;
		6282: rom = 1'b0;
		6283: rom = 1'b0;
		6284: rom = 1'b0;
		6285: rom = 1'b0;
		6286: rom = 1'b0;
		6287: rom = 1'b0;
		6288: rom = 1'b0;
		6289: rom = 1'b0;
		6290: rom = 1'b0;
		6291: rom = 1'b0;
		6292: rom = 1'b0;
		6293: rom = 1'b0;
		6294: rom = 1'b0;
		6295: rom = 1'b0;
		6296: rom = 1'b0;
		6297: rom = 1'b0;
		6298: rom = 1'b0;
		6299: rom = 1'b1;
		6300: rom = 1'b1;
		6301: rom = 1'b1;
		6302: rom = 1'b1;
		6303: rom = 1'b1;
		6304: rom = 1'b1;
		6305: rom = 1'b0;
		6306: rom = 1'b0;
		6307: rom = 1'b0;
		6308: rom = 1'b0;
		6309: rom = 1'b0;
		6310: rom = 1'b0;
		6311: rom = 1'b0;
		6312: rom = 1'b0;
		6313: rom = 1'b1;
		6314: rom = 1'b1;
		6315: rom = 1'b1;
		6316: rom = 1'b1;
		6317: rom = 1'b1;
		6318: rom = 1'b1;
		6319: rom = 1'b1;
		6320: rom = 1'b1;
		6321: rom = 1'b1;
		6322: rom = 1'b1;
		6323: rom = 1'b1;
		6324: rom = 1'b1;
		6325: rom = 1'b1;
		6326: rom = 1'b1;
		6327: rom = 1'b1;
		6328: rom = 1'b1;
		6329: rom = 1'b0;
		6330: rom = 1'b0;
		6331: rom = 1'b0;
		6332: rom = 1'b0;
		6333: rom = 1'b0;
		6334: rom = 1'b0;
		6335: rom = 1'b1;
		6336: rom = 1'b1;
		6337: rom = 1'b1;
		6338: rom = 1'b1;
		6339: rom = 1'b1;
		6340: rom = 1'b1;
		6341: rom = 1'b1;
		6342: rom = 1'b1;
		6343: rom = 1'b1;
		6344: rom = 1'b1;
		6345: rom = 1'b1;
		6346: rom = 1'b1;
		6347: rom = 1'b1;
		6348: rom = 1'b1;
		6349: rom = 1'b1;
		6350: rom = 1'b1;
		6351: rom = 1'b1;
		6352: rom = 1'b1;
		6353: rom = 1'b1;
		6354: rom = 1'b1;
		6355: rom = 1'b1;
		6356: rom = 1'b1;
		6357: rom = 1'b1;
		6358: rom = 1'b1;
		6359: rom = 1'b1;
		6360: rom = 1'b1;
		6361: rom = 1'b1;
		6362: rom = 1'b1;
		6363: rom = 1'b1;
		6364: rom = 1'b1;
		6365: rom = 1'b1;
		6366: rom = 1'b1;
		6367: rom = 1'b1;
		6368: rom = 1'b1;
		6369: rom = 1'b1;
		6370: rom = 1'b1;
		6371: rom = 1'b1;
		6372: rom = 1'b1;
		6373: rom = 1'b1;
		6374: rom = 1'b1;
		6375: rom = 1'b1;
		6376: rom = 1'b0;
		6377: rom = 1'b1;
		6378: rom = 1'b0;
		6379: rom = 1'b0;
		6380: rom = 1'b1;
		6381: rom = 1'b1;
		6382: rom = 1'b1;
		6383: rom = 1'b1;
		6384: rom = 1'b1;
		6385: rom = 1'b1;
		6386: rom = 1'b1;
		6387: rom = 1'b1;
		6388: rom = 1'b1;
		6389: rom = 1'b1;
		6390: rom = 1'b1;
		6391: rom = 1'b0;
		6392: rom = 1'b0;
		6393: rom = 1'b0;
		6394: rom = 1'b0;
		6395: rom = 1'b0;
		6396: rom = 1'b0;
		6397: rom = 1'b0;
		6398: rom = 1'b0;
		6399: rom = 1'b0;
		6400: rom = 1'b0;
		6401: rom = 1'b0;
		6402: rom = 1'b0;
		6403: rom = 1'b0;
		6404: rom = 1'b0;
		6405: rom = 1'b0;
		6406: rom = 1'b0;
		6407: rom = 1'b0;
		6408: rom = 1'b0;
		6409: rom = 1'b0;
		6410: rom = 1'b0;
		6411: rom = 1'b0;
		6412: rom = 1'b0;
		6413: rom = 1'b0;
		6414: rom = 1'b0;
		6415: rom = 1'b0;
		6416: rom = 1'b0;
		6417: rom = 1'b0;
		6418: rom = 1'b0;
		6419: rom = 1'b0;
		6420: rom = 1'b0;
		6421: rom = 1'b0;
		6422: rom = 1'b0;
		6423: rom = 1'b0;
		6424: rom = 1'b0;
		6425: rom = 1'b0;
		6426: rom = 1'b0;
		6427: rom = 1'b1;
		6428: rom = 1'b1;
		6429: rom = 1'b1;
		6430: rom = 1'b1;
		6431: rom = 1'b1;
		6432: rom = 1'b1;
		6433: rom = 1'b0;
		6434: rom = 1'b0;
		6435: rom = 1'b0;
		6436: rom = 1'b0;
		6437: rom = 1'b0;
		6438: rom = 1'b0;
		6439: rom = 1'b0;
		6440: rom = 1'b0;
		6441: rom = 1'b1;
		6442: rom = 1'b1;
		6443: rom = 1'b1;
		6444: rom = 1'b1;
		6445: rom = 1'b1;
		6446: rom = 1'b1;
		6447: rom = 1'b1;
		6448: rom = 1'b1;
		6449: rom = 1'b1;
		6450: rom = 1'b1;
		6451: rom = 1'b1;
		6452: rom = 1'b1;
		6453: rom = 1'b1;
		6454: rom = 1'b1;
		6455: rom = 1'b1;
		6456: rom = 1'b1;
		6457: rom = 1'b1;
		6458: rom = 1'b0;
		6459: rom = 1'b0;
		6460: rom = 1'b0;
		6461: rom = 1'b0;
		6462: rom = 1'b1;
		6463: rom = 1'b1;
		6464: rom = 1'b1;
		6465: rom = 1'b1;
		6466: rom = 1'b1;
		6467: rom = 1'b1;
		6468: rom = 1'b1;
		6469: rom = 1'b1;
		6470: rom = 1'b1;
		6471: rom = 1'b1;
		6472: rom = 1'b1;
		6473: rom = 1'b1;
		6474: rom = 1'b1;
		6475: rom = 1'b1;
		6476: rom = 1'b1;
		6477: rom = 1'b1;
		6478: rom = 1'b1;
		6479: rom = 1'b1;
		6480: rom = 1'b1;
		6481: rom = 1'b1;
		6482: rom = 1'b1;
		6483: rom = 1'b1;
		6484: rom = 1'b1;
		6485: rom = 1'b1;
		6486: rom = 1'b1;
		6487: rom = 1'b1;
		6488: rom = 1'b1;
		6489: rom = 1'b1;
		6490: rom = 1'b1;
		6491: rom = 1'b1;
		6492: rom = 1'b1;
		6493: rom = 1'b1;
		6494: rom = 1'b1;
		6495: rom = 1'b1;
		6496: rom = 1'b1;
		6497: rom = 1'b1;
		6498: rom = 1'b1;
		6499: rom = 1'b1;
		6500: rom = 1'b1;
		6501: rom = 1'b1;
		6502: rom = 1'b1;
		6503: rom = 1'b0;
		6504: rom = 1'b1;
		6505: rom = 1'b1;
		6506: rom = 1'b0;
		6507: rom = 1'b1;
		6508: rom = 1'b1;
		6509: rom = 1'b1;
		6510: rom = 1'b1;
		6511: rom = 1'b1;
		6512: rom = 1'b1;
		6513: rom = 1'b1;
		6514: rom = 1'b1;
		6515: rom = 1'b1;
		6516: rom = 1'b1;
		6517: rom = 1'b1;
		6518: rom = 1'b1;
		6519: rom = 1'b0;
		6520: rom = 1'b0;
		6521: rom = 1'b0;
		6522: rom = 1'b0;
		6523: rom = 1'b0;
		6524: rom = 1'b0;
		6525: rom = 1'b0;
		6526: rom = 1'b0;
		6527: rom = 1'b0;
		6528: rom = 1'b0;
		6529: rom = 1'b0;
		6530: rom = 1'b0;
		6531: rom = 1'b0;
		6532: rom = 1'b0;
		6533: rom = 1'b0;
		6534: rom = 1'b0;
		6535: rom = 1'b0;
		6536: rom = 1'b0;
		6537: rom = 1'b0;
		6538: rom = 1'b0;
		6539: rom = 1'b0;
		6540: rom = 1'b0;
		6541: rom = 1'b0;
		6542: rom = 1'b0;
		6543: rom = 1'b0;
		6544: rom = 1'b0;
		6545: rom = 1'b0;
		6546: rom = 1'b0;
		6547: rom = 1'b0;
		6548: rom = 1'b0;
		6549: rom = 1'b0;
		6550: rom = 1'b0;
		6551: rom = 1'b0;
		6552: rom = 1'b0;
		6553: rom = 1'b0;
		6554: rom = 1'b0;
		6555: rom = 1'b1;
		6556: rom = 1'b1;
		6557: rom = 1'b1;
		6558: rom = 1'b1;
		6559: rom = 1'b1;
		6560: rom = 1'b0;
		6561: rom = 1'b0;
		6562: rom = 1'b0;
		6563: rom = 1'b0;
		6564: rom = 1'b0;
		6565: rom = 1'b0;
		6566: rom = 1'b0;
		6567: rom = 1'b0;
		6568: rom = 1'b1;
		6569: rom = 1'b1;
		6570: rom = 1'b1;
		6571: rom = 1'b1;
		6572: rom = 1'b1;
		6573: rom = 1'b1;
		6574: rom = 1'b1;
		6575: rom = 1'b1;
		6576: rom = 1'b1;
		6577: rom = 1'b1;
		6578: rom = 1'b1;
		6579: rom = 1'b1;
		6580: rom = 1'b1;
		6581: rom = 1'b1;
		6582: rom = 1'b1;
		6583: rom = 1'b1;
		6584: rom = 1'b1;
		6585: rom = 1'b1;
		6586: rom = 1'b0;
		6587: rom = 1'b0;
		6588: rom = 1'b0;
		6589: rom = 1'b0;
		6590: rom = 1'b1;
		6591: rom = 1'b1;
		6592: rom = 1'b1;
		6593: rom = 1'b1;
		6594: rom = 1'b1;
		6595: rom = 1'b1;
		6596: rom = 1'b1;
		6597: rom = 1'b1;
		6598: rom = 1'b1;
		6599: rom = 1'b1;
		6600: rom = 1'b1;
		6601: rom = 1'b1;
		6602: rom = 1'b1;
		6603: rom = 1'b1;
		6604: rom = 1'b1;
		6605: rom = 1'b1;
		6606: rom = 1'b1;
		6607: rom = 1'b1;
		6608: rom = 1'b1;
		6609: rom = 1'b1;
		6610: rom = 1'b1;
		6611: rom = 1'b1;
		6612: rom = 1'b1;
		6613: rom = 1'b1;
		6614: rom = 1'b1;
		6615: rom = 1'b1;
		6616: rom = 1'b1;
		6617: rom = 1'b1;
		6618: rom = 1'b1;
		6619: rom = 1'b1;
		6620: rom = 1'b1;
		6621: rom = 1'b1;
		6622: rom = 1'b1;
		6623: rom = 1'b1;
		6624: rom = 1'b1;
		6625: rom = 1'b1;
		6626: rom = 1'b1;
		6627: rom = 1'b1;
		6628: rom = 1'b1;
		6629: rom = 1'b1;
		6630: rom = 1'b0;
		6631: rom = 1'b1;
		6632: rom = 1'b1;
		6633: rom = 1'b0;
		6634: rom = 1'b1;
		6635: rom = 1'b1;
		6636: rom = 1'b1;
		6637: rom = 1'b1;
		6638: rom = 1'b1;
		6639: rom = 1'b1;
		6640: rom = 1'b1;
		6641: rom = 1'b1;
		6642: rom = 1'b1;
		6643: rom = 1'b1;
		6644: rom = 1'b1;
		6645: rom = 1'b1;
		6646: rom = 1'b1;
		6647: rom = 1'b0;
		6648: rom = 1'b0;
		6649: rom = 1'b0;
		6650: rom = 1'b0;
		6651: rom = 1'b0;
		6652: rom = 1'b0;
		6653: rom = 1'b0;
		6654: rom = 1'b0;
		6655: rom = 1'b0;
		6656: rom = 1'b0;
		6657: rom = 1'b0;
		6658: rom = 1'b0;
		6659: rom = 1'b0;
		6660: rom = 1'b0;
		6661: rom = 1'b0;
		6662: rom = 1'b0;
		6663: rom = 1'b0;
		6664: rom = 1'b0;
		6665: rom = 1'b0;
		6666: rom = 1'b0;
		6667: rom = 1'b0;
		6668: rom = 1'b0;
		6669: rom = 1'b0;
		6670: rom = 1'b0;
		6671: rom = 1'b0;
		6672: rom = 1'b0;
		6673: rom = 1'b0;
		6674: rom = 1'b0;
		6675: rom = 1'b0;
		6676: rom = 1'b0;
		6677: rom = 1'b0;
		6678: rom = 1'b0;
		6679: rom = 1'b0;
		6680: rom = 1'b0;
		6681: rom = 1'b0;
		6682: rom = 1'b0;
		6683: rom = 1'b1;
		6684: rom = 1'b1;
		6685: rom = 1'b1;
		6686: rom = 1'b1;
		6687: rom = 1'b1;
		6688: rom = 1'b0;
		6689: rom = 1'b0;
		6690: rom = 1'b0;
		6691: rom = 1'b0;
		6692: rom = 1'b0;
		6693: rom = 1'b0;
		6694: rom = 1'b0;
		6695: rom = 1'b0;
		6696: rom = 1'b1;
		6697: rom = 1'b1;
		6698: rom = 1'b1;
		6699: rom = 1'b1;
		6700: rom = 1'b1;
		6701: rom = 1'b1;
		6702: rom = 1'b1;
		6703: rom = 1'b1;
		6704: rom = 1'b1;
		6705: rom = 1'b1;
		6706: rom = 1'b1;
		6707: rom = 1'b1;
		6708: rom = 1'b1;
		6709: rom = 1'b1;
		6710: rom = 1'b1;
		6711: rom = 1'b1;
		6712: rom = 1'b1;
		6713: rom = 1'b1;
		6714: rom = 1'b0;
		6715: rom = 1'b0;
		6716: rom = 1'b0;
		6717: rom = 1'b1;
		6718: rom = 1'b1;
		6719: rom = 1'b1;
		6720: rom = 1'b1;
		6721: rom = 1'b1;
		6722: rom = 1'b1;
		6723: rom = 1'b1;
		6724: rom = 1'b1;
		6725: rom = 1'b1;
		6726: rom = 1'b1;
		6727: rom = 1'b1;
		6728: rom = 1'b1;
		6729: rom = 1'b1;
		6730: rom = 1'b1;
		6731: rom = 1'b1;
		6732: rom = 1'b0;
		6733: rom = 1'b0;
		6734: rom = 1'b0;
		6735: rom = 1'b0;
		6736: rom = 1'b0;
		6737: rom = 1'b0;
		6738: rom = 1'b1;
		6739: rom = 1'b1;
		6740: rom = 1'b1;
		6741: rom = 1'b1;
		6742: rom = 1'b1;
		6743: rom = 1'b1;
		6744: rom = 1'b1;
		6745: rom = 1'b1;
		6746: rom = 1'b1;
		6747: rom = 1'b1;
		6748: rom = 1'b1;
		6749: rom = 1'b1;
		6750: rom = 1'b1;
		6751: rom = 1'b1;
		6752: rom = 1'b1;
		6753: rom = 1'b1;
		6754: rom = 1'b1;
		6755: rom = 1'b1;
		6756: rom = 1'b0;
		6757: rom = 1'b0;
		6758: rom = 1'b1;
		6759: rom = 1'b1;
		6760: rom = 1'b0;
		6761: rom = 1'b0;
		6762: rom = 1'b1;
		6763: rom = 1'b1;
		6764: rom = 1'b1;
		6765: rom = 1'b1;
		6766: rom = 1'b1;
		6767: rom = 1'b1;
		6768: rom = 1'b1;
		6769: rom = 1'b1;
		6770: rom = 1'b1;
		6771: rom = 1'b1;
		6772: rom = 1'b1;
		6773: rom = 1'b1;
		6774: rom = 1'b1;
		6775: rom = 1'b0;
		6776: rom = 1'b0;
		6777: rom = 1'b0;
		6778: rom = 1'b0;
		6779: rom = 1'b0;
		6780: rom = 1'b0;
		6781: rom = 1'b0;
		6782: rom = 1'b0;
		6783: rom = 1'b0;
		6784: rom = 1'b0;
		6785: rom = 1'b0;
		6786: rom = 1'b0;
		6787: rom = 1'b0;
		6788: rom = 1'b0;
		6789: rom = 1'b0;
		6790: rom = 1'b0;
		6791: rom = 1'b0;
		6792: rom = 1'b0;
		6793: rom = 1'b0;
		6794: rom = 1'b0;
		6795: rom = 1'b0;
		6796: rom = 1'b0;
		6797: rom = 1'b0;
		6798: rom = 1'b0;
		6799: rom = 1'b0;
		6800: rom = 1'b0;
		6801: rom = 1'b0;
		6802: rom = 1'b0;
		6803: rom = 1'b0;
		6804: rom = 1'b0;
		6805: rom = 1'b0;
		6806: rom = 1'b0;
		6807: rom = 1'b0;
		6808: rom = 1'b0;
		6809: rom = 1'b0;
		6810: rom = 1'b0;
		6811: rom = 1'b1;
		6812: rom = 1'b1;
		6813: rom = 1'b1;
		6814: rom = 1'b1;
		6815: rom = 1'b1;
		6816: rom = 1'b0;
		6817: rom = 1'b0;
		6818: rom = 1'b0;
		6819: rom = 1'b0;
		6820: rom = 1'b0;
		6821: rom = 1'b0;
		6822: rom = 1'b0;
		6823: rom = 1'b1;
		6824: rom = 1'b1;
		6825: rom = 1'b1;
		6826: rom = 1'b1;
		6827: rom = 1'b1;
		6828: rom = 1'b1;
		6829: rom = 1'b1;
		6830: rom = 1'b1;
		6831: rom = 1'b1;
		6832: rom = 1'b1;
		6833: rom = 1'b1;
		6834: rom = 1'b1;
		6835: rom = 1'b1;
		6836: rom = 1'b1;
		6837: rom = 1'b1;
		6838: rom = 1'b1;
		6839: rom = 1'b1;
		6840: rom = 1'b1;
		6841: rom = 1'b1;
		6842: rom = 1'b1;
		6843: rom = 1'b0;
		6844: rom = 1'b0;
		6845: rom = 1'b1;
		6846: rom = 1'b1;
		6847: rom = 1'b1;
		6848: rom = 1'b1;
		6849: rom = 1'b1;
		6850: rom = 1'b1;
		6851: rom = 1'b1;
		6852: rom = 1'b1;
		6853: rom = 1'b1;
		6854: rom = 1'b1;
		6855: rom = 1'b1;
		6856: rom = 1'b0;
		6857: rom = 1'b0;
		6858: rom = 1'b0;
		6859: rom = 1'b0;
		6860: rom = 1'b0;
		6861: rom = 1'b0;
		6862: rom = 1'b0;
		6863: rom = 1'b0;
		6864: rom = 1'b0;
		6865: rom = 1'b0;
		6866: rom = 1'b0;
		6867: rom = 1'b0;
		6868: rom = 1'b0;
		6869: rom = 1'b0;
		6870: rom = 1'b1;
		6871: rom = 1'b1;
		6872: rom = 1'b1;
		6873: rom = 1'b1;
		6874: rom = 1'b1;
		6875: rom = 1'b1;
		6876: rom = 1'b1;
		6877: rom = 1'b1;
		6878: rom = 1'b1;
		6879: rom = 1'b1;
		6880: rom = 1'b1;
		6881: rom = 1'b1;
		6882: rom = 1'b1;
		6883: rom = 1'b1;
		6884: rom = 1'b0;
		6885: rom = 1'b1;
		6886: rom = 1'b1;
		6887: rom = 1'b1;
		6888: rom = 1'b0;
		6889: rom = 1'b1;
		6890: rom = 1'b1;
		6891: rom = 1'b1;
		6892: rom = 1'b1;
		6893: rom = 1'b1;
		6894: rom = 1'b1;
		6895: rom = 1'b1;
		6896: rom = 1'b1;
		6897: rom = 1'b1;
		6898: rom = 1'b1;
		6899: rom = 1'b1;
		6900: rom = 1'b1;
		6901: rom = 1'b1;
		6902: rom = 1'b1;
		6903: rom = 1'b0;
		6904: rom = 1'b0;
		6905: rom = 1'b0;
		6906: rom = 1'b0;
		6907: rom = 1'b0;
		6908: rom = 1'b0;
		6909: rom = 1'b0;
		6910: rom = 1'b0;
		6911: rom = 1'b0;
		6912: rom = 1'b0;
		6913: rom = 1'b0;
		6914: rom = 1'b0;
		6915: rom = 1'b0;
		6916: rom = 1'b0;
		6917: rom = 1'b0;
		6918: rom = 1'b0;
		6919: rom = 1'b0;
		6920: rom = 1'b0;
		6921: rom = 1'b0;
		6922: rom = 1'b0;
		6923: rom = 1'b0;
		6924: rom = 1'b0;
		6925: rom = 1'b0;
		6926: rom = 1'b0;
		6927: rom = 1'b0;
		6928: rom = 1'b0;
		6929: rom = 1'b0;
		6930: rom = 1'b0;
		6931: rom = 1'b0;
		6932: rom = 1'b0;
		6933: rom = 1'b0;
		6934: rom = 1'b0;
		6935: rom = 1'b0;
		6936: rom = 1'b0;
		6937: rom = 1'b0;
		6938: rom = 1'b0;
		6939: rom = 1'b0;
		6940: rom = 1'b1;
		6941: rom = 1'b1;
		6942: rom = 1'b1;
		6943: rom = 1'b0;
		6944: rom = 1'b0;
		6945: rom = 1'b0;
		6946: rom = 1'b0;
		6947: rom = 1'b0;
		6948: rom = 1'b0;
		6949: rom = 1'b0;
		6950: rom = 1'b0;
		6951: rom = 1'b1;
		6952: rom = 1'b1;
		6953: rom = 1'b1;
		6954: rom = 1'b1;
		6955: rom = 1'b1;
		6956: rom = 1'b1;
		6957: rom = 1'b1;
		6958: rom = 1'b1;
		6959: rom = 1'b1;
		6960: rom = 1'b1;
		6961: rom = 1'b1;
		6962: rom = 1'b1;
		6963: rom = 1'b1;
		6964: rom = 1'b1;
		6965: rom = 1'b1;
		6966: rom = 1'b1;
		6967: rom = 1'b1;
		6968: rom = 1'b1;
		6969: rom = 1'b1;
		6970: rom = 1'b1;
		6971: rom = 1'b0;
		6972: rom = 1'b1;
		6973: rom = 1'b1;
		6974: rom = 1'b1;
		6975: rom = 1'b1;
		6976: rom = 1'b1;
		6977: rom = 1'b1;
		6978: rom = 1'b1;
		6979: rom = 1'b1;
		6980: rom = 1'b1;
		6981: rom = 1'b0;
		6982: rom = 1'b0;
		6983: rom = 1'b0;
		6984: rom = 1'b1;
		6985: rom = 1'b1;
		6986: rom = 1'b1;
		6987: rom = 1'b1;
		6988: rom = 1'b1;
		6989: rom = 1'b1;
		6990: rom = 1'b1;
		6991: rom = 1'b1;
		6992: rom = 1'b1;
		6993: rom = 1'b1;
		6994: rom = 1'b1;
		6995: rom = 1'b1;
		6996: rom = 1'b1;
		6997: rom = 1'b0;
		6998: rom = 1'b0;
		6999: rom = 1'b0;
		7000: rom = 1'b0;
		7001: rom = 1'b1;
		7002: rom = 1'b1;
		7003: rom = 1'b1;
		7004: rom = 1'b1;
		7005: rom = 1'b1;
		7006: rom = 1'b1;
		7007: rom = 1'b1;
		7008: rom = 1'b1;
		7009: rom = 1'b1;
		7010: rom = 1'b1;
		7011: rom = 1'b0;
		7012: rom = 1'b1;
		7013: rom = 1'b1;
		7014: rom = 1'b1;
		7015: rom = 1'b0;
		7016: rom = 1'b1;
		7017: rom = 1'b1;
		7018: rom = 1'b1;
		7019: rom = 1'b1;
		7020: rom = 1'b1;
		7021: rom = 1'b1;
		7022: rom = 1'b1;
		7023: rom = 1'b1;
		7024: rom = 1'b1;
		7025: rom = 1'b1;
		7026: rom = 1'b1;
		7027: rom = 1'b1;
		7028: rom = 1'b1;
		7029: rom = 1'b1;
		7030: rom = 1'b1;
		7031: rom = 1'b0;
		7032: rom = 1'b0;
		7033: rom = 1'b0;
		7034: rom = 1'b0;
		7035: rom = 1'b0;
		7036: rom = 1'b0;
		7037: rom = 1'b0;
		7038: rom = 1'b0;
		7039: rom = 1'b0;
		7040: rom = 1'b0;
		7041: rom = 1'b0;
		7042: rom = 1'b0;
		7043: rom = 1'b0;
		7044: rom = 1'b0;
		7045: rom = 1'b0;
		7046: rom = 1'b0;
		7047: rom = 1'b0;
		7048: rom = 1'b0;
		7049: rom = 1'b0;
		7050: rom = 1'b0;
		7051: rom = 1'b0;
		7052: rom = 1'b0;
		7053: rom = 1'b0;
		7054: rom = 1'b0;
		7055: rom = 1'b0;
		7056: rom = 1'b0;
		7057: rom = 1'b0;
		7058: rom = 1'b0;
		7059: rom = 1'b0;
		7060: rom = 1'b0;
		7061: rom = 1'b0;
		7062: rom = 1'b0;
		7063: rom = 1'b0;
		7064: rom = 1'b0;
		7065: rom = 1'b0;
		7066: rom = 1'b0;
		7067: rom = 1'b0;
		7068: rom = 1'b1;
		7069: rom = 1'b1;
		7070: rom = 1'b1;
		7071: rom = 1'b0;
		7072: rom = 1'b0;
		7073: rom = 1'b0;
		7074: rom = 1'b0;
		7075: rom = 1'b0;
		7076: rom = 1'b0;
		7077: rom = 1'b0;
		7078: rom = 1'b0;
		7079: rom = 1'b1;
		7080: rom = 1'b1;
		7081: rom = 1'b1;
		7082: rom = 1'b1;
		7083: rom = 1'b1;
		7084: rom = 1'b1;
		7085: rom = 1'b1;
		7086: rom = 1'b1;
		7087: rom = 1'b1;
		7088: rom = 1'b1;
		7089: rom = 1'b1;
		7090: rom = 1'b1;
		7091: rom = 1'b1;
		7092: rom = 1'b1;
		7093: rom = 1'b1;
		7094: rom = 1'b1;
		7095: rom = 1'b1;
		7096: rom = 1'b1;
		7097: rom = 1'b1;
		7098: rom = 1'b1;
		7099: rom = 1'b1;
		7100: rom = 1'b1;
		7101: rom = 1'b1;
		7102: rom = 1'b1;
		7103: rom = 1'b1;
		7104: rom = 1'b1;
		7105: rom = 1'b1;
		7106: rom = 1'b0;
		7107: rom = 1'b0;
		7108: rom = 1'b0;
		7109: rom = 1'b1;
		7110: rom = 1'b1;
		7111: rom = 1'b1;
		7112: rom = 1'b1;
		7113: rom = 1'b1;
		7114: rom = 1'b1;
		7115: rom = 1'b1;
		7116: rom = 1'b1;
		7117: rom = 1'b1;
		7118: rom = 1'b1;
		7119: rom = 1'b1;
		7120: rom = 1'b1;
		7121: rom = 1'b1;
		7122: rom = 1'b1;
		7123: rom = 1'b1;
		7124: rom = 1'b1;
		7125: rom = 1'b1;
		7126: rom = 1'b1;
		7127: rom = 1'b1;
		7128: rom = 1'b0;
		7129: rom = 1'b0;
		7130: rom = 1'b0;
		7131: rom = 1'b0;
		7132: rom = 1'b1;
		7133: rom = 1'b1;
		7134: rom = 1'b1;
		7135: rom = 1'b1;
		7136: rom = 1'b1;
		7137: rom = 1'b0;
		7138: rom = 1'b0;
		7139: rom = 1'b1;
		7140: rom = 1'b1;
		7141: rom = 1'b1;
		7142: rom = 1'b0;
		7143: rom = 1'b1;
		7144: rom = 1'b1;
		7145: rom = 1'b1;
		7146: rom = 1'b1;
		7147: rom = 1'b1;
		7148: rom = 1'b1;
		7149: rom = 1'b1;
		7150: rom = 1'b1;
		7151: rom = 1'b1;
		7152: rom = 1'b1;
		7153: rom = 1'b1;
		7154: rom = 1'b1;
		7155: rom = 1'b1;
		7156: rom = 1'b1;
		7157: rom = 1'b1;
		7158: rom = 1'b1;
		7159: rom = 1'b0;
		7160: rom = 1'b0;
		7161: rom = 1'b0;
		7162: rom = 1'b0;
		7163: rom = 1'b0;
		7164: rom = 1'b0;
		7165: rom = 1'b0;
		7166: rom = 1'b0;
		7167: rom = 1'b0;
		7168: rom = 1'b0;
		7169: rom = 1'b0;
		7170: rom = 1'b0;
		7171: rom = 1'b0;
		7172: rom = 1'b0;
		7173: rom = 1'b0;
		7174: rom = 1'b0;
		7175: rom = 1'b0;
		7176: rom = 1'b0;
		7177: rom = 1'b0;
		7178: rom = 1'b0;
		7179: rom = 1'b0;
		7180: rom = 1'b0;
		7181: rom = 1'b0;
		7182: rom = 1'b0;
		7183: rom = 1'b0;
		7184: rom = 1'b0;
		7185: rom = 1'b0;
		7186: rom = 1'b0;
		7187: rom = 1'b0;
		7188: rom = 1'b0;
		7189: rom = 1'b0;
		7190: rom = 1'b0;
		7191: rom = 1'b0;
		7192: rom = 1'b0;
		7193: rom = 1'b0;
		7194: rom = 1'b0;
		7195: rom = 1'b0;
		7196: rom = 1'b1;
		7197: rom = 1'b1;
		7198: rom = 1'b1;
		7199: rom = 1'b0;
		7200: rom = 1'b0;
		7201: rom = 1'b0;
		7202: rom = 1'b0;
		7203: rom = 1'b0;
		7204: rom = 1'b0;
		7205: rom = 1'b0;
		7206: rom = 1'b1;
		7207: rom = 1'b1;
		7208: rom = 1'b1;
		7209: rom = 1'b1;
		7210: rom = 1'b1;
		7211: rom = 1'b1;
		7212: rom = 1'b1;
		7213: rom = 1'b1;
		7214: rom = 1'b1;
		7215: rom = 1'b1;
		7216: rom = 1'b1;
		7217: rom = 1'b1;
		7218: rom = 1'b1;
		7219: rom = 1'b1;
		7220: rom = 1'b1;
		7221: rom = 1'b1;
		7222: rom = 1'b1;
		7223: rom = 1'b1;
		7224: rom = 1'b1;
		7225: rom = 1'b1;
		7226: rom = 1'b1;
		7227: rom = 1'b1;
		7228: rom = 1'b1;
		7229: rom = 1'b1;
		7230: rom = 1'b1;
		7231: rom = 1'b1;
		7232: rom = 1'b1;
		7233: rom = 1'b0;
		7234: rom = 1'b0;
		7235: rom = 1'b1;
		7236: rom = 1'b1;
		7237: rom = 1'b1;
		7238: rom = 1'b1;
		7239: rom = 1'b1;
		7240: rom = 1'b1;
		7241: rom = 1'b1;
		7242: rom = 1'b1;
		7243: rom = 1'b1;
		7244: rom = 1'b1;
		7245: rom = 1'b1;
		7246: rom = 1'b1;
		7247: rom = 1'b1;
		7248: rom = 1'b1;
		7249: rom = 1'b1;
		7250: rom = 1'b1;
		7251: rom = 1'b1;
		7252: rom = 1'b1;
		7253: rom = 1'b1;
		7254: rom = 1'b1;
		7255: rom = 1'b1;
		7256: rom = 1'b1;
		7257: rom = 1'b1;
		7258: rom = 1'b1;
		7259: rom = 1'b0;
		7260: rom = 1'b0;
		7261: rom = 1'b0;
		7262: rom = 1'b1;
		7263: rom = 1'b1;
		7264: rom = 1'b0;
		7265: rom = 1'b0;
		7266: rom = 1'b1;
		7267: rom = 1'b1;
		7268: rom = 1'b1;
		7269: rom = 1'b1;
		7270: rom = 1'b0;
		7271: rom = 1'b1;
		7272: rom = 1'b1;
		7273: rom = 1'b1;
		7274: rom = 1'b1;
		7275: rom = 1'b1;
		7276: rom = 1'b1;
		7277: rom = 1'b1;
		7278: rom = 1'b1;
		7279: rom = 1'b1;
		7280: rom = 1'b1;
		7281: rom = 1'b1;
		7282: rom = 1'b1;
		7283: rom = 1'b1;
		7284: rom = 1'b1;
		7285: rom = 1'b1;
		7286: rom = 1'b1;
		7287: rom = 1'b0;
		7288: rom = 1'b0;
		7289: rom = 1'b0;
		7290: rom = 1'b0;
		7291: rom = 1'b0;
		7292: rom = 1'b0;
		7293: rom = 1'b0;
		7294: rom = 1'b0;
		7295: rom = 1'b0;
		7296: rom = 1'b0;
		7297: rom = 1'b0;
		7298: rom = 1'b0;
		7299: rom = 1'b0;
		7300: rom = 1'b0;
		7301: rom = 1'b0;
		7302: rom = 1'b0;
		7303: rom = 1'b0;
		7304: rom = 1'b0;
		7305: rom = 1'b0;
		7306: rom = 1'b0;
		7307: rom = 1'b0;
		7308: rom = 1'b0;
		7309: rom = 1'b0;
		7310: rom = 1'b0;
		7311: rom = 1'b0;
		7312: rom = 1'b0;
		7313: rom = 1'b0;
		7314: rom = 1'b0;
		7315: rom = 1'b0;
		7316: rom = 1'b0;
		7317: rom = 1'b0;
		7318: rom = 1'b0;
		7319: rom = 1'b0;
		7320: rom = 1'b0;
		7321: rom = 1'b0;
		7322: rom = 1'b0;
		7323: rom = 1'b0;
		7324: rom = 1'b1;
		7325: rom = 1'b1;
		7326: rom = 1'b1;
		7327: rom = 1'b0;
		7328: rom = 1'b0;
		7329: rom = 1'b0;
		7330: rom = 1'b0;
		7331: rom = 1'b0;
		7332: rom = 1'b0;
		7333: rom = 1'b1;
		7334: rom = 1'b1;
		7335: rom = 1'b1;
		7336: rom = 1'b1;
		7337: rom = 1'b1;
		7338: rom = 1'b1;
		7339: rom = 1'b1;
		7340: rom = 1'b1;
		7341: rom = 1'b1;
		7342: rom = 1'b1;
		7343: rom = 1'b1;
		7344: rom = 1'b1;
		7345: rom = 1'b1;
		7346: rom = 1'b1;
		7347: rom = 1'b1;
		7348: rom = 1'b1;
		7349: rom = 1'b1;
		7350: rom = 1'b1;
		7351: rom = 1'b1;
		7352: rom = 1'b1;
		7353: rom = 1'b1;
		7354: rom = 1'b1;
		7355: rom = 1'b1;
		7356: rom = 1'b1;
		7357: rom = 1'b1;
		7358: rom = 1'b1;
		7359: rom = 1'b0;
		7360: rom = 1'b0;
		7361: rom = 1'b1;
		7362: rom = 1'b1;
		7363: rom = 1'b1;
		7364: rom = 1'b1;
		7365: rom = 1'b1;
		7366: rom = 1'b1;
		7367: rom = 1'b1;
		7368: rom = 1'b1;
		7369: rom = 1'b1;
		7370: rom = 1'b1;
		7371: rom = 1'b1;
		7372: rom = 1'b1;
		7373: rom = 1'b1;
		7374: rom = 1'b1;
		7375: rom = 1'b1;
		7376: rom = 1'b1;
		7377: rom = 1'b1;
		7378: rom = 1'b1;
		7379: rom = 1'b1;
		7380: rom = 1'b1;
		7381: rom = 1'b1;
		7382: rom = 1'b1;
		7383: rom = 1'b1;
		7384: rom = 1'b1;
		7385: rom = 1'b1;
		7386: rom = 1'b1;
		7387: rom = 1'b1;
		7388: rom = 1'b1;
		7389: rom = 1'b0;
		7390: rom = 1'b0;
		7391: rom = 1'b0;
		7392: rom = 1'b0;
		7393: rom = 1'b1;
		7394: rom = 1'b1;
		7395: rom = 1'b1;
		7396: rom = 1'b1;
		7397: rom = 1'b0;
		7398: rom = 1'b1;
		7399: rom = 1'b1;
		7400: rom = 1'b1;
		7401: rom = 1'b1;
		7402: rom = 1'b1;
		7403: rom = 1'b1;
		7404: rom = 1'b1;
		7405: rom = 1'b1;
		7406: rom = 1'b1;
		7407: rom = 1'b1;
		7408: rom = 1'b1;
		7409: rom = 1'b1;
		7410: rom = 1'b1;
		7411: rom = 1'b1;
		7412: rom = 1'b1;
		7413: rom = 1'b1;
		7414: rom = 1'b1;
		7415: rom = 1'b0;
		7416: rom = 1'b0;
		7417: rom = 1'b0;
		7418: rom = 1'b0;
		7419: rom = 1'b0;
		7420: rom = 1'b0;
		7421: rom = 1'b0;
		7422: rom = 1'b0;
		7423: rom = 1'b0;
		7424: rom = 1'b0;
		7425: rom = 1'b0;
		7426: rom = 1'b0;
		7427: rom = 1'b0;
		7428: rom = 1'b0;
		7429: rom = 1'b0;
		7430: rom = 1'b0;
		7431: rom = 1'b0;
		7432: rom = 1'b0;
		7433: rom = 1'b0;
		7434: rom = 1'b0;
		7435: rom = 1'b0;
		7436: rom = 1'b0;
		7437: rom = 1'b0;
		7438: rom = 1'b0;
		7439: rom = 1'b0;
		7440: rom = 1'b0;
		7441: rom = 1'b0;
		7442: rom = 1'b0;
		7443: rom = 1'b0;
		7444: rom = 1'b0;
		7445: rom = 1'b0;
		7446: rom = 1'b0;
		7447: rom = 1'b0;
		7448: rom = 1'b0;
		7449: rom = 1'b0;
		7450: rom = 1'b0;
		7451: rom = 1'b0;
		7452: rom = 1'b1;
		7453: rom = 1'b1;
		7454: rom = 1'b0;
		7455: rom = 1'b0;
		7456: rom = 1'b0;
		7457: rom = 1'b0;
		7458: rom = 1'b0;
		7459: rom = 1'b0;
		7460: rom = 1'b0;
		7461: rom = 1'b1;
		7462: rom = 1'b1;
		7463: rom = 1'b1;
		7464: rom = 1'b1;
		7465: rom = 1'b1;
		7466: rom = 1'b1;
		7467: rom = 1'b1;
		7468: rom = 1'b1;
		7469: rom = 1'b1;
		7470: rom = 1'b1;
		7471: rom = 1'b1;
		7472: rom = 1'b1;
		7473: rom = 1'b1;
		7474: rom = 1'b1;
		7475: rom = 1'b1;
		7476: rom = 1'b1;
		7477: rom = 1'b1;
		7478: rom = 1'b1;
		7479: rom = 1'b1;
		7480: rom = 1'b1;
		7481: rom = 1'b1;
		7482: rom = 1'b1;
		7483: rom = 1'b1;
		7484: rom = 1'b1;
		7485: rom = 1'b1;
		7486: rom = 1'b0;
		7487: rom = 1'b0;
		7488: rom = 1'b1;
		7489: rom = 1'b1;
		7490: rom = 1'b1;
		7491: rom = 1'b1;
		7492: rom = 1'b1;
		7493: rom = 1'b1;
		7494: rom = 1'b1;
		7495: rom = 1'b1;
		7496: rom = 1'b1;
		7497: rom = 1'b1;
		7498: rom = 1'b1;
		7499: rom = 1'b1;
		7500: rom = 1'b1;
		7501: rom = 1'b1;
		7502: rom = 1'b1;
		7503: rom = 1'b1;
		7504: rom = 1'b1;
		7505: rom = 1'b1;
		7506: rom = 1'b1;
		7507: rom = 1'b1;
		7508: rom = 1'b1;
		7509: rom = 1'b1;
		7510: rom = 1'b1;
		7511: rom = 1'b1;
		7512: rom = 1'b1;
		7513: rom = 1'b1;
		7514: rom = 1'b1;
		7515: rom = 1'b1;
		7516: rom = 1'b1;
		7517: rom = 1'b1;
		7518: rom = 1'b0;
		7519: rom = 1'b0;
		7520: rom = 1'b1;
		7521: rom = 1'b1;
		7522: rom = 1'b1;
		7523: rom = 1'b1;
		7524: rom = 1'b0;
		7525: rom = 1'b0;
		7526: rom = 1'b1;
		7527: rom = 1'b1;
		7528: rom = 1'b1;
		7529: rom = 1'b1;
		7530: rom = 1'b1;
		7531: rom = 1'b1;
		7532: rom = 1'b1;
		7533: rom = 1'b1;
		7534: rom = 1'b1;
		7535: rom = 1'b1;
		7536: rom = 1'b1;
		7537: rom = 1'b1;
		7538: rom = 1'b1;
		7539: rom = 1'b1;
		7540: rom = 1'b1;
		7541: rom = 1'b1;
		7542: rom = 1'b1;
		7543: rom = 1'b0;
		7544: rom = 1'b0;
		7545: rom = 1'b0;
		7546: rom = 1'b0;
		7547: rom = 1'b0;
		7548: rom = 1'b0;
		7549: rom = 1'b0;
		7550: rom = 1'b0;
		7551: rom = 1'b0;
		7552: rom = 1'b0;
		7553: rom = 1'b0;
		7554: rom = 1'b0;
		7555: rom = 1'b0;
		7556: rom = 1'b0;
		7557: rom = 1'b0;
		7558: rom = 1'b0;
		7559: rom = 1'b0;
		7560: rom = 1'b0;
		7561: rom = 1'b0;
		7562: rom = 1'b0;
		7563: rom = 1'b0;
		7564: rom = 1'b0;
		7565: rom = 1'b0;
		7566: rom = 1'b0;
		7567: rom = 1'b0;
		7568: rom = 1'b0;
		7569: rom = 1'b0;
		7570: rom = 1'b0;
		7571: rom = 1'b0;
		7572: rom = 1'b0;
		7573: rom = 1'b0;
		7574: rom = 1'b0;
		7575: rom = 1'b0;
		7576: rom = 1'b0;
		7577: rom = 1'b0;
		7578: rom = 1'b0;
		7579: rom = 1'b0;
		7580: rom = 1'b1;
		7581: rom = 1'b1;
		7582: rom = 1'b0;
		7583: rom = 1'b0;
		7584: rom = 1'b0;
		7585: rom = 1'b0;
		7586: rom = 1'b0;
		7587: rom = 1'b0;
		7588: rom = 1'b0;
		7589: rom = 1'b1;
		7590: rom = 1'b1;
		7591: rom = 1'b1;
		7592: rom = 1'b1;
		7593: rom = 1'b1;
		7594: rom = 1'b1;
		7595: rom = 1'b1;
		7596: rom = 1'b1;
		7597: rom = 1'b1;
		7598: rom = 1'b1;
		7599: rom = 1'b1;
		7600: rom = 1'b1;
		7601: rom = 1'b1;
		7602: rom = 1'b1;
		7603: rom = 1'b1;
		7604: rom = 1'b1;
		7605: rom = 1'b1;
		7606: rom = 1'b1;
		7607: rom = 1'b1;
		7608: rom = 1'b1;
		7609: rom = 1'b1;
		7610: rom = 1'b1;
		7611: rom = 1'b1;
		7612: rom = 1'b1;
		7613: rom = 1'b0;
		7614: rom = 1'b1;
		7615: rom = 1'b1;
		7616: rom = 1'b1;
		7617: rom = 1'b1;
		7618: rom = 1'b1;
		7619: rom = 1'b1;
		7620: rom = 1'b1;
		7621: rom = 1'b1;
		7622: rom = 1'b1;
		7623: rom = 1'b1;
		7624: rom = 1'b1;
		7625: rom = 1'b1;
		7626: rom = 1'b1;
		7627: rom = 1'b1;
		7628: rom = 1'b1;
		7629: rom = 1'b1;
		7630: rom = 1'b1;
		7631: rom = 1'b1;
		7632: rom = 1'b1;
		7633: rom = 1'b1;
		7634: rom = 1'b1;
		7635: rom = 1'b1;
		7636: rom = 1'b1;
		7637: rom = 1'b1;
		7638: rom = 1'b1;
		7639: rom = 1'b1;
		7640: rom = 1'b1;
		7641: rom = 1'b1;
		7642: rom = 1'b1;
		7643: rom = 1'b1;
		7644: rom = 1'b1;
		7645: rom = 1'b1;
		7646: rom = 1'b1;
		7647: rom = 1'b1;
		7648: rom = 1'b0;
		7649: rom = 1'b0;
		7650: rom = 1'b1;
		7651: rom = 1'b1;
		7652: rom = 1'b0;
		7653: rom = 1'b1;
		7654: rom = 1'b1;
		7655: rom = 1'b1;
		7656: rom = 1'b1;
		7657: rom = 1'b1;
		7658: rom = 1'b1;
		7659: rom = 1'b1;
		7660: rom = 1'b1;
		7661: rom = 1'b1;
		7662: rom = 1'b1;
		7663: rom = 1'b1;
		7664: rom = 1'b1;
		7665: rom = 1'b1;
		7666: rom = 1'b1;
		7667: rom = 1'b1;
		7668: rom = 1'b1;
		7669: rom = 1'b1;
		7670: rom = 1'b1;
		7671: rom = 1'b0;
		7672: rom = 1'b0;
		7673: rom = 1'b0;
		7674: rom = 1'b0;
		7675: rom = 1'b0;
		7676: rom = 1'b0;
		7677: rom = 1'b0;
		7678: rom = 1'b0;
		7679: rom = 1'b0;
		7680: rom = 1'b0;
		7681: rom = 1'b0;
		7682: rom = 1'b0;
		7683: rom = 1'b0;
		7684: rom = 1'b0;
		7685: rom = 1'b0;
		7686: rom = 1'b0;
		7687: rom = 1'b0;
		7688: rom = 1'b0;
		7689: rom = 1'b0;
		7690: rom = 1'b0;
		7691: rom = 1'b0;
		7692: rom = 1'b0;
		7693: rom = 1'b0;
		7694: rom = 1'b0;
		7695: rom = 1'b0;
		7696: rom = 1'b0;
		7697: rom = 1'b0;
		7698: rom = 1'b0;
		7699: rom = 1'b0;
		7700: rom = 1'b0;
		7701: rom = 1'b0;
		7702: rom = 1'b0;
		7703: rom = 1'b0;
		7704: rom = 1'b0;
		7705: rom = 1'b0;
		7706: rom = 1'b0;
		7707: rom = 1'b0;
		7708: rom = 1'b0;
		7709: rom = 1'b1;
		7710: rom = 1'b0;
		7711: rom = 1'b0;
		7712: rom = 1'b0;
		7713: rom = 1'b0;
		7714: rom = 1'b0;
		7715: rom = 1'b0;
		7716: rom = 1'b1;
		7717: rom = 1'b1;
		7718: rom = 1'b1;
		7719: rom = 1'b1;
		7720: rom = 1'b1;
		7721: rom = 1'b1;
		7722: rom = 1'b1;
		7723: rom = 1'b1;
		7724: rom = 1'b1;
		7725: rom = 1'b1;
		7726: rom = 1'b1;
		7727: rom = 1'b1;
		7728: rom = 1'b1;
		7729: rom = 1'b1;
		7730: rom = 1'b1;
		7731: rom = 1'b1;
		7732: rom = 1'b1;
		7733: rom = 1'b1;
		7734: rom = 1'b1;
		7735: rom = 1'b1;
		7736: rom = 1'b1;
		7737: rom = 1'b1;
		7738: rom = 1'b1;
		7739: rom = 1'b1;
		7740: rom = 1'b0;
		7741: rom = 1'b1;
		7742: rom = 1'b1;
		7743: rom = 1'b1;
		7744: rom = 1'b1;
		7745: rom = 1'b1;
		7746: rom = 1'b1;
		7747: rom = 1'b1;
		7748: rom = 1'b1;
		7749: rom = 1'b1;
		7750: rom = 1'b1;
		7751: rom = 1'b1;
		7752: rom = 1'b1;
		7753: rom = 1'b1;
		7754: rom = 1'b1;
		7755: rom = 1'b1;
		7756: rom = 1'b1;
		7757: rom = 1'b1;
		7758: rom = 1'b1;
		7759: rom = 1'b1;
		7760: rom = 1'b1;
		7761: rom = 1'b1;
		7762: rom = 1'b1;
		7763: rom = 1'b1;
		7764: rom = 1'b1;
		7765: rom = 1'b1;
		7766: rom = 1'b1;
		7767: rom = 1'b1;
		7768: rom = 1'b1;
		7769: rom = 1'b1;
		7770: rom = 1'b1;
		7771: rom = 1'b1;
		7772: rom = 1'b1;
		7773: rom = 1'b1;
		7774: rom = 1'b1;
		7775: rom = 1'b1;
		7776: rom = 1'b0;
		7777: rom = 1'b0;
		7778: rom = 1'b0;
		7779: rom = 1'b0;
		7780: rom = 1'b1;
		7781: rom = 1'b1;
		7782: rom = 1'b1;
		7783: rom = 1'b1;
		7784: rom = 1'b1;
		7785: rom = 1'b1;
		7786: rom = 1'b1;
		7787: rom = 1'b1;
		7788: rom = 1'b1;
		7789: rom = 1'b1;
		7790: rom = 1'b1;
		7791: rom = 1'b1;
		7792: rom = 1'b1;
		7793: rom = 1'b1;
		7794: rom = 1'b1;
		7795: rom = 1'b1;
		7796: rom = 1'b1;
		7797: rom = 1'b1;
		7798: rom = 1'b0;
		7799: rom = 1'b0;
		7800: rom = 1'b0;
		7801: rom = 1'b0;
		7802: rom = 1'b0;
		7803: rom = 1'b0;
		7804: rom = 1'b0;
		7805: rom = 1'b0;
		7806: rom = 1'b0;
		7807: rom = 1'b0;
		7808: rom = 1'b0;
		7809: rom = 1'b0;
		7810: rom = 1'b0;
		7811: rom = 1'b0;
		7812: rom = 1'b0;
		7813: rom = 1'b0;
		7814: rom = 1'b0;
		7815: rom = 1'b0;
		7816: rom = 1'b0;
		7817: rom = 1'b0;
		7818: rom = 1'b0;
		7819: rom = 1'b0;
		7820: rom = 1'b0;
		7821: rom = 1'b0;
		7822: rom = 1'b0;
		7823: rom = 1'b0;
		7824: rom = 1'b0;
		7825: rom = 1'b0;
		7826: rom = 1'b0;
		7827: rom = 1'b0;
		7828: rom = 1'b0;
		7829: rom = 1'b0;
		7830: rom = 1'b0;
		7831: rom = 1'b0;
		7832: rom = 1'b0;
		7833: rom = 1'b0;
		7834: rom = 1'b0;
		7835: rom = 1'b0;
		7836: rom = 1'b0;
		7837: rom = 1'b0;
		7838: rom = 1'b0;
		7839: rom = 1'b0;
		7840: rom = 1'b0;
		7841: rom = 1'b0;
		7842: rom = 1'b0;
		7843: rom = 1'b0;
		7844: rom = 1'b1;
		7845: rom = 1'b1;
		7846: rom = 1'b1;
		7847: rom = 1'b1;
		7848: rom = 1'b1;
		7849: rom = 1'b1;
		7850: rom = 1'b1;
		7851: rom = 1'b1;
		7852: rom = 1'b1;
		7853: rom = 1'b1;
		7854: rom = 1'b1;
		7855: rom = 1'b1;
		7856: rom = 1'b1;
		7857: rom = 1'b1;
		7858: rom = 1'b1;
		7859: rom = 1'b1;
		7860: rom = 1'b1;
		7861: rom = 1'b1;
		7862: rom = 1'b1;
		7863: rom = 1'b1;
		7864: rom = 1'b1;
		7865: rom = 1'b1;
		7866: rom = 1'b1;
		7867: rom = 1'b0;
		7868: rom = 1'b1;
		7869: rom = 1'b1;
		7870: rom = 1'b1;
		7871: rom = 1'b1;
		7872: rom = 1'b1;
		7873: rom = 1'b1;
		7874: rom = 1'b1;
		7875: rom = 1'b1;
		7876: rom = 1'b1;
		7877: rom = 1'b1;
		7878: rom = 1'b1;
		7879: rom = 1'b1;
		7880: rom = 1'b1;
		7881: rom = 1'b1;
		7882: rom = 1'b1;
		7883: rom = 1'b1;
		7884: rom = 1'b1;
		7885: rom = 1'b1;
		7886: rom = 1'b1;
		7887: rom = 1'b1;
		7888: rom = 1'b1;
		7889: rom = 1'b1;
		7890: rom = 1'b1;
		7891: rom = 1'b1;
		7892: rom = 1'b1;
		7893: rom = 1'b1;
		7894: rom = 1'b1;
		7895: rom = 1'b1;
		7896: rom = 1'b1;
		7897: rom = 1'b1;
		7898: rom = 1'b1;
		7899: rom = 1'b1;
		7900: rom = 1'b1;
		7901: rom = 1'b1;
		7902: rom = 1'b1;
		7903: rom = 1'b1;
		7904: rom = 1'b1;
		7905: rom = 1'b1;
		7906: rom = 1'b0;
		7907: rom = 1'b0;
		7908: rom = 1'b1;
		7909: rom = 1'b1;
		7910: rom = 1'b1;
		7911: rom = 1'b1;
		7912: rom = 1'b1;
		7913: rom = 1'b1;
		7914: rom = 1'b1;
		7915: rom = 1'b1;
		7916: rom = 1'b1;
		7917: rom = 1'b1;
		7918: rom = 1'b1;
		7919: rom = 1'b1;
		7920: rom = 1'b1;
		7921: rom = 1'b1;
		7922: rom = 1'b1;
		7923: rom = 1'b1;
		7924: rom = 1'b1;
		7925: rom = 1'b1;
		7926: rom = 1'b0;
		7927: rom = 1'b0;
		7928: rom = 1'b0;
		7929: rom = 1'b0;
		7930: rom = 1'b0;
		7931: rom = 1'b0;
		7932: rom = 1'b0;
		7933: rom = 1'b0;
		7934: rom = 1'b0;
		7935: rom = 1'b0;
		7936: rom = 1'b0;
		7937: rom = 1'b0;
		7938: rom = 1'b0;
		7939: rom = 1'b0;
		7940: rom = 1'b0;
		7941: rom = 1'b0;
		7942: rom = 1'b0;
		7943: rom = 1'b0;
		7944: rom = 1'b0;
		7945: rom = 1'b0;
		7946: rom = 1'b0;
		7947: rom = 1'b0;
		7948: rom = 1'b0;
		7949: rom = 1'b0;
		7950: rom = 1'b0;
		7951: rom = 1'b0;
		7952: rom = 1'b0;
		7953: rom = 1'b0;
		7954: rom = 1'b0;
		7955: rom = 1'b0;
		7956: rom = 1'b0;
		7957: rom = 1'b0;
		7958: rom = 1'b0;
		7959: rom = 1'b0;
		7960: rom = 1'b0;
		7961: rom = 1'b0;
		7962: rom = 1'b0;
		7963: rom = 1'b0;
		7964: rom = 1'b0;
		7965: rom = 1'b0;
		7966: rom = 1'b0;
		7967: rom = 1'b0;
		7968: rom = 1'b0;
		7969: rom = 1'b0;
		7970: rom = 1'b0;
		7971: rom = 1'b0;
		7972: rom = 1'b1;
		7973: rom = 1'b1;
		7974: rom = 1'b1;
		7975: rom = 1'b1;
		7976: rom = 1'b1;
		7977: rom = 1'b1;
		7978: rom = 1'b1;
		7979: rom = 1'b1;
		7980: rom = 1'b1;
		7981: rom = 1'b1;
		7982: rom = 1'b1;
		7983: rom = 1'b1;
		7984: rom = 1'b1;
		7985: rom = 1'b1;
		7986: rom = 1'b1;
		7987: rom = 1'b1;
		7988: rom = 1'b1;
		7989: rom = 1'b1;
		7990: rom = 1'b1;
		7991: rom = 1'b1;
		7992: rom = 1'b1;
		7993: rom = 1'b1;
		7994: rom = 1'b0;
		7995: rom = 1'b1;
		7996: rom = 1'b1;
		7997: rom = 1'b1;
		7998: rom = 1'b1;
		7999: rom = 1'b1;
		8000: rom = 1'b1;
		8001: rom = 1'b1;
		8002: rom = 1'b1;
		8003: rom = 1'b1;
		8004: rom = 1'b1;
		8005: rom = 1'b1;
		8006: rom = 1'b1;
		8007: rom = 1'b1;
		8008: rom = 1'b1;
		8009: rom = 1'b1;
		8010: rom = 1'b1;
		8011: rom = 1'b1;
		8012: rom = 1'b1;
		8013: rom = 1'b1;
		8014: rom = 1'b1;
		8015: rom = 1'b1;
		8016: rom = 1'b1;
		8017: rom = 1'b1;
		8018: rom = 1'b1;
		8019: rom = 1'b1;
		8020: rom = 1'b1;
		8021: rom = 1'b1;
		8022: rom = 1'b1;
		8023: rom = 1'b1;
		8024: rom = 1'b1;
		8025: rom = 1'b1;
		8026: rom = 1'b1;
		8027: rom = 1'b1;
		8028: rom = 1'b1;
		8029: rom = 1'b1;
		8030: rom = 1'b1;
		8031: rom = 1'b1;
		8032: rom = 1'b1;
		8033: rom = 1'b1;
		8034: rom = 1'b0;
		8035: rom = 1'b1;
		8036: rom = 1'b1;
		8037: rom = 1'b1;
		8038: rom = 1'b1;
		8039: rom = 1'b1;
		8040: rom = 1'b1;
		8041: rom = 1'b1;
		8042: rom = 1'b1;
		8043: rom = 1'b1;
		8044: rom = 1'b1;
		8045: rom = 1'b1;
		8046: rom = 1'b1;
		8047: rom = 1'b1;
		8048: rom = 1'b1;
		8049: rom = 1'b1;
		8050: rom = 1'b1;
		8051: rom = 1'b1;
		8052: rom = 1'b1;
		8053: rom = 1'b1;
		8054: rom = 1'b0;
		8055: rom = 1'b0;
		8056: rom = 1'b0;
		8057: rom = 1'b0;
		8058: rom = 1'b0;
		8059: rom = 1'b0;
		8060: rom = 1'b0;
		8061: rom = 1'b0;
		8062: rom = 1'b0;
		8063: rom = 1'b0;
		8064: rom = 1'b0;
		8065: rom = 1'b0;
		8066: rom = 1'b0;
		8067: rom = 1'b0;
		8068: rom = 1'b0;
		8069: rom = 1'b0;
		8070: rom = 1'b0;
		8071: rom = 1'b0;
		8072: rom = 1'b0;
		8073: rom = 1'b0;
		8074: rom = 1'b0;
		8075: rom = 1'b0;
		8076: rom = 1'b0;
		8077: rom = 1'b0;
		8078: rom = 1'b0;
		8079: rom = 1'b0;
		8080: rom = 1'b0;
		8081: rom = 1'b0;
		8082: rom = 1'b0;
		8083: rom = 1'b0;
		8084: rom = 1'b0;
		8085: rom = 1'b0;
		8086: rom = 1'b0;
		8087: rom = 1'b0;
		8088: rom = 1'b0;
		8089: rom = 1'b0;
		8090: rom = 1'b0;
		8091: rom = 1'b0;
		8092: rom = 1'b0;
		8093: rom = 1'b0;
		8094: rom = 1'b0;
		8095: rom = 1'b0;
		8096: rom = 1'b0;
		8097: rom = 1'b0;
		8098: rom = 1'b0;
		8099: rom = 1'b1;
		8100: rom = 1'b1;
		8101: rom = 1'b1;
		8102: rom = 1'b1;
		8103: rom = 1'b1;
		8104: rom = 1'b1;
		8105: rom = 1'b1;
		8106: rom = 1'b1;
		8107: rom = 1'b1;
		8108: rom = 1'b1;
		8109: rom = 1'b1;
		8110: rom = 1'b1;
		8111: rom = 1'b1;
		8112: rom = 1'b1;
		8113: rom = 1'b1;
		8114: rom = 1'b1;
		8115: rom = 1'b1;
		8116: rom = 1'b1;
		8117: rom = 1'b1;
		8118: rom = 1'b1;
		8119: rom = 1'b1;
		8120: rom = 1'b1;
		8121: rom = 1'b0;
		8122: rom = 1'b1;
		8123: rom = 1'b1;
		8124: rom = 1'b1;
		8125: rom = 1'b1;
		8126: rom = 1'b1;
		8127: rom = 1'b1;
		8128: rom = 1'b1;
		8129: rom = 1'b1;
		8130: rom = 1'b1;
		8131: rom = 1'b1;
		8132: rom = 1'b1;
		8133: rom = 1'b1;
		8134: rom = 1'b1;
		8135: rom = 1'b1;
		8136: rom = 1'b1;
		8137: rom = 1'b1;
		8138: rom = 1'b1;
		8139: rom = 1'b1;
		8140: rom = 1'b1;
		8141: rom = 1'b1;
		8142: rom = 1'b1;
		8143: rom = 1'b1;
		8144: rom = 1'b1;
		8145: rom = 1'b1;
		8146: rom = 1'b1;
		8147: rom = 1'b1;
		8148: rom = 1'b1;
		8149: rom = 1'b1;
		8150: rom = 1'b1;
		8151: rom = 1'b1;
		8152: rom = 1'b1;
		8153: rom = 1'b1;
		8154: rom = 1'b1;
		8155: rom = 1'b1;
		8156: rom = 1'b1;
		8157: rom = 1'b1;
		8158: rom = 1'b1;
		8159: rom = 1'b1;
		8160: rom = 1'b1;
		8161: rom = 1'b0;
		8162: rom = 1'b1;
		8163: rom = 1'b1;
		8164: rom = 1'b1;
		8165: rom = 1'b1;
		8166: rom = 1'b1;
		8167: rom = 1'b1;
		8168: rom = 1'b1;
		8169: rom = 1'b1;
		8170: rom = 1'b1;
		8171: rom = 1'b1;
		8172: rom = 1'b1;
		8173: rom = 1'b1;
		8174: rom = 1'b1;
		8175: rom = 1'b1;
		8176: rom = 1'b1;
		8177: rom = 1'b1;
		8178: rom = 1'b1;
		8179: rom = 1'b1;
		8180: rom = 1'b1;
		8181: rom = 1'b1;
		8182: rom = 1'b0;
		8183: rom = 1'b0;
		8184: rom = 1'b0;
		8185: rom = 1'b0;
		8186: rom = 1'b0;
		8187: rom = 1'b0;
		8188: rom = 1'b0;
		8189: rom = 1'b0;
		8190: rom = 1'b0;
		8191: rom = 1'b0;
		8192: rom = 1'b0;
		8193: rom = 1'b0;
		8194: rom = 1'b0;
		8195: rom = 1'b0;
		8196: rom = 1'b0;
		8197: rom = 1'b0;
		8198: rom = 1'b0;
		8199: rom = 1'b0;
		8200: rom = 1'b0;
		8201: rom = 1'b0;
		8202: rom = 1'b0;
		8203: rom = 1'b0;
		8204: rom = 1'b0;
		8205: rom = 1'b0;
		8206: rom = 1'b0;
		8207: rom = 1'b0;
		8208: rom = 1'b0;
		8209: rom = 1'b0;
		8210: rom = 1'b0;
		8211: rom = 1'b0;
		8212: rom = 1'b0;
		8213: rom = 1'b0;
		8214: rom = 1'b0;
		8215: rom = 1'b0;
		8216: rom = 1'b0;
		8217: rom = 1'b0;
		8218: rom = 1'b0;
		8219: rom = 1'b0;
		8220: rom = 1'b0;
		8221: rom = 1'b0;
		8222: rom = 1'b0;
		8223: rom = 1'b0;
		8224: rom = 1'b0;
		8225: rom = 1'b0;
		8226: rom = 1'b0;
		8227: rom = 1'b1;
		8228: rom = 1'b1;
		8229: rom = 1'b1;
		8230: rom = 1'b1;
		8231: rom = 1'b1;
		8232: rom = 1'b1;
		8233: rom = 1'b1;
		8234: rom = 1'b1;
		8235: rom = 1'b1;
		8236: rom = 1'b1;
		8237: rom = 1'b1;
		8238: rom = 1'b1;
		8239: rom = 1'b1;
		8240: rom = 1'b1;
		8241: rom = 1'b1;
		8242: rom = 1'b1;
		8243: rom = 1'b1;
		8244: rom = 1'b1;
		8245: rom = 1'b1;
		8246: rom = 1'b1;
		8247: rom = 1'b1;
		8248: rom = 1'b0;
		8249: rom = 1'b1;
		8250: rom = 1'b1;
		8251: rom = 1'b1;
		8252: rom = 1'b1;
		8253: rom = 1'b1;
		8254: rom = 1'b1;
		8255: rom = 1'b1;
		8256: rom = 1'b1;
		8257: rom = 1'b1;
		8258: rom = 1'b1;
		8259: rom = 1'b1;
		8260: rom = 1'b1;
		8261: rom = 1'b1;
		8262: rom = 1'b1;
		8263: rom = 1'b1;
		8264: rom = 1'b1;
		8265: rom = 1'b1;
		8266: rom = 1'b1;
		8267: rom = 1'b1;
		8268: rom = 1'b1;
		8269: rom = 1'b1;
		8270: rom = 1'b1;
		8271: rom = 1'b1;
		8272: rom = 1'b1;
		8273: rom = 1'b1;
		8274: rom = 1'b1;
		8275: rom = 1'b1;
		8276: rom = 1'b1;
		8277: rom = 1'b1;
		8278: rom = 1'b1;
		8279: rom = 1'b1;
		8280: rom = 1'b1;
		8281: rom = 1'b1;
		8282: rom = 1'b1;
		8283: rom = 1'b1;
		8284: rom = 1'b1;
		8285: rom = 1'b1;
		8286: rom = 1'b1;
		8287: rom = 1'b1;
		8288: rom = 1'b0;
		8289: rom = 1'b1;
		8290: rom = 1'b1;
		8291: rom = 1'b1;
		8292: rom = 1'b1;
		8293: rom = 1'b1;
		8294: rom = 1'b1;
		8295: rom = 1'b1;
		8296: rom = 1'b1;
		8297: rom = 1'b1;
		8298: rom = 1'b1;
		8299: rom = 1'b1;
		8300: rom = 1'b1;
		8301: rom = 1'b1;
		8302: rom = 1'b1;
		8303: rom = 1'b1;
		8304: rom = 1'b1;
		8305: rom = 1'b1;
		8306: rom = 1'b1;
		8307: rom = 1'b1;
		8308: rom = 1'b1;
		8309: rom = 1'b1;
		8310: rom = 1'b0;
		8311: rom = 1'b0;
		8312: rom = 1'b0;
		8313: rom = 1'b0;
		8314: rom = 1'b0;
		8315: rom = 1'b0;
		8316: rom = 1'b0;
		8317: rom = 1'b0;
		8318: rom = 1'b0;
		8319: rom = 1'b0;
		8320: rom = 1'b0;
		8321: rom = 1'b0;
		8322: rom = 1'b0;
		8323: rom = 1'b0;
		8324: rom = 1'b0;
		8325: rom = 1'b0;
		8326: rom = 1'b0;
		8327: rom = 1'b0;
		8328: rom = 1'b0;
		8329: rom = 1'b0;
		8330: rom = 1'b0;
		8331: rom = 1'b0;
		8332: rom = 1'b0;
		8333: rom = 1'b0;
		8334: rom = 1'b0;
		8335: rom = 1'b0;
		8336: rom = 1'b0;
		8337: rom = 1'b0;
		8338: rom = 1'b0;
		8339: rom = 1'b0;
		8340: rom = 1'b0;
		8341: rom = 1'b0;
		8342: rom = 1'b0;
		8343: rom = 1'b0;
		8344: rom = 1'b0;
		8345: rom = 1'b0;
		8346: rom = 1'b0;
		8347: rom = 1'b0;
		8348: rom = 1'b0;
		8349: rom = 1'b0;
		8350: rom = 1'b0;
		8351: rom = 1'b0;
		8352: rom = 1'b0;
		8353: rom = 1'b0;
		8354: rom = 1'b0;
		8355: rom = 1'b1;
		8356: rom = 1'b1;
		8357: rom = 1'b1;
		8358: rom = 1'b1;
		8359: rom = 1'b1;
		8360: rom = 1'b1;
		8361: rom = 1'b1;
		8362: rom = 1'b1;
		8363: rom = 1'b1;
		8364: rom = 1'b1;
		8365: rom = 1'b1;
		8366: rom = 1'b1;
		8367: rom = 1'b1;
		8368: rom = 1'b1;
		8369: rom = 1'b1;
		8370: rom = 1'b1;
		8371: rom = 1'b1;
		8372: rom = 1'b1;
		8373: rom = 1'b1;
		8374: rom = 1'b1;
		8375: rom = 1'b1;
		8376: rom = 1'b0;
		8377: rom = 1'b1;
		8378: rom = 1'b1;
		8379: rom = 1'b1;
		8380: rom = 1'b1;
		8381: rom = 1'b1;
		8382: rom = 1'b1;
		8383: rom = 1'b1;
		8384: rom = 1'b1;
		8385: rom = 1'b1;
		8386: rom = 1'b1;
		8387: rom = 1'b1;
		8388: rom = 1'b1;
		8389: rom = 1'b1;
		8390: rom = 1'b1;
		8391: rom = 1'b1;
		8392: rom = 1'b1;
		8393: rom = 1'b1;
		8394: rom = 1'b1;
		8395: rom = 1'b1;
		8396: rom = 1'b1;
		8397: rom = 1'b1;
		8398: rom = 1'b1;
		8399: rom = 1'b1;
		8400: rom = 1'b1;
		8401: rom = 1'b1;
		8402: rom = 1'b1;
		8403: rom = 1'b1;
		8404: rom = 1'b1;
		8405: rom = 1'b1;
		8406: rom = 1'b1;
		8407: rom = 1'b1;
		8408: rom = 1'b1;
		8409: rom = 1'b1;
		8410: rom = 1'b1;
		8411: rom = 1'b1;
		8412: rom = 1'b1;
		8413: rom = 1'b1;
		8414: rom = 1'b1;
		8415: rom = 1'b0;
		8416: rom = 1'b0;
		8417: rom = 1'b1;
		8418: rom = 1'b1;
		8419: rom = 1'b1;
		8420: rom = 1'b1;
		8421: rom = 1'b1;
		8422: rom = 1'b1;
		8423: rom = 1'b1;
		8424: rom = 1'b1;
		8425: rom = 1'b1;
		8426: rom = 1'b1;
		8427: rom = 1'b1;
		8428: rom = 1'b1;
		8429: rom = 1'b1;
		8430: rom = 1'b1;
		8431: rom = 1'b1;
		8432: rom = 1'b1;
		8433: rom = 1'b1;
		8434: rom = 1'b1;
		8435: rom = 1'b1;
		8436: rom = 1'b1;
		8437: rom = 1'b1;
		8438: rom = 1'b0;
		8439: rom = 1'b0;
		8440: rom = 1'b0;
		8441: rom = 1'b0;
		8442: rom = 1'b0;
		8443: rom = 1'b0;
		8444: rom = 1'b0;
		8445: rom = 1'b0;
		8446: rom = 1'b0;
		8447: rom = 1'b0;
		8448: rom = 1'b0;
		8449: rom = 1'b0;
		8450: rom = 1'b0;
		8451: rom = 1'b0;
		8452: rom = 1'b0;
		8453: rom = 1'b0;
		8454: rom = 1'b0;
		8455: rom = 1'b0;
		8456: rom = 1'b0;
		8457: rom = 1'b0;
		8458: rom = 1'b0;
		8459: rom = 1'b0;
		8460: rom = 1'b0;
		8461: rom = 1'b0;
		8462: rom = 1'b0;
		8463: rom = 1'b0;
		8464: rom = 1'b0;
		8465: rom = 1'b0;
		8466: rom = 1'b0;
		8467: rom = 1'b0;
		8468: rom = 1'b0;
		8469: rom = 1'b0;
		8470: rom = 1'b0;
		8471: rom = 1'b0;
		8472: rom = 1'b0;
		8473: rom = 1'b0;
		8474: rom = 1'b0;
		8475: rom = 1'b0;
		8476: rom = 1'b0;
		8477: rom = 1'b0;
		8478: rom = 1'b0;
		8479: rom = 1'b0;
		8480: rom = 1'b0;
		8481: rom = 1'b0;
		8482: rom = 1'b0;
		8483: rom = 1'b1;
		8484: rom = 1'b1;
		8485: rom = 1'b1;
		8486: rom = 1'b1;
		8487: rom = 1'b1;
		8488: rom = 1'b1;
		8489: rom = 1'b1;
		8490: rom = 1'b1;
		8491: rom = 1'b1;
		8492: rom = 1'b1;
		8493: rom = 1'b1;
		8494: rom = 1'b1;
		8495: rom = 1'b1;
		8496: rom = 1'b1;
		8497: rom = 1'b1;
		8498: rom = 1'b1;
		8499: rom = 1'b1;
		8500: rom = 1'b1;
		8501: rom = 1'b1;
		8502: rom = 1'b1;
		8503: rom = 1'b0;
		8504: rom = 1'b1;
		8505: rom = 1'b1;
		8506: rom = 1'b1;
		8507: rom = 1'b1;
		8508: rom = 1'b1;
		8509: rom = 1'b1;
		8510: rom = 1'b1;
		8511: rom = 1'b1;
		8512: rom = 1'b1;
		8513: rom = 1'b1;
		8514: rom = 1'b1;
		8515: rom = 1'b1;
		8516: rom = 1'b1;
		8517: rom = 1'b1;
		8518: rom = 1'b1;
		8519: rom = 1'b1;
		8520: rom = 1'b1;
		8521: rom = 1'b1;
		8522: rom = 1'b1;
		8523: rom = 1'b1;
		8524: rom = 1'b1;
		8525: rom = 1'b1;
		8526: rom = 1'b1;
		8527: rom = 1'b1;
		8528: rom = 1'b1;
		8529: rom = 1'b1;
		8530: rom = 1'b1;
		8531: rom = 1'b1;
		8532: rom = 1'b1;
		8533: rom = 1'b1;
		8534: rom = 1'b1;
		8535: rom = 1'b1;
		8536: rom = 1'b1;
		8537: rom = 1'b1;
		8538: rom = 1'b1;
		8539: rom = 1'b1;
		8540: rom = 1'b1;
		8541: rom = 1'b1;
		8542: rom = 1'b1;
		8543: rom = 1'b0;
		8544: rom = 1'b1;
		8545: rom = 1'b1;
		8546: rom = 1'b1;
		8547: rom = 1'b1;
		8548: rom = 1'b1;
		8549: rom = 1'b1;
		8550: rom = 1'b1;
		8551: rom = 1'b1;
		8552: rom = 1'b1;
		8553: rom = 1'b1;
		8554: rom = 1'b1;
		8555: rom = 1'b1;
		8556: rom = 1'b1;
		8557: rom = 1'b1;
		8558: rom = 1'b1;
		8559: rom = 1'b1;
		8560: rom = 1'b1;
		8561: rom = 1'b1;
		8562: rom = 1'b1;
		8563: rom = 1'b1;
		8564: rom = 1'b1;
		8565: rom = 1'b1;
		8566: rom = 1'b0;
		8567: rom = 1'b0;
		8568: rom = 1'b0;
		8569: rom = 1'b0;
		8570: rom = 1'b0;
		8571: rom = 1'b0;
		8572: rom = 1'b0;
		8573: rom = 1'b0;
		8574: rom = 1'b0;
		8575: rom = 1'b0;
		8576: rom = 1'b0;
		8577: rom = 1'b0;
		8578: rom = 1'b0;
		8579: rom = 1'b0;
		8580: rom = 1'b0;
		8581: rom = 1'b0;
		8582: rom = 1'b0;
		8583: rom = 1'b0;
		8584: rom = 1'b0;
		8585: rom = 1'b0;
		8586: rom = 1'b0;
		8587: rom = 1'b0;
		8588: rom = 1'b0;
		8589: rom = 1'b0;
		8590: rom = 1'b0;
		8591: rom = 1'b0;
		8592: rom = 1'b0;
		8593: rom = 1'b0;
		8594: rom = 1'b0;
		8595: rom = 1'b0;
		8596: rom = 1'b0;
		8597: rom = 1'b0;
		8598: rom = 1'b0;
		8599: rom = 1'b0;
		8600: rom = 1'b0;
		8601: rom = 1'b0;
		8602: rom = 1'b0;
		8603: rom = 1'b0;
		8604: rom = 1'b0;
		8605: rom = 1'b0;
		8606: rom = 1'b0;
		8607: rom = 1'b0;
		8608: rom = 1'b0;
		8609: rom = 1'b0;
		8610: rom = 1'b1;
		8611: rom = 1'b1;
		8612: rom = 1'b1;
		8613: rom = 1'b1;
		8614: rom = 1'b1;
		8615: rom = 1'b1;
		8616: rom = 1'b1;
		8617: rom = 1'b1;
		8618: rom = 1'b1;
		8619: rom = 1'b1;
		8620: rom = 1'b1;
		8621: rom = 1'b1;
		8622: rom = 1'b1;
		8623: rom = 1'b1;
		8624: rom = 1'b1;
		8625: rom = 1'b1;
		8626: rom = 1'b1;
		8627: rom = 1'b1;
		8628: rom = 1'b1;
		8629: rom = 1'b1;
		8630: rom = 1'b0;
		8631: rom = 1'b0;
		8632: rom = 1'b1;
		8633: rom = 1'b1;
		8634: rom = 1'b1;
		8635: rom = 1'b1;
		8636: rom = 1'b1;
		8637: rom = 1'b1;
		8638: rom = 1'b1;
		8639: rom = 1'b1;
		8640: rom = 1'b1;
		8641: rom = 1'b1;
		8642: rom = 1'b1;
		8643: rom = 1'b1;
		8644: rom = 1'b1;
		8645: rom = 1'b1;
		8646: rom = 1'b1;
		8647: rom = 1'b1;
		8648: rom = 1'b1;
		8649: rom = 1'b1;
		8650: rom = 1'b1;
		8651: rom = 1'b1;
		8652: rom = 1'b1;
		8653: rom = 1'b1;
		8654: rom = 1'b1;
		8655: rom = 1'b1;
		8656: rom = 1'b1;
		8657: rom = 1'b1;
		8658: rom = 1'b1;
		8659: rom = 1'b1;
		8660: rom = 1'b1;
		8661: rom = 1'b1;
		8662: rom = 1'b1;
		8663: rom = 1'b1;
		8664: rom = 1'b1;
		8665: rom = 1'b1;
		8666: rom = 1'b1;
		8667: rom = 1'b1;
		8668: rom = 1'b1;
		8669: rom = 1'b1;
		8670: rom = 1'b0;
		8671: rom = 1'b1;
		8672: rom = 1'b1;
		8673: rom = 1'b1;
		8674: rom = 1'b1;
		8675: rom = 1'b1;
		8676: rom = 1'b1;
		8677: rom = 1'b1;
		8678: rom = 1'b1;
		8679: rom = 1'b1;
		8680: rom = 1'b1;
		8681: rom = 1'b1;
		8682: rom = 1'b1;
		8683: rom = 1'b1;
		8684: rom = 1'b1;
		8685: rom = 1'b1;
		8686: rom = 1'b1;
		8687: rom = 1'b1;
		8688: rom = 1'b1;
		8689: rom = 1'b1;
		8690: rom = 1'b1;
		8691: rom = 1'b1;
		8692: rom = 1'b1;
		8693: rom = 1'b0;
		8694: rom = 1'b0;
		8695: rom = 1'b0;
		8696: rom = 1'b0;
		8697: rom = 1'b0;
		8698: rom = 1'b0;
		8699: rom = 1'b0;
		8700: rom = 1'b0;
		8701: rom = 1'b0;
		8702: rom = 1'b0;
		8703: rom = 1'b0;
		8704: rom = 1'b0;
		8705: rom = 1'b0;
		8706: rom = 1'b0;
		8707: rom = 1'b0;
		8708: rom = 1'b0;
		8709: rom = 1'b0;
		8710: rom = 1'b0;
		8711: rom = 1'b0;
		8712: rom = 1'b0;
		8713: rom = 1'b0;
		8714: rom = 1'b0;
		8715: rom = 1'b0;
		8716: rom = 1'b0;
		8717: rom = 1'b0;
		8718: rom = 1'b0;
		8719: rom = 1'b0;
		8720: rom = 1'b0;
		8721: rom = 1'b0;
		8722: rom = 1'b0;
		8723: rom = 1'b0;
		8724: rom = 1'b0;
		8725: rom = 1'b0;
		8726: rom = 1'b0;
		8727: rom = 1'b0;
		8728: rom = 1'b0;
		8729: rom = 1'b0;
		8730: rom = 1'b0;
		8731: rom = 1'b0;
		8732: rom = 1'b0;
		8733: rom = 1'b0;
		8734: rom = 1'b0;
		8735: rom = 1'b0;
		8736: rom = 1'b0;
		8737: rom = 1'b0;
		8738: rom = 1'b1;
		8739: rom = 1'b1;
		8740: rom = 1'b1;
		8741: rom = 1'b1;
		8742: rom = 1'b1;
		8743: rom = 1'b1;
		8744: rom = 1'b1;
		8745: rom = 1'b1;
		8746: rom = 1'b1;
		8747: rom = 1'b1;
		8748: rom = 1'b1;
		8749: rom = 1'b1;
		8750: rom = 1'b1;
		8751: rom = 1'b1;
		8752: rom = 1'b1;
		8753: rom = 1'b1;
		8754: rom = 1'b1;
		8755: rom = 1'b1;
		8756: rom = 1'b1;
		8757: rom = 1'b1;
		8758: rom = 1'b0;
		8759: rom = 1'b1;
		8760: rom = 1'b1;
		8761: rom = 1'b1;
		8762: rom = 1'b1;
		8763: rom = 1'b1;
		8764: rom = 1'b1;
		8765: rom = 1'b1;
		8766: rom = 1'b1;
		8767: rom = 1'b1;
		8768: rom = 1'b1;
		8769: rom = 1'b1;
		8770: rom = 1'b1;
		8771: rom = 1'b1;
		8772: rom = 1'b1;
		8773: rom = 1'b1;
		8774: rom = 1'b1;
		8775: rom = 1'b1;
		8776: rom = 1'b1;
		8777: rom = 1'b1;
		8778: rom = 1'b1;
		8779: rom = 1'b1;
		8780: rom = 1'b1;
		8781: rom = 1'b1;
		8782: rom = 1'b1;
		8783: rom = 1'b1;
		8784: rom = 1'b1;
		8785: rom = 1'b1;
		8786: rom = 1'b1;
		8787: rom = 1'b1;
		8788: rom = 1'b1;
		8789: rom = 1'b1;
		8790: rom = 1'b1;
		8791: rom = 1'b1;
		8792: rom = 1'b1;
		8793: rom = 1'b1;
		8794: rom = 1'b1;
		8795: rom = 1'b1;
		8796: rom = 1'b1;
		8797: rom = 1'b1;
		8798: rom = 1'b0;
		8799: rom = 1'b1;
		8800: rom = 1'b1;
		8801: rom = 1'b1;
		8802: rom = 1'b1;
		8803: rom = 1'b1;
		8804: rom = 1'b1;
		8805: rom = 1'b1;
		8806: rom = 1'b1;
		8807: rom = 1'b1;
		8808: rom = 1'b1;
		8809: rom = 1'b1;
		8810: rom = 1'b1;
		8811: rom = 1'b1;
		8812: rom = 1'b1;
		8813: rom = 1'b1;
		8814: rom = 1'b1;
		8815: rom = 1'b1;
		8816: rom = 1'b1;
		8817: rom = 1'b1;
		8818: rom = 1'b1;
		8819: rom = 1'b1;
		8820: rom = 1'b1;
		8821: rom = 1'b0;
		8822: rom = 1'b0;
		8823: rom = 1'b0;
		8824: rom = 1'b0;
		8825: rom = 1'b0;
		8826: rom = 1'b0;
		8827: rom = 1'b0;
		8828: rom = 1'b0;
		8829: rom = 1'b0;
		8830: rom = 1'b0;
		8831: rom = 1'b0;
		8832: rom = 1'b0;
		8833: rom = 1'b0;
		8834: rom = 1'b0;
		8835: rom = 1'b0;
		8836: rom = 1'b0;
		8837: rom = 1'b0;
		8838: rom = 1'b0;
		8839: rom = 1'b0;
		8840: rom = 1'b0;
		8841: rom = 1'b0;
		8842: rom = 1'b0;
		8843: rom = 1'b0;
		8844: rom = 1'b0;
		8845: rom = 1'b0;
		8846: rom = 1'b0;
		8847: rom = 1'b0;
		8848: rom = 1'b0;
		8849: rom = 1'b0;
		8850: rom = 1'b0;
		8851: rom = 1'b0;
		8852: rom = 1'b0;
		8853: rom = 1'b0;
		8854: rom = 1'b0;
		8855: rom = 1'b0;
		8856: rom = 1'b0;
		8857: rom = 1'b0;
		8858: rom = 1'b0;
		8859: rom = 1'b0;
		8860: rom = 1'b0;
		8861: rom = 1'b0;
		8862: rom = 1'b0;
		8863: rom = 1'b0;
		8864: rom = 1'b0;
		8865: rom = 1'b0;
		8866: rom = 1'b1;
		8867: rom = 1'b1;
		8868: rom = 1'b1;
		8869: rom = 1'b1;
		8870: rom = 1'b1;
		8871: rom = 1'b1;
		8872: rom = 1'b1;
		8873: rom = 1'b1;
		8874: rom = 1'b1;
		8875: rom = 1'b1;
		8876: rom = 1'b1;
		8877: rom = 1'b1;
		8878: rom = 1'b1;
		8879: rom = 1'b1;
		8880: rom = 1'b1;
		8881: rom = 1'b1;
		8882: rom = 1'b1;
		8883: rom = 1'b1;
		8884: rom = 1'b1;
		8885: rom = 1'b1;
		8886: rom = 1'b0;
		8887: rom = 1'b1;
		8888: rom = 1'b1;
		8889: rom = 1'b1;
		8890: rom = 1'b1;
		8891: rom = 1'b1;
		8892: rom = 1'b1;
		8893: rom = 1'b1;
		8894: rom = 1'b1;
		8895: rom = 1'b1;
		8896: rom = 1'b1;
		8897: rom = 1'b1;
		8898: rom = 1'b1;
		8899: rom = 1'b1;
		8900: rom = 1'b1;
		8901: rom = 1'b1;
		8902: rom = 1'b1;
		8903: rom = 1'b1;
		8904: rom = 1'b1;
		8905: rom = 1'b1;
		8906: rom = 1'b1;
		8907: rom = 1'b1;
		8908: rom = 1'b1;
		8909: rom = 1'b1;
		8910: rom = 1'b1;
		8911: rom = 1'b1;
		8912: rom = 1'b1;
		8913: rom = 1'b1;
		8914: rom = 1'b1;
		8915: rom = 1'b1;
		8916: rom = 1'b1;
		8917: rom = 1'b1;
		8918: rom = 1'b1;
		8919: rom = 1'b1;
		8920: rom = 1'b1;
		8921: rom = 1'b1;
		8922: rom = 1'b1;
		8923: rom = 1'b1;
		8924: rom = 1'b1;
		8925: rom = 1'b0;
		8926: rom = 1'b1;
		8927: rom = 1'b1;
		8928: rom = 1'b1;
		8929: rom = 1'b1;
		8930: rom = 1'b1;
		8931: rom = 1'b1;
		8932: rom = 1'b1;
		8933: rom = 1'b1;
		8934: rom = 1'b1;
		8935: rom = 1'b1;
		8936: rom = 1'b1;
		8937: rom = 1'b1;
		8938: rom = 1'b1;
		8939: rom = 1'b1;
		8940: rom = 1'b1;
		8941: rom = 1'b1;
		8942: rom = 1'b1;
		8943: rom = 1'b1;
		8944: rom = 1'b1;
		8945: rom = 1'b1;
		8946: rom = 1'b1;
		8947: rom = 1'b1;
		8948: rom = 1'b1;
		8949: rom = 1'b0;
		8950: rom = 1'b0;
		8951: rom = 1'b0;
		8952: rom = 1'b0;
		8953: rom = 1'b0;
		8954: rom = 1'b0;
		8955: rom = 1'b0;
		8956: rom = 1'b0;
		8957: rom = 1'b0;
		8958: rom = 1'b0;
		8959: rom = 1'b0;
		8960: rom = 1'b0;
		8961: rom = 1'b0;
		8962: rom = 1'b0;
		8963: rom = 1'b0;
		8964: rom = 1'b0;
		8965: rom = 1'b0;
		8966: rom = 1'b0;
		8967: rom = 1'b0;
		8968: rom = 1'b0;
		8969: rom = 1'b0;
		8970: rom = 1'b0;
		8971: rom = 1'b0;
		8972: rom = 1'b0;
		8973: rom = 1'b0;
		8974: rom = 1'b0;
		8975: rom = 1'b0;
		8976: rom = 1'b0;
		8977: rom = 1'b0;
		8978: rom = 1'b0;
		8979: rom = 1'b0;
		8980: rom = 1'b0;
		8981: rom = 1'b0;
		8982: rom = 1'b0;
		8983: rom = 1'b0;
		8984: rom = 1'b0;
		8985: rom = 1'b0;
		8986: rom = 1'b0;
		8987: rom = 1'b0;
		8988: rom = 1'b0;
		8989: rom = 1'b0;
		8990: rom = 1'b0;
		8991: rom = 1'b0;
		8992: rom = 1'b0;
		8993: rom = 1'b0;
		8994: rom = 1'b1;
		8995: rom = 1'b1;
		8996: rom = 1'b1;
		8997: rom = 1'b1;
		8998: rom = 1'b1;
		8999: rom = 1'b1;
		9000: rom = 1'b1;
		9001: rom = 1'b1;
		9002: rom = 1'b1;
		9003: rom = 1'b1;
		9004: rom = 1'b1;
		9005: rom = 1'b1;
		9006: rom = 1'b1;
		9007: rom = 1'b1;
		9008: rom = 1'b1;
		9009: rom = 1'b1;
		9010: rom = 1'b1;
		9011: rom = 1'b1;
		9012: rom = 1'b1;
		9013: rom = 1'b0;
		9014: rom = 1'b1;
		9015: rom = 1'b1;
		9016: rom = 1'b1;
		9017: rom = 1'b1;
		9018: rom = 1'b1;
		9019: rom = 1'b1;
		9020: rom = 1'b1;
		9021: rom = 1'b1;
		9022: rom = 1'b1;
		9023: rom = 1'b1;
		9024: rom = 1'b1;
		9025: rom = 1'b1;
		9026: rom = 1'b1;
		9027: rom = 1'b1;
		9028: rom = 1'b1;
		9029: rom = 1'b1;
		9030: rom = 1'b1;
		9031: rom = 1'b1;
		9032: rom = 1'b1;
		9033: rom = 1'b1;
		9034: rom = 1'b1;
		9035: rom = 1'b1;
		9036: rom = 1'b1;
		9037: rom = 1'b1;
		9038: rom = 1'b1;
		9039: rom = 1'b1;
		9040: rom = 1'b1;
		9041: rom = 1'b1;
		9042: rom = 1'b1;
		9043: rom = 1'b1;
		9044: rom = 1'b1;
		9045: rom = 1'b1;
		9046: rom = 1'b1;
		9047: rom = 1'b1;
		9048: rom = 1'b1;
		9049: rom = 1'b1;
		9050: rom = 1'b1;
		9051: rom = 1'b1;
		9052: rom = 1'b0;
		9053: rom = 1'b0;
		9054: rom = 1'b1;
		9055: rom = 1'b1;
		9056: rom = 1'b1;
		9057: rom = 1'b1;
		9058: rom = 1'b1;
		9059: rom = 1'b1;
		9060: rom = 1'b1;
		9061: rom = 1'b1;
		9062: rom = 1'b1;
		9063: rom = 1'b1;
		9064: rom = 1'b1;
		9065: rom = 1'b1;
		9066: rom = 1'b1;
		9067: rom = 1'b1;
		9068: rom = 1'b1;
		9069: rom = 1'b1;
		9070: rom = 1'b1;
		9071: rom = 1'b1;
		9072: rom = 1'b1;
		9073: rom = 1'b1;
		9074: rom = 1'b1;
		9075: rom = 1'b1;
		9076: rom = 1'b1;
		9077: rom = 1'b0;
		9078: rom = 1'b0;
		9079: rom = 1'b0;
		9080: rom = 1'b0;
		9081: rom = 1'b0;
		9082: rom = 1'b0;
		9083: rom = 1'b0;
		9084: rom = 1'b0;
		9085: rom = 1'b0;
		9086: rom = 1'b0;
		9087: rom = 1'b0;
		9088: rom = 1'b0;
		9089: rom = 1'b0;
		9090: rom = 1'b0;
		9091: rom = 1'b0;
		9092: rom = 1'b0;
		9093: rom = 1'b0;
		9094: rom = 1'b0;
		9095: rom = 1'b0;
		9096: rom = 1'b0;
		9097: rom = 1'b0;
		9098: rom = 1'b0;
		9099: rom = 1'b0;
		9100: rom = 1'b0;
		9101: rom = 1'b0;
		9102: rom = 1'b0;
		9103: rom = 1'b0;
		9104: rom = 1'b0;
		9105: rom = 1'b0;
		9106: rom = 1'b0;
		9107: rom = 1'b0;
		9108: rom = 1'b0;
		9109: rom = 1'b0;
		9110: rom = 1'b0;
		9111: rom = 1'b0;
		9112: rom = 1'b0;
		9113: rom = 1'b0;
		9114: rom = 1'b0;
		9115: rom = 1'b0;
		9116: rom = 1'b0;
		9117: rom = 1'b0;
		9118: rom = 1'b0;
		9119: rom = 1'b0;
		9120: rom = 1'b0;
		9121: rom = 1'b1;
		9122: rom = 1'b1;
		9123: rom = 1'b1;
		9124: rom = 1'b1;
		9125: rom = 1'b1;
		9126: rom = 1'b1;
		9127: rom = 1'b1;
		9128: rom = 1'b1;
		9129: rom = 1'b1;
		9130: rom = 1'b1;
		9131: rom = 1'b1;
		9132: rom = 1'b1;
		9133: rom = 1'b1;
		9134: rom = 1'b1;
		9135: rom = 1'b1;
		9136: rom = 1'b1;
		9137: rom = 1'b1;
		9138: rom = 1'b1;
		9139: rom = 1'b1;
		9140: rom = 1'b1;
		9141: rom = 1'b0;
		9142: rom = 1'b1;
		9143: rom = 1'b1;
		9144: rom = 1'b1;
		9145: rom = 1'b1;
		9146: rom = 1'b1;
		9147: rom = 1'b1;
		9148: rom = 1'b1;
		9149: rom = 1'b1;
		9150: rom = 1'b1;
		9151: rom = 1'b1;
		9152: rom = 1'b1;
		9153: rom = 1'b1;
		9154: rom = 1'b1;
		9155: rom = 1'b1;
		9156: rom = 1'b1;
		9157: rom = 1'b1;
		9158: rom = 1'b1;
		9159: rom = 1'b1;
		9160: rom = 1'b1;
		9161: rom = 1'b1;
		9162: rom = 1'b1;
		9163: rom = 1'b1;
		9164: rom = 1'b1;
		9165: rom = 1'b1;
		9166: rom = 1'b1;
		9167: rom = 1'b1;
		9168: rom = 1'b1;
		9169: rom = 1'b1;
		9170: rom = 1'b1;
		9171: rom = 1'b1;
		9172: rom = 1'b1;
		9173: rom = 1'b1;
		9174: rom = 1'b1;
		9175: rom = 1'b1;
		9176: rom = 1'b1;
		9177: rom = 1'b1;
		9178: rom = 1'b1;
		9179: rom = 1'b1;
		9180: rom = 1'b0;
		9181: rom = 1'b1;
		9182: rom = 1'b1;
		9183: rom = 1'b1;
		9184: rom = 1'b1;
		9185: rom = 1'b1;
		9186: rom = 1'b1;
		9187: rom = 1'b1;
		9188: rom = 1'b1;
		9189: rom = 1'b1;
		9190: rom = 1'b1;
		9191: rom = 1'b1;
		9192: rom = 1'b1;
		9193: rom = 1'b1;
		9194: rom = 1'b1;
		9195: rom = 1'b1;
		9196: rom = 1'b1;
		9197: rom = 1'b1;
		9198: rom = 1'b1;
		9199: rom = 1'b1;
		9200: rom = 1'b1;
		9201: rom = 1'b1;
		9202: rom = 1'b1;
		9203: rom = 1'b1;
		9204: rom = 1'b0;
		9205: rom = 1'b0;
		9206: rom = 1'b0;
		9207: rom = 1'b0;
		9208: rom = 1'b0;
		9209: rom = 1'b0;
		9210: rom = 1'b0;
		9211: rom = 1'b0;
		9212: rom = 1'b0;
		9213: rom = 1'b0;
		9214: rom = 1'b0;
		9215: rom = 1'b0;
		9216: rom = 1'b0;
		9217: rom = 1'b0;
		9218: rom = 1'b0;
		9219: rom = 1'b0;
		9220: rom = 1'b0;
		9221: rom = 1'b0;
		9222: rom = 1'b0;
		9223: rom = 1'b0;
		9224: rom = 1'b0;
		9225: rom = 1'b0;
		9226: rom = 1'b0;
		9227: rom = 1'b0;
		9228: rom = 1'b0;
		9229: rom = 1'b0;
		9230: rom = 1'b0;
		9231: rom = 1'b0;
		9232: rom = 1'b0;
		9233: rom = 1'b0;
		9234: rom = 1'b0;
		9235: rom = 1'b0;
		9236: rom = 1'b0;
		9237: rom = 1'b0;
		9238: rom = 1'b0;
		9239: rom = 1'b0;
		9240: rom = 1'b0;
		9241: rom = 1'b0;
		9242: rom = 1'b0;
		9243: rom = 1'b0;
		9244: rom = 1'b0;
		9245: rom = 1'b0;
		9246: rom = 1'b0;
		9247: rom = 1'b0;
		9248: rom = 1'b0;
		9249: rom = 1'b0;
		9250: rom = 1'b1;
		9251: rom = 1'b1;
		9252: rom = 1'b1;
		9253: rom = 1'b1;
		9254: rom = 1'b1;
		9255: rom = 1'b1;
		9256: rom = 1'b1;
		9257: rom = 1'b1;
		9258: rom = 1'b1;
		9259: rom = 1'b1;
		9260: rom = 1'b1;
		9261: rom = 1'b1;
		9262: rom = 1'b1;
		9263: rom = 1'b1;
		9264: rom = 1'b1;
		9265: rom = 1'b1;
		9266: rom = 1'b1;
		9267: rom = 1'b1;
		9268: rom = 1'b0;
		9269: rom = 1'b0;
		9270: rom = 1'b1;
		9271: rom = 1'b1;
		9272: rom = 1'b1;
		9273: rom = 1'b1;
		9274: rom = 1'b1;
		9275: rom = 1'b1;
		9276: rom = 1'b1;
		9277: rom = 1'b1;
		9278: rom = 1'b1;
		9279: rom = 1'b1;
		9280: rom = 1'b1;
		9281: rom = 1'b1;
		9282: rom = 1'b1;
		9283: rom = 1'b1;
		9284: rom = 1'b1;
		9285: rom = 1'b1;
		9286: rom = 1'b1;
		9287: rom = 1'b1;
		9288: rom = 1'b1;
		9289: rom = 1'b1;
		9290: rom = 1'b1;
		9291: rom = 1'b1;
		9292: rom = 1'b1;
		9293: rom = 1'b1;
		9294: rom = 1'b1;
		9295: rom = 1'b1;
		9296: rom = 1'b1;
		9297: rom = 1'b1;
		9298: rom = 1'b1;
		9299: rom = 1'b1;
		9300: rom = 1'b1;
		9301: rom = 1'b1;
		9302: rom = 1'b1;
		9303: rom = 1'b1;
		9304: rom = 1'b1;
		9305: rom = 1'b1;
		9306: rom = 1'b1;
		9307: rom = 1'b0;
		9308: rom = 1'b1;
		9309: rom = 1'b1;
		9310: rom = 1'b1;
		9311: rom = 1'b1;
		9312: rom = 1'b1;
		9313: rom = 1'b1;
		9314: rom = 1'b1;
		9315: rom = 1'b1;
		9316: rom = 1'b1;
		9317: rom = 1'b1;
		9318: rom = 1'b1;
		9319: rom = 1'b1;
		9320: rom = 1'b1;
		9321: rom = 1'b1;
		9322: rom = 1'b1;
		9323: rom = 1'b1;
		9324: rom = 1'b1;
		9325: rom = 1'b1;
		9326: rom = 1'b1;
		9327: rom = 1'b1;
		9328: rom = 1'b1;
		9329: rom = 1'b1;
		9330: rom = 1'b1;
		9331: rom = 1'b1;
		9332: rom = 1'b0;
		9333: rom = 1'b0;
		9334: rom = 1'b0;
		9335: rom = 1'b0;
		9336: rom = 1'b0;
		9337: rom = 1'b0;
		9338: rom = 1'b0;
		9339: rom = 1'b0;
		9340: rom = 1'b0;
		9341: rom = 1'b0;
		9342: rom = 1'b0;
		9343: rom = 1'b0;
		9344: rom = 1'b0;
		9345: rom = 1'b0;
		9346: rom = 1'b0;
		9347: rom = 1'b0;
		9348: rom = 1'b0;
		9349: rom = 1'b0;
		9350: rom = 1'b0;
		9351: rom = 1'b0;
		9352: rom = 1'b0;
		9353: rom = 1'b0;
		9354: rom = 1'b0;
		9355: rom = 1'b0;
		9356: rom = 1'b0;
		9357: rom = 1'b0;
		9358: rom = 1'b0;
		9359: rom = 1'b0;
		9360: rom = 1'b0;
		9361: rom = 1'b0;
		9362: rom = 1'b0;
		9363: rom = 1'b0;
		9364: rom = 1'b0;
		9365: rom = 1'b0;
		9366: rom = 1'b0;
		9367: rom = 1'b0;
		9368: rom = 1'b0;
		9369: rom = 1'b0;
		9370: rom = 1'b0;
		9371: rom = 1'b0;
		9372: rom = 1'b0;
		9373: rom = 1'b0;
		9374: rom = 1'b0;
		9375: rom = 1'b0;
		9376: rom = 1'b0;
		9377: rom = 1'b0;
		9378: rom = 1'b1;
		9379: rom = 1'b1;
		9380: rom = 1'b1;
		9381: rom = 1'b1;
		9382: rom = 1'b1;
		9383: rom = 1'b1;
		9384: rom = 1'b1;
		9385: rom = 1'b1;
		9386: rom = 1'b1;
		9387: rom = 1'b1;
		9388: rom = 1'b1;
		9389: rom = 1'b1;
		9390: rom = 1'b1;
		9391: rom = 1'b1;
		9392: rom = 1'b1;
		9393: rom = 1'b1;
		9394: rom = 1'b1;
		9395: rom = 1'b1;
		9396: rom = 1'b0;
		9397: rom = 1'b1;
		9398: rom = 1'b1;
		9399: rom = 1'b1;
		9400: rom = 1'b1;
		9401: rom = 1'b1;
		9402: rom = 1'b1;
		9403: rom = 1'b1;
		9404: rom = 1'b1;
		9405: rom = 1'b1;
		9406: rom = 1'b1;
		9407: rom = 1'b1;
		9408: rom = 1'b1;
		9409: rom = 1'b1;
		9410: rom = 1'b1;
		9411: rom = 1'b1;
		9412: rom = 1'b1;
		9413: rom = 1'b1;
		9414: rom = 1'b1;
		9415: rom = 1'b1;
		9416: rom = 1'b1;
		9417: rom = 1'b1;
		9418: rom = 1'b1;
		9419: rom = 1'b1;
		9420: rom = 1'b1;
		9421: rom = 1'b1;
		9422: rom = 1'b1;
		9423: rom = 1'b1;
		9424: rom = 1'b1;
		9425: rom = 1'b1;
		9426: rom = 1'b1;
		9427: rom = 1'b1;
		9428: rom = 1'b1;
		9429: rom = 1'b1;
		9430: rom = 1'b1;
		9431: rom = 1'b1;
		9432: rom = 1'b1;
		9433: rom = 1'b1;
		9434: rom = 1'b0;
		9435: rom = 1'b0;
		9436: rom = 1'b1;
		9437: rom = 1'b1;
		9438: rom = 1'b1;
		9439: rom = 1'b1;
		9440: rom = 1'b1;
		9441: rom = 1'b1;
		9442: rom = 1'b1;
		9443: rom = 1'b1;
		9444: rom = 1'b1;
		9445: rom = 1'b1;
		9446: rom = 1'b1;
		9447: rom = 1'b1;
		9448: rom = 1'b1;
		9449: rom = 1'b1;
		9450: rom = 1'b1;
		9451: rom = 1'b1;
		9452: rom = 1'b1;
		9453: rom = 1'b1;
		9454: rom = 1'b1;
		9455: rom = 1'b1;
		9456: rom = 1'b1;
		9457: rom = 1'b1;
		9458: rom = 1'b1;
		9459: rom = 1'b1;
		9460: rom = 1'b0;
		9461: rom = 1'b0;
		9462: rom = 1'b0;
		9463: rom = 1'b0;
		9464: rom = 1'b0;
		9465: rom = 1'b0;
		9466: rom = 1'b0;
		9467: rom = 1'b0;
		9468: rom = 1'b0;
		9469: rom = 1'b0;
		9470: rom = 1'b0;
		9471: rom = 1'b0;
		9472: rom = 1'b0;
		9473: rom = 1'b0;
		9474: rom = 1'b0;
		9475: rom = 1'b0;
		9476: rom = 1'b0;
		9477: rom = 1'b0;
		9478: rom = 1'b0;
		9479: rom = 1'b0;
		9480: rom = 1'b0;
		9481: rom = 1'b0;
		9482: rom = 1'b0;
		9483: rom = 1'b0;
		9484: rom = 1'b0;
		9485: rom = 1'b0;
		9486: rom = 1'b0;
		9487: rom = 1'b0;
		9488: rom = 1'b0;
		9489: rom = 1'b0;
		9490: rom = 1'b0;
		9491: rom = 1'b0;
		9492: rom = 1'b0;
		9493: rom = 1'b0;
		9494: rom = 1'b0;
		9495: rom = 1'b0;
		9496: rom = 1'b0;
		9497: rom = 1'b0;
		9498: rom = 1'b0;
		9499: rom = 1'b0;
		9500: rom = 1'b0;
		9501: rom = 1'b0;
		9502: rom = 1'b0;
		9503: rom = 1'b0;
		9504: rom = 1'b0;
		9505: rom = 1'b0;
		9506: rom = 1'b0;
		9507: rom = 1'b1;
		9508: rom = 1'b1;
		9509: rom = 1'b1;
		9510: rom = 1'b1;
		9511: rom = 1'b1;
		9512: rom = 1'b1;
		9513: rom = 1'b1;
		9514: rom = 1'b1;
		9515: rom = 1'b1;
		9516: rom = 1'b1;
		9517: rom = 1'b1;
		9518: rom = 1'b1;
		9519: rom = 1'b1;
		9520: rom = 1'b1;
		9521: rom = 1'b1;
		9522: rom = 1'b1;
		9523: rom = 1'b1;
		9524: rom = 1'b0;
		9525: rom = 1'b1;
		9526: rom = 1'b1;
		9527: rom = 1'b1;
		9528: rom = 1'b1;
		9529: rom = 1'b1;
		9530: rom = 1'b1;
		9531: rom = 1'b1;
		9532: rom = 1'b1;
		9533: rom = 1'b1;
		9534: rom = 1'b1;
		9535: rom = 1'b1;
		9536: rom = 1'b1;
		9537: rom = 1'b1;
		9538: rom = 1'b1;
		9539: rom = 1'b1;
		9540: rom = 1'b1;
		9541: rom = 1'b1;
		9542: rom = 1'b1;
		9543: rom = 1'b1;
		9544: rom = 1'b1;
		9545: rom = 1'b1;
		9546: rom = 1'b1;
		9547: rom = 1'b1;
		9548: rom = 1'b1;
		9549: rom = 1'b1;
		9550: rom = 1'b1;
		9551: rom = 1'b1;
		9552: rom = 1'b1;
		9553: rom = 1'b1;
		9554: rom = 1'b1;
		9555: rom = 1'b1;
		9556: rom = 1'b1;
		9557: rom = 1'b1;
		9558: rom = 1'b1;
		9559: rom = 1'b1;
		9560: rom = 1'b1;
		9561: rom = 1'b0;
		9562: rom = 1'b0;
		9563: rom = 1'b1;
		9564: rom = 1'b1;
		9565: rom = 1'b1;
		9566: rom = 1'b1;
		9567: rom = 1'b1;
		9568: rom = 1'b1;
		9569: rom = 1'b1;
		9570: rom = 1'b1;
		9571: rom = 1'b1;
		9572: rom = 1'b1;
		9573: rom = 1'b1;
		9574: rom = 1'b1;
		9575: rom = 1'b1;
		9576: rom = 1'b1;
		9577: rom = 1'b1;
		9578: rom = 1'b1;
		9579: rom = 1'b1;
		9580: rom = 1'b1;
		9581: rom = 1'b1;
		9582: rom = 1'b1;
		9583: rom = 1'b1;
		9584: rom = 1'b1;
		9585: rom = 1'b1;
		9586: rom = 1'b1;
		9587: rom = 1'b1;
		9588: rom = 1'b0;
		9589: rom = 1'b0;
		9590: rom = 1'b0;
		9591: rom = 1'b0;
		9592: rom = 1'b0;
		9593: rom = 1'b0;
		9594: rom = 1'b0;
		9595: rom = 1'b0;
		9596: rom = 1'b0;
		9597: rom = 1'b0;
		9598: rom = 1'b0;
		9599: rom = 1'b0;
		9600: rom = 1'b0;
		9601: rom = 1'b0;
		9602: rom = 1'b0;
		9603: rom = 1'b0;
		9604: rom = 1'b0;
		9605: rom = 1'b0;
		9606: rom = 1'b0;
		9607: rom = 1'b0;
		9608: rom = 1'b0;
		9609: rom = 1'b0;
		9610: rom = 1'b0;
		9611: rom = 1'b0;
		9612: rom = 1'b0;
		9613: rom = 1'b0;
		9614: rom = 1'b0;
		9615: rom = 1'b0;
		9616: rom = 1'b0;
		9617: rom = 1'b0;
		9618: rom = 1'b0;
		9619: rom = 1'b0;
		9620: rom = 1'b0;
		9621: rom = 1'b0;
		9622: rom = 1'b0;
		9623: rom = 1'b0;
		9624: rom = 1'b0;
		9625: rom = 1'b0;
		9626: rom = 1'b0;
		9627: rom = 1'b0;
		9628: rom = 1'b0;
		9629: rom = 1'b0;
		9630: rom = 1'b0;
		9631: rom = 1'b0;
		9632: rom = 1'b0;
		9633: rom = 1'b0;
		9634: rom = 1'b0;
		9635: rom = 1'b1;
		9636: rom = 1'b1;
		9637: rom = 1'b1;
		9638: rom = 1'b1;
		9639: rom = 1'b1;
		9640: rom = 1'b1;
		9641: rom = 1'b1;
		9642: rom = 1'b1;
		9643: rom = 1'b1;
		9644: rom = 1'b1;
		9645: rom = 1'b1;
		9646: rom = 1'b1;
		9647: rom = 1'b1;
		9648: rom = 1'b1;
		9649: rom = 1'b1;
		9650: rom = 1'b1;
		9651: rom = 1'b1;
		9652: rom = 1'b0;
		9653: rom = 1'b1;
		9654: rom = 1'b1;
		9655: rom = 1'b1;
		9656: rom = 1'b1;
		9657: rom = 1'b1;
		9658: rom = 1'b1;
		9659: rom = 1'b1;
		9660: rom = 1'b1;
		9661: rom = 1'b1;
		9662: rom = 1'b1;
		9663: rom = 1'b1;
		9664: rom = 1'b1;
		9665: rom = 1'b1;
		9666: rom = 1'b1;
		9667: rom = 1'b1;
		9668: rom = 1'b1;
		9669: rom = 1'b1;
		9670: rom = 1'b1;
		9671: rom = 1'b1;
		9672: rom = 1'b1;
		9673: rom = 1'b1;
		9674: rom = 1'b1;
		9675: rom = 1'b1;
		9676: rom = 1'b1;
		9677: rom = 1'b1;
		9678: rom = 1'b1;
		9679: rom = 1'b1;
		9680: rom = 1'b1;
		9681: rom = 1'b1;
		9682: rom = 1'b1;
		9683: rom = 1'b1;
		9684: rom = 1'b1;
		9685: rom = 1'b1;
		9686: rom = 1'b1;
		9687: rom = 1'b1;
		9688: rom = 1'b1;
		9689: rom = 1'b0;
		9690: rom = 1'b0;
		9691: rom = 1'b1;
		9692: rom = 1'b1;
		9693: rom = 1'b1;
		9694: rom = 1'b1;
		9695: rom = 1'b1;
		9696: rom = 1'b1;
		9697: rom = 1'b1;
		9698: rom = 1'b1;
		9699: rom = 1'b1;
		9700: rom = 1'b1;
		9701: rom = 1'b1;
		9702: rom = 1'b1;
		9703: rom = 1'b1;
		9704: rom = 1'b1;
		9705: rom = 1'b1;
		9706: rom = 1'b1;
		9707: rom = 1'b1;
		9708: rom = 1'b1;
		9709: rom = 1'b1;
		9710: rom = 1'b1;
		9711: rom = 1'b1;
		9712: rom = 1'b1;
		9713: rom = 1'b1;
		9714: rom = 1'b1;
		9715: rom = 1'b0;
		9716: rom = 1'b0;
		9717: rom = 1'b0;
		9718: rom = 1'b0;
		9719: rom = 1'b0;
		9720: rom = 1'b0;
		9721: rom = 1'b0;
		9722: rom = 1'b0;
		9723: rom = 1'b0;
		9724: rom = 1'b0;
		9725: rom = 1'b0;
		9726: rom = 1'b0;
		9727: rom = 1'b0;
		9728: rom = 1'b0;
		9729: rom = 1'b0;
		9730: rom = 1'b0;
		9731: rom = 1'b0;
		9732: rom = 1'b0;
		9733: rom = 1'b0;
		9734: rom = 1'b0;
		9735: rom = 1'b0;
		9736: rom = 1'b0;
		9737: rom = 1'b0;
		9738: rom = 1'b0;
		9739: rom = 1'b0;
		9740: rom = 1'b0;
		9741: rom = 1'b0;
		9742: rom = 1'b0;
		9743: rom = 1'b0;
		9744: rom = 1'b0;
		9745: rom = 1'b0;
		9746: rom = 1'b0;
		9747: rom = 1'b0;
		9748: rom = 1'b0;
		9749: rom = 1'b0;
		9750: rom = 1'b0;
		9751: rom = 1'b0;
		9752: rom = 1'b0;
		9753: rom = 1'b0;
		9754: rom = 1'b0;
		9755: rom = 1'b0;
		9756: rom = 1'b0;
		9757: rom = 1'b0;
		9758: rom = 1'b0;
		9759: rom = 1'b0;
		9760: rom = 1'b0;
		9761: rom = 1'b0;
		9762: rom = 1'b0;
		9763: rom = 1'b0;
		9764: rom = 1'b1;
		9765: rom = 1'b1;
		9766: rom = 1'b1;
		9767: rom = 1'b1;
		9768: rom = 1'b1;
		9769: rom = 1'b1;
		9770: rom = 1'b1;
		9771: rom = 1'b1;
		9772: rom = 1'b1;
		9773: rom = 1'b1;
		9774: rom = 1'b1;
		9775: rom = 1'b1;
		9776: rom = 1'b1;
		9777: rom = 1'b1;
		9778: rom = 1'b1;
		9779: rom = 1'b1;
		9780: rom = 1'b0;
		9781: rom = 1'b1;
		9782: rom = 1'b1;
		9783: rom = 1'b1;
		9784: rom = 1'b1;
		9785: rom = 1'b1;
		9786: rom = 1'b1;
		9787: rom = 1'b1;
		9788: rom = 1'b1;
		9789: rom = 1'b1;
		9790: rom = 1'b1;
		9791: rom = 1'b1;
		9792: rom = 1'b1;
		9793: rom = 1'b1;
		9794: rom = 1'b1;
		9795: rom = 1'b1;
		9796: rom = 1'b1;
		9797: rom = 1'b1;
		9798: rom = 1'b1;
		9799: rom = 1'b1;
		9800: rom = 1'b1;
		9801: rom = 1'b1;
		9802: rom = 1'b1;
		9803: rom = 1'b1;
		9804: rom = 1'b1;
		9805: rom = 1'b1;
		9806: rom = 1'b1;
		9807: rom = 1'b1;
		9808: rom = 1'b1;
		9809: rom = 1'b1;
		9810: rom = 1'b1;
		9811: rom = 1'b1;
		9812: rom = 1'b1;
		9813: rom = 1'b1;
		9814: rom = 1'b1;
		9815: rom = 1'b1;
		9816: rom = 1'b0;
		9817: rom = 1'b0;
		9818: rom = 1'b1;
		9819: rom = 1'b1;
		9820: rom = 1'b1;
		9821: rom = 1'b1;
		9822: rom = 1'b1;
		9823: rom = 1'b1;
		9824: rom = 1'b1;
		9825: rom = 1'b1;
		9826: rom = 1'b1;
		9827: rom = 1'b1;
		9828: rom = 1'b1;
		9829: rom = 1'b1;
		9830: rom = 1'b1;
		9831: rom = 1'b1;
		9832: rom = 1'b1;
		9833: rom = 1'b1;
		9834: rom = 1'b1;
		9835: rom = 1'b1;
		9836: rom = 1'b1;
		9837: rom = 1'b1;
		9838: rom = 1'b1;
		9839: rom = 1'b1;
		9840: rom = 1'b1;
		9841: rom = 1'b1;
		9842: rom = 1'b1;
		9843: rom = 1'b0;
		9844: rom = 1'b0;
		9845: rom = 1'b0;
		9846: rom = 1'b0;
		9847: rom = 1'b0;
		9848: rom = 1'b0;
		9849: rom = 1'b0;
		9850: rom = 1'b0;
		9851: rom = 1'b0;
		9852: rom = 1'b0;
		9853: rom = 1'b0;
		9854: rom = 1'b0;
		9855: rom = 1'b0;
		9856: rom = 1'b0;
		9857: rom = 1'b0;
		9858: rom = 1'b0;
		9859: rom = 1'b0;
		9860: rom = 1'b0;
		9861: rom = 1'b0;
		9862: rom = 1'b0;
		9863: rom = 1'b0;
		9864: rom = 1'b0;
		9865: rom = 1'b0;
		9866: rom = 1'b0;
		9867: rom = 1'b0;
		9868: rom = 1'b0;
		9869: rom = 1'b0;
		9870: rom = 1'b0;
		9871: rom = 1'b0;
		9872: rom = 1'b0;
		9873: rom = 1'b0;
		9874: rom = 1'b0;
		9875: rom = 1'b0;
		9876: rom = 1'b0;
		9877: rom = 1'b0;
		9878: rom = 1'b0;
		9879: rom = 1'b0;
		9880: rom = 1'b0;
		9881: rom = 1'b0;
		9882: rom = 1'b0;
		9883: rom = 1'b0;
		9884: rom = 1'b0;
		9885: rom = 1'b0;
		9886: rom = 1'b0;
		9887: rom = 1'b0;
		9888: rom = 1'b0;
		9889: rom = 1'b0;
		9890: rom = 1'b0;
		9891: rom = 1'b0;
		9892: rom = 1'b0;
		9893: rom = 1'b1;
		9894: rom = 1'b1;
		9895: rom = 1'b1;
		9896: rom = 1'b1;
		9897: rom = 1'b1;
		9898: rom = 1'b1;
		9899: rom = 1'b1;
		9900: rom = 1'b1;
		9901: rom = 1'b1;
		9902: rom = 1'b1;
		9903: rom = 1'b1;
		9904: rom = 1'b1;
		9905: rom = 1'b1;
		9906: rom = 1'b1;
		9907: rom = 1'b0;
		9908: rom = 1'b1;
		9909: rom = 1'b1;
		9910: rom = 1'b1;
		9911: rom = 1'b1;
		9912: rom = 1'b1;
		9913: rom = 1'b1;
		9914: rom = 1'b1;
		9915: rom = 1'b1;
		9916: rom = 1'b1;
		9917: rom = 1'b1;
		9918: rom = 1'b1;
		9919: rom = 1'b1;
		9920: rom = 1'b1;
		9921: rom = 1'b1;
		9922: rom = 1'b1;
		9923: rom = 1'b1;
		9924: rom = 1'b1;
		9925: rom = 1'b1;
		9926: rom = 1'b1;
		9927: rom = 1'b1;
		9928: rom = 1'b1;
		9929: rom = 1'b1;
		9930: rom = 1'b1;
		9931: rom = 1'b1;
		9932: rom = 1'b1;
		9933: rom = 1'b1;
		9934: rom = 1'b1;
		9935: rom = 1'b1;
		9936: rom = 1'b1;
		9937: rom = 1'b1;
		9938: rom = 1'b1;
		9939: rom = 1'b1;
		9940: rom = 1'b1;
		9941: rom = 1'b1;
		9942: rom = 1'b1;
		9943: rom = 1'b1;
		9944: rom = 1'b0;
		9945: rom = 1'b1;
		9946: rom = 1'b1;
		9947: rom = 1'b1;
		9948: rom = 1'b1;
		9949: rom = 1'b1;
		9950: rom = 1'b1;
		9951: rom = 1'b1;
		9952: rom = 1'b1;
		9953: rom = 1'b1;
		9954: rom = 1'b1;
		9955: rom = 1'b1;
		9956: rom = 1'b1;
		9957: rom = 1'b1;
		9958: rom = 1'b1;
		9959: rom = 1'b1;
		9960: rom = 1'b1;
		9961: rom = 1'b1;
		9962: rom = 1'b1;
		9963: rom = 1'b1;
		9964: rom = 1'b1;
		9965: rom = 1'b1;
		9966: rom = 1'b1;
		9967: rom = 1'b1;
		9968: rom = 1'b1;
		9969: rom = 1'b1;
		9970: rom = 1'b1;
		9971: rom = 1'b0;
		9972: rom = 1'b0;
		9973: rom = 1'b0;
		9974: rom = 1'b0;
		9975: rom = 1'b0;
		9976: rom = 1'b0;
		9977: rom = 1'b0;
		9978: rom = 1'b0;
		9979: rom = 1'b0;
		9980: rom = 1'b0;
		9981: rom = 1'b0;
		9982: rom = 1'b0;
		9983: rom = 1'b0;
		9984: rom = 1'b0;
		9985: rom = 1'b0;
		9986: rom = 1'b0;
		9987: rom = 1'b0;
		9988: rom = 1'b0;
		9989: rom = 1'b0;
		9990: rom = 1'b0;
		9991: rom = 1'b0;
		9992: rom = 1'b0;
		9993: rom = 1'b0;
		9994: rom = 1'b0;
		9995: rom = 1'b0;
		9996: rom = 1'b0;
		9997: rom = 1'b0;
		9998: rom = 1'b0;
		9999: rom = 1'b0;
		10000: rom = 1'b0;
		10001: rom = 1'b0;
		10002: rom = 1'b0;
		10003: rom = 1'b0;
		10004: rom = 1'b0;
		10005: rom = 1'b0;
		10006: rom = 1'b0;
		10007: rom = 1'b0;
		10008: rom = 1'b0;
		10009: rom = 1'b0;
		10010: rom = 1'b0;
		10011: rom = 1'b0;
		10012: rom = 1'b0;
		10013: rom = 1'b0;
		10014: rom = 1'b0;
		10015: rom = 1'b0;
		10016: rom = 1'b0;
		10017: rom = 1'b0;
		10018: rom = 1'b0;
		10019: rom = 1'b0;
		10020: rom = 1'b0;
		10021: rom = 1'b0;
		10022: rom = 1'b1;
		10023: rom = 1'b1;
		10024: rom = 1'b1;
		10025: rom = 1'b1;
		10026: rom = 1'b1;
		10027: rom = 1'b1;
		10028: rom = 1'b1;
		10029: rom = 1'b1;
		10030: rom = 1'b1;
		10031: rom = 1'b1;
		10032: rom = 1'b1;
		10033: rom = 1'b1;
		10034: rom = 1'b1;
		10035: rom = 1'b0;
		10036: rom = 1'b1;
		10037: rom = 1'b1;
		10038: rom = 1'b1;
		10039: rom = 1'b1;
		10040: rom = 1'b1;
		10041: rom = 1'b1;
		10042: rom = 1'b1;
		10043: rom = 1'b1;
		10044: rom = 1'b1;
		10045: rom = 1'b1;
		10046: rom = 1'b1;
		10047: rom = 1'b1;
		10048: rom = 1'b1;
		10049: rom = 1'b1;
		10050: rom = 1'b1;
		10051: rom = 1'b1;
		10052: rom = 1'b1;
		10053: rom = 1'b1;
		10054: rom = 1'b1;
		10055: rom = 1'b1;
		10056: rom = 1'b1;
		10057: rom = 1'b1;
		10058: rom = 1'b1;
		10059: rom = 1'b1;
		10060: rom = 1'b1;
		10061: rom = 1'b1;
		10062: rom = 1'b1;
		10063: rom = 1'b1;
		10064: rom = 1'b1;
		10065: rom = 1'b1;
		10066: rom = 1'b1;
		10067: rom = 1'b1;
		10068: rom = 1'b1;
		10069: rom = 1'b1;
		10070: rom = 1'b1;
		10071: rom = 1'b0;
		10072: rom = 1'b1;
		10073: rom = 1'b1;
		10074: rom = 1'b1;
		10075: rom = 1'b1;
		10076: rom = 1'b1;
		10077: rom = 1'b1;
		10078: rom = 1'b1;
		10079: rom = 1'b1;
		10080: rom = 1'b1;
		10081: rom = 1'b1;
		10082: rom = 1'b1;
		10083: rom = 1'b1;
		10084: rom = 1'b1;
		10085: rom = 1'b1;
		10086: rom = 1'b1;
		10087: rom = 1'b1;
		10088: rom = 1'b1;
		10089: rom = 1'b1;
		10090: rom = 1'b1;
		10091: rom = 1'b1;
		10092: rom = 1'b1;
		10093: rom = 1'b1;
		10094: rom = 1'b1;
		10095: rom = 1'b1;
		10096: rom = 1'b1;
		10097: rom = 1'b1;
		10098: rom = 1'b1;
		10099: rom = 1'b0;
		10100: rom = 1'b0;
		10101: rom = 1'b0;
		10102: rom = 1'b0;
		10103: rom = 1'b0;
		10104: rom = 1'b0;
		10105: rom = 1'b0;
		10106: rom = 1'b0;
		10107: rom = 1'b0;
		10108: rom = 1'b0;
		10109: rom = 1'b0;
		10110: rom = 1'b0;
		10111: rom = 1'b0;
		10112: rom = 1'b0;
		10113: rom = 1'b0;
		10114: rom = 1'b0;
		10115: rom = 1'b0;
		10116: rom = 1'b0;
		10117: rom = 1'b0;
		10118: rom = 1'b0;
		10119: rom = 1'b0;
		10120: rom = 1'b0;
		10121: rom = 1'b0;
		10122: rom = 1'b0;
		10123: rom = 1'b0;
		10124: rom = 1'b0;
		10125: rom = 1'b0;
		10126: rom = 1'b0;
		10127: rom = 1'b0;
		10128: rom = 1'b0;
		10129: rom = 1'b0;
		10130: rom = 1'b0;
		10131: rom = 1'b0;
		10132: rom = 1'b0;
		10133: rom = 1'b0;
		10134: rom = 1'b0;
		10135: rom = 1'b0;
		10136: rom = 1'b0;
		10137: rom = 1'b0;
		10138: rom = 1'b0;
		10139: rom = 1'b0;
		10140: rom = 1'b0;
		10141: rom = 1'b0;
		10142: rom = 1'b0;
		10143: rom = 1'b0;
		10144: rom = 1'b0;
		10145: rom = 1'b0;
		10146: rom = 1'b0;
		10147: rom = 1'b0;
		10148: rom = 1'b1;
		10149: rom = 1'b0;
		10150: rom = 1'b0;
		10151: rom = 1'b1;
		10152: rom = 1'b1;
		10153: rom = 1'b1;
		10154: rom = 1'b1;
		10155: rom = 1'b1;
		10156: rom = 1'b1;
		10157: rom = 1'b1;
		10158: rom = 1'b1;
		10159: rom = 1'b1;
		10160: rom = 1'b1;
		10161: rom = 1'b1;
		10162: rom = 1'b1;
		10163: rom = 1'b0;
		10164: rom = 1'b1;
		10165: rom = 1'b1;
		10166: rom = 1'b1;
		10167: rom = 1'b1;
		10168: rom = 1'b1;
		10169: rom = 1'b1;
		10170: rom = 1'b1;
		10171: rom = 1'b1;
		10172: rom = 1'b1;
		10173: rom = 1'b1;
		10174: rom = 1'b1;
		10175: rom = 1'b1;
		10176: rom = 1'b1;
		10177: rom = 1'b1;
		10178: rom = 1'b1;
		10179: rom = 1'b1;
		10180: rom = 1'b1;
		10181: rom = 1'b1;
		10182: rom = 1'b1;
		10183: rom = 1'b1;
		10184: rom = 1'b1;
		10185: rom = 1'b1;
		10186: rom = 1'b1;
		10187: rom = 1'b1;
		10188: rom = 1'b1;
		10189: rom = 1'b1;
		10190: rom = 1'b1;
		10191: rom = 1'b1;
		10192: rom = 1'b1;
		10193: rom = 1'b1;
		10194: rom = 1'b1;
		10195: rom = 1'b1;
		10196: rom = 1'b1;
		10197: rom = 1'b1;
		10198: rom = 1'b1;
		10199: rom = 1'b0;
		10200: rom = 1'b1;
		10201: rom = 1'b1;
		10202: rom = 1'b1;
		10203: rom = 1'b1;
		10204: rom = 1'b1;
		10205: rom = 1'b1;
		10206: rom = 1'b1;
		10207: rom = 1'b1;
		10208: rom = 1'b1;
		10209: rom = 1'b1;
		10210: rom = 1'b1;
		10211: rom = 1'b1;
		10212: rom = 1'b1;
		10213: rom = 1'b1;
		10214: rom = 1'b1;
		10215: rom = 1'b1;
		10216: rom = 1'b1;
		10217: rom = 1'b1;
		10218: rom = 1'b1;
		10219: rom = 1'b1;
		10220: rom = 1'b1;
		10221: rom = 1'b1;
		10222: rom = 1'b1;
		10223: rom = 1'b1;
		10224: rom = 1'b1;
		10225: rom = 1'b1;
		10226: rom = 1'b0;
		10227: rom = 1'b0;
		10228: rom = 1'b0;
		10229: rom = 1'b0;
		10230: rom = 1'b0;
		10231: rom = 1'b0;
		10232: rom = 1'b0;
		10233: rom = 1'b0;
		10234: rom = 1'b0;
		10235: rom = 1'b0;
		10236: rom = 1'b0;
		10237: rom = 1'b0;
		10238: rom = 1'b0;
		10239: rom = 1'b0;
		10240: rom = 1'b0;
		10241: rom = 1'b0;
		10242: rom = 1'b0;
		10243: rom = 1'b0;
		10244: rom = 1'b0;
		10245: rom = 1'b0;
		10246: rom = 1'b0;
		10247: rom = 1'b0;
		10248: rom = 1'b0;
		10249: rom = 1'b0;
		10250: rom = 1'b0;
		10251: rom = 1'b0;
		10252: rom = 1'b0;
		10253: rom = 1'b0;
		10254: rom = 1'b0;
		10255: rom = 1'b0;
		10256: rom = 1'b0;
		10257: rom = 1'b0;
		10258: rom = 1'b0;
		10259: rom = 1'b0;
		10260: rom = 1'b0;
		10261: rom = 1'b0;
		10262: rom = 1'b0;
		10263: rom = 1'b0;
		10264: rom = 1'b0;
		10265: rom = 1'b0;
		10266: rom = 1'b0;
		10267: rom = 1'b0;
		10268: rom = 1'b0;
		10269: rom = 1'b0;
		10270: rom = 1'b0;
		10271: rom = 1'b0;
		10272: rom = 1'b0;
		10273: rom = 1'b0;
		10274: rom = 1'b0;
		10275: rom = 1'b1;
		10276: rom = 1'b1;
		10277: rom = 1'b0;
		10278: rom = 1'b0;
		10279: rom = 1'b0;
		10280: rom = 1'b1;
		10281: rom = 1'b1;
		10282: rom = 1'b1;
		10283: rom = 1'b1;
		10284: rom = 1'b1;
		10285: rom = 1'b1;
		10286: rom = 1'b1;
		10287: rom = 1'b1;
		10288: rom = 1'b1;
		10289: rom = 1'b1;
		10290: rom = 1'b1;
		10291: rom = 1'b0;
		10292: rom = 1'b1;
		10293: rom = 1'b1;
		10294: rom = 1'b1;
		10295: rom = 1'b1;
		10296: rom = 1'b1;
		10297: rom = 1'b1;
		10298: rom = 1'b1;
		10299: rom = 1'b1;
		10300: rom = 1'b1;
		10301: rom = 1'b1;
		10302: rom = 1'b1;
		10303: rom = 1'b1;
		10304: rom = 1'b1;
		10305: rom = 1'b1;
		10306: rom = 1'b1;
		10307: rom = 1'b1;
		10308: rom = 1'b1;
		10309: rom = 1'b1;
		10310: rom = 1'b1;
		10311: rom = 1'b1;
		10312: rom = 1'b1;
		10313: rom = 1'b1;
		10314: rom = 1'b1;
		10315: rom = 1'b1;
		10316: rom = 1'b1;
		10317: rom = 1'b1;
		10318: rom = 1'b1;
		10319: rom = 1'b1;
		10320: rom = 1'b1;
		10321: rom = 1'b1;
		10322: rom = 1'b1;
		10323: rom = 1'b1;
		10324: rom = 1'b1;
		10325: rom = 1'b1;
		10326: rom = 1'b0;
		10327: rom = 1'b1;
		10328: rom = 1'b1;
		10329: rom = 1'b1;
		10330: rom = 1'b1;
		10331: rom = 1'b1;
		10332: rom = 1'b1;
		10333: rom = 1'b1;
		10334: rom = 1'b1;
		10335: rom = 1'b1;
		10336: rom = 1'b1;
		10337: rom = 1'b1;
		10338: rom = 1'b1;
		10339: rom = 1'b1;
		10340: rom = 1'b1;
		10341: rom = 1'b1;
		10342: rom = 1'b1;
		10343: rom = 1'b1;
		10344: rom = 1'b1;
		10345: rom = 1'b1;
		10346: rom = 1'b1;
		10347: rom = 1'b1;
		10348: rom = 1'b1;
		10349: rom = 1'b1;
		10350: rom = 1'b1;
		10351: rom = 1'b1;
		10352: rom = 1'b1;
		10353: rom = 1'b1;
		10354: rom = 1'b0;
		10355: rom = 1'b0;
		10356: rom = 1'b0;
		10357: rom = 1'b0;
		10358: rom = 1'b0;
		10359: rom = 1'b0;
		10360: rom = 1'b0;
		10361: rom = 1'b0;
		10362: rom = 1'b0;
		10363: rom = 1'b0;
		10364: rom = 1'b0;
		10365: rom = 1'b0;
		10366: rom = 1'b0;
		10367: rom = 1'b0;
		10368: rom = 1'b0;
		10369: rom = 1'b0;
		10370: rom = 1'b0;
		10371: rom = 1'b0;
		10372: rom = 1'b0;
		10373: rom = 1'b0;
		10374: rom = 1'b0;
		10375: rom = 1'b0;
		10376: rom = 1'b0;
		10377: rom = 1'b0;
		10378: rom = 1'b0;
		10379: rom = 1'b0;
		10380: rom = 1'b0;
		10381: rom = 1'b0;
		10382: rom = 1'b0;
		10383: rom = 1'b0;
		10384: rom = 1'b0;
		10385: rom = 1'b0;
		10386: rom = 1'b0;
		10387: rom = 1'b0;
		10388: rom = 1'b0;
		10389: rom = 1'b0;
		10390: rom = 1'b0;
		10391: rom = 1'b0;
		10392: rom = 1'b0;
		10393: rom = 1'b0;
		10394: rom = 1'b0;
		10395: rom = 1'b0;
		10396: rom = 1'b0;
		10397: rom = 1'b0;
		10398: rom = 1'b0;
		10399: rom = 1'b0;
		10400: rom = 1'b0;
		10401: rom = 1'b1;
		10402: rom = 1'b1;
		10403: rom = 1'b1;
		10404: rom = 1'b1;
		10405: rom = 1'b1;
		10406: rom = 1'b1;
		10407: rom = 1'b0;
		10408: rom = 1'b0;
		10409: rom = 1'b1;
		10410: rom = 1'b1;
		10411: rom = 1'b1;
		10412: rom = 1'b1;
		10413: rom = 1'b1;
		10414: rom = 1'b1;
		10415: rom = 1'b1;
		10416: rom = 1'b1;
		10417: rom = 1'b1;
		10418: rom = 1'b1;
		10419: rom = 1'b0;
		10420: rom = 1'b1;
		10421: rom = 1'b1;
		10422: rom = 1'b1;
		10423: rom = 1'b1;
		10424: rom = 1'b1;
		10425: rom = 1'b1;
		10426: rom = 1'b1;
		10427: rom = 1'b1;
		10428: rom = 1'b1;
		10429: rom = 1'b1;
		10430: rom = 1'b1;
		10431: rom = 1'b1;
		10432: rom = 1'b1;
		10433: rom = 1'b1;
		10434: rom = 1'b1;
		10435: rom = 1'b1;
		10436: rom = 1'b1;
		10437: rom = 1'b1;
		10438: rom = 1'b1;
		10439: rom = 1'b1;
		10440: rom = 1'b1;
		10441: rom = 1'b1;
		10442: rom = 1'b1;
		10443: rom = 1'b1;
		10444: rom = 1'b1;
		10445: rom = 1'b1;
		10446: rom = 1'b1;
		10447: rom = 1'b1;
		10448: rom = 1'b1;
		10449: rom = 1'b1;
		10450: rom = 1'b1;
		10451: rom = 1'b1;
		10452: rom = 1'b1;
		10453: rom = 1'b0;
		10454: rom = 1'b0;
		10455: rom = 1'b1;
		10456: rom = 1'b1;
		10457: rom = 1'b1;
		10458: rom = 1'b1;
		10459: rom = 1'b1;
		10460: rom = 1'b1;
		10461: rom = 1'b1;
		10462: rom = 1'b1;
		10463: rom = 1'b1;
		10464: rom = 1'b1;
		10465: rom = 1'b1;
		10466: rom = 1'b1;
		10467: rom = 1'b1;
		10468: rom = 1'b1;
		10469: rom = 1'b1;
		10470: rom = 1'b1;
		10471: rom = 1'b1;
		10472: rom = 1'b1;
		10473: rom = 1'b1;
		10474: rom = 1'b1;
		10475: rom = 1'b1;
		10476: rom = 1'b1;
		10477: rom = 1'b1;
		10478: rom = 1'b1;
		10479: rom = 1'b1;
		10480: rom = 1'b1;
		10481: rom = 1'b1;
		10482: rom = 1'b0;
		10483: rom = 1'b0;
		10484: rom = 1'b0;
		10485: rom = 1'b0;
		10486: rom = 1'b0;
		10487: rom = 1'b0;
		10488: rom = 1'b0;
		10489: rom = 1'b0;
		10490: rom = 1'b0;
		10491: rom = 1'b0;
		10492: rom = 1'b0;
		10493: rom = 1'b0;
		10494: rom = 1'b0;
		10495: rom = 1'b0;
		10496: rom = 1'b0;
		10497: rom = 1'b0;
		10498: rom = 1'b0;
		10499: rom = 1'b0;
		10500: rom = 1'b0;
		10501: rom = 1'b0;
		10502: rom = 1'b0;
		10503: rom = 1'b0;
		10504: rom = 1'b0;
		10505: rom = 1'b0;
		10506: rom = 1'b0;
		10507: rom = 1'b0;
		10508: rom = 1'b0;
		10509: rom = 1'b0;
		10510: rom = 1'b0;
		10511: rom = 1'b0;
		10512: rom = 1'b0;
		10513: rom = 1'b0;
		10514: rom = 1'b0;
		10515: rom = 1'b0;
		10516: rom = 1'b0;
		10517: rom = 1'b0;
		10518: rom = 1'b0;
		10519: rom = 1'b0;
		10520: rom = 1'b0;
		10521: rom = 1'b0;
		10522: rom = 1'b0;
		10523: rom = 1'b0;
		10524: rom = 1'b0;
		10525: rom = 1'b0;
		10526: rom = 1'b0;
		10527: rom = 1'b0;
		10528: rom = 1'b1;
		10529: rom = 1'b1;
		10530: rom = 1'b1;
		10531: rom = 1'b1;
		10532: rom = 1'b1;
		10533: rom = 1'b1;
		10534: rom = 1'b1;
		10535: rom = 1'b1;
		10536: rom = 1'b0;
		10537: rom = 1'b0;
		10538: rom = 1'b1;
		10539: rom = 1'b1;
		10540: rom = 1'b1;
		10541: rom = 1'b1;
		10542: rom = 1'b1;
		10543: rom = 1'b1;
		10544: rom = 1'b1;
		10545: rom = 1'b1;
		10546: rom = 1'b1;
		10547: rom = 1'b0;
		10548: rom = 1'b1;
		10549: rom = 1'b1;
		10550: rom = 1'b1;
		10551: rom = 1'b1;
		10552: rom = 1'b1;
		10553: rom = 1'b1;
		10554: rom = 1'b1;
		10555: rom = 1'b1;
		10556: rom = 1'b1;
		10557: rom = 1'b1;
		10558: rom = 1'b1;
		10559: rom = 1'b1;
		10560: rom = 1'b1;
		10561: rom = 1'b1;
		10562: rom = 1'b1;
		10563: rom = 1'b1;
		10564: rom = 1'b1;
		10565: rom = 1'b1;
		10566: rom = 1'b1;
		10567: rom = 1'b1;
		10568: rom = 1'b1;
		10569: rom = 1'b1;
		10570: rom = 1'b1;
		10571: rom = 1'b1;
		10572: rom = 1'b1;
		10573: rom = 1'b1;
		10574: rom = 1'b1;
		10575: rom = 1'b1;
		10576: rom = 1'b1;
		10577: rom = 1'b1;
		10578: rom = 1'b1;
		10579: rom = 1'b1;
		10580: rom = 1'b1;
		10581: rom = 1'b0;
		10582: rom = 1'b1;
		10583: rom = 1'b1;
		10584: rom = 1'b1;
		10585: rom = 1'b1;
		10586: rom = 1'b1;
		10587: rom = 1'b1;
		10588: rom = 1'b1;
		10589: rom = 1'b1;
		10590: rom = 1'b1;
		10591: rom = 1'b1;
		10592: rom = 1'b1;
		10593: rom = 1'b1;
		10594: rom = 1'b1;
		10595: rom = 1'b1;
		10596: rom = 1'b1;
		10597: rom = 1'b1;
		10598: rom = 1'b1;
		10599: rom = 1'b1;
		10600: rom = 1'b1;
		10601: rom = 1'b1;
		10602: rom = 1'b1;
		10603: rom = 1'b1;
		10604: rom = 1'b1;
		10605: rom = 1'b1;
		10606: rom = 1'b1;
		10607: rom = 1'b1;
		10608: rom = 1'b1;
		10609: rom = 1'b0;
		10610: rom = 1'b0;
		10611: rom = 1'b0;
		10612: rom = 1'b0;
		10613: rom = 1'b0;
		10614: rom = 1'b0;
		10615: rom = 1'b0;
		10616: rom = 1'b0;
		10617: rom = 1'b0;
		10618: rom = 1'b0;
		10619: rom = 1'b0;
		10620: rom = 1'b0;
		10621: rom = 1'b0;
		10622: rom = 1'b0;
		10623: rom = 1'b0;
		10624: rom = 1'b0;
		10625: rom = 1'b0;
		10626: rom = 1'b0;
		10627: rom = 1'b0;
		10628: rom = 1'b0;
		10629: rom = 1'b0;
		10630: rom = 1'b0;
		10631: rom = 1'b0;
		10632: rom = 1'b0;
		10633: rom = 1'b0;
		10634: rom = 1'b0;
		10635: rom = 1'b0;
		10636: rom = 1'b0;
		10637: rom = 1'b0;
		10638: rom = 1'b0;
		10639: rom = 1'b0;
		10640: rom = 1'b0;
		10641: rom = 1'b0;
		10642: rom = 1'b0;
		10643: rom = 1'b0;
		10644: rom = 1'b0;
		10645: rom = 1'b0;
		10646: rom = 1'b0;
		10647: rom = 1'b0;
		10648: rom = 1'b0;
		10649: rom = 1'b0;
		10650: rom = 1'b0;
		10651: rom = 1'b0;
		10652: rom = 1'b0;
		10653: rom = 1'b0;
		10654: rom = 1'b0;
		10655: rom = 1'b1;
		10656: rom = 1'b1;
		10657: rom = 1'b1;
		10658: rom = 1'b1;
		10659: rom = 1'b1;
		10660: rom = 1'b1;
		10661: rom = 1'b1;
		10662: rom = 1'b1;
		10663: rom = 1'b1;
		10664: rom = 1'b0;
		10665: rom = 1'b0;
		10666: rom = 1'b1;
		10667: rom = 1'b1;
		10668: rom = 1'b1;
		10669: rom = 1'b1;
		10670: rom = 1'b1;
		10671: rom = 1'b1;
		10672: rom = 1'b1;
		10673: rom = 1'b1;
		10674: rom = 1'b1;
		10675: rom = 1'b0;
		10676: rom = 1'b1;
		10677: rom = 1'b1;
		10678: rom = 1'b1;
		10679: rom = 1'b1;
		10680: rom = 1'b1;
		10681: rom = 1'b1;
		10682: rom = 1'b1;
		10683: rom = 1'b1;
		10684: rom = 1'b1;
		10685: rom = 1'b1;
		10686: rom = 1'b1;
		10687: rom = 1'b1;
		10688: rom = 1'b1;
		10689: rom = 1'b1;
		10690: rom = 1'b1;
		10691: rom = 1'b1;
		10692: rom = 1'b1;
		10693: rom = 1'b1;
		10694: rom = 1'b1;
		10695: rom = 1'b1;
		10696: rom = 1'b1;
		10697: rom = 1'b1;
		10698: rom = 1'b1;
		10699: rom = 1'b1;
		10700: rom = 1'b1;
		10701: rom = 1'b1;
		10702: rom = 1'b1;
		10703: rom = 1'b1;
		10704: rom = 1'b1;
		10705: rom = 1'b1;
		10706: rom = 1'b1;
		10707: rom = 1'b1;
		10708: rom = 1'b1;
		10709: rom = 1'b0;
		10710: rom = 1'b1;
		10711: rom = 1'b1;
		10712: rom = 1'b1;
		10713: rom = 1'b1;
		10714: rom = 1'b1;
		10715: rom = 1'b1;
		10716: rom = 1'b1;
		10717: rom = 1'b1;
		10718: rom = 1'b1;
		10719: rom = 1'b1;
		10720: rom = 1'b1;
		10721: rom = 1'b1;
		10722: rom = 1'b1;
		10723: rom = 1'b1;
		10724: rom = 1'b1;
		10725: rom = 1'b1;
		10726: rom = 1'b1;
		10727: rom = 1'b1;
		10728: rom = 1'b1;
		10729: rom = 1'b1;
		10730: rom = 1'b1;
		10731: rom = 1'b1;
		10732: rom = 1'b1;
		10733: rom = 1'b1;
		10734: rom = 1'b1;
		10735: rom = 1'b1;
		10736: rom = 1'b1;
		10737: rom = 1'b0;
		10738: rom = 1'b0;
		10739: rom = 1'b0;
		10740: rom = 1'b0;
		10741: rom = 1'b0;
		10742: rom = 1'b0;
		10743: rom = 1'b0;
		10744: rom = 1'b0;
		10745: rom = 1'b0;
		10746: rom = 1'b0;
		10747: rom = 1'b0;
		10748: rom = 1'b0;
		10749: rom = 1'b0;
		10750: rom = 1'b0;
		10751: rom = 1'b0;
		10752: rom = 1'b0;
		10753: rom = 1'b0;
		10754: rom = 1'b0;
		10755: rom = 1'b0;
		10756: rom = 1'b0;
		10757: rom = 1'b0;
		10758: rom = 1'b0;
		10759: rom = 1'b0;
		10760: rom = 1'b0;
		10761: rom = 1'b0;
		10762: rom = 1'b0;
		10763: rom = 1'b0;
		10764: rom = 1'b0;
		10765: rom = 1'b0;
		10766: rom = 1'b0;
		10767: rom = 1'b0;
		10768: rom = 1'b0;
		10769: rom = 1'b0;
		10770: rom = 1'b0;
		10771: rom = 1'b0;
		10772: rom = 1'b0;
		10773: rom = 1'b0;
		10774: rom = 1'b0;
		10775: rom = 1'b0;
		10776: rom = 1'b0;
		10777: rom = 1'b0;
		10778: rom = 1'b0;
		10779: rom = 1'b0;
		10780: rom = 1'b0;
		10781: rom = 1'b0;
		10782: rom = 1'b1;
		10783: rom = 1'b1;
		10784: rom = 1'b1;
		10785: rom = 1'b1;
		10786: rom = 1'b1;
		10787: rom = 1'b1;
		10788: rom = 1'b1;
		10789: rom = 1'b1;
		10790: rom = 1'b1;
		10791: rom = 1'b1;
		10792: rom = 1'b1;
		10793: rom = 1'b1;
		10794: rom = 1'b0;
		10795: rom = 1'b0;
		10796: rom = 1'b1;
		10797: rom = 1'b1;
		10798: rom = 1'b1;
		10799: rom = 1'b1;
		10800: rom = 1'b1;
		10801: rom = 1'b1;
		10802: rom = 1'b1;
		10803: rom = 1'b1;
		10804: rom = 1'b0;
		10805: rom = 1'b1;
		10806: rom = 1'b1;
		10807: rom = 1'b1;
		10808: rom = 1'b1;
		10809: rom = 1'b1;
		10810: rom = 1'b1;
		10811: rom = 1'b1;
		10812: rom = 1'b1;
		10813: rom = 1'b1;
		10814: rom = 1'b1;
		10815: rom = 1'b1;
		10816: rom = 1'b1;
		10817: rom = 1'b1;
		10818: rom = 1'b1;
		10819: rom = 1'b1;
		10820: rom = 1'b1;
		10821: rom = 1'b1;
		10822: rom = 1'b1;
		10823: rom = 1'b1;
		10824: rom = 1'b1;
		10825: rom = 1'b1;
		10826: rom = 1'b1;
		10827: rom = 1'b1;
		10828: rom = 1'b1;
		10829: rom = 1'b1;
		10830: rom = 1'b1;
		10831: rom = 1'b1;
		10832: rom = 1'b1;
		10833: rom = 1'b1;
		10834: rom = 1'b1;
		10835: rom = 1'b1;
		10836: rom = 1'b0;
		10837: rom = 1'b1;
		10838: rom = 1'b1;
		10839: rom = 1'b1;
		10840: rom = 1'b1;
		10841: rom = 1'b1;
		10842: rom = 1'b1;
		10843: rom = 1'b1;
		10844: rom = 1'b1;
		10845: rom = 1'b1;
		10846: rom = 1'b1;
		10847: rom = 1'b1;
		10848: rom = 1'b1;
		10849: rom = 1'b1;
		10850: rom = 1'b1;
		10851: rom = 1'b1;
		10852: rom = 1'b1;
		10853: rom = 1'b1;
		10854: rom = 1'b1;
		10855: rom = 1'b1;
		10856: rom = 1'b1;
		10857: rom = 1'b1;
		10858: rom = 1'b1;
		10859: rom = 1'b1;
		10860: rom = 1'b1;
		10861: rom = 1'b1;
		10862: rom = 1'b1;
		10863: rom = 1'b1;
		10864: rom = 1'b0;
		10865: rom = 1'b0;
		10866: rom = 1'b0;
		10867: rom = 1'b0;
		10868: rom = 1'b0;
		10869: rom = 1'b0;
		10870: rom = 1'b0;
		10871: rom = 1'b0;
		10872: rom = 1'b0;
		10873: rom = 1'b0;
		10874: rom = 1'b0;
		10875: rom = 1'b0;
		10876: rom = 1'b0;
		10877: rom = 1'b0;
		10878: rom = 1'b0;
		10879: rom = 1'b0;
		10880: rom = 1'b0;
		10881: rom = 1'b0;
		10882: rom = 1'b0;
		10883: rom = 1'b0;
		10884: rom = 1'b0;
		10885: rom = 1'b0;
		10886: rom = 1'b0;
		10887: rom = 1'b0;
		10888: rom = 1'b0;
		10889: rom = 1'b0;
		10890: rom = 1'b0;
		10891: rom = 1'b0;
		10892: rom = 1'b0;
		10893: rom = 1'b0;
		10894: rom = 1'b0;
		10895: rom = 1'b0;
		10896: rom = 1'b0;
		10897: rom = 1'b0;
		10898: rom = 1'b0;
		10899: rom = 1'b0;
		10900: rom = 1'b0;
		10901: rom = 1'b0;
		10902: rom = 1'b0;
		10903: rom = 1'b0;
		10904: rom = 1'b0;
		10905: rom = 1'b0;
		10906: rom = 1'b0;
		10907: rom = 1'b0;
		10908: rom = 1'b0;
		10909: rom = 1'b1;
		10910: rom = 1'b1;
		10911: rom = 1'b1;
		10912: rom = 1'b1;
		10913: rom = 1'b1;
		10914: rom = 1'b1;
		10915: rom = 1'b1;
		10916: rom = 1'b1;
		10917: rom = 1'b1;
		10918: rom = 1'b1;
		10919: rom = 1'b1;
		10920: rom = 1'b1;
		10921: rom = 1'b1;
		10922: rom = 1'b1;
		10923: rom = 1'b0;
		10924: rom = 1'b0;
		10925: rom = 1'b1;
		10926: rom = 1'b1;
		10927: rom = 1'b1;
		10928: rom = 1'b1;
		10929: rom = 1'b1;
		10930: rom = 1'b1;
		10931: rom = 1'b1;
		10932: rom = 1'b0;
		10933: rom = 1'b1;
		10934: rom = 1'b1;
		10935: rom = 1'b1;
		10936: rom = 1'b1;
		10937: rom = 1'b1;
		10938: rom = 1'b1;
		10939: rom = 1'b1;
		10940: rom = 1'b1;
		10941: rom = 1'b1;
		10942: rom = 1'b1;
		10943: rom = 1'b1;
		10944: rom = 1'b1;
		10945: rom = 1'b1;
		10946: rom = 1'b1;
		10947: rom = 1'b1;
		10948: rom = 1'b1;
		10949: rom = 1'b1;
		10950: rom = 1'b1;
		10951: rom = 1'b1;
		10952: rom = 1'b1;
		10953: rom = 1'b1;
		10954: rom = 1'b1;
		10955: rom = 1'b1;
		10956: rom = 1'b1;
		10957: rom = 1'b1;
		10958: rom = 1'b1;
		10959: rom = 1'b1;
		10960: rom = 1'b1;
		10961: rom = 1'b1;
		10962: rom = 1'b1;
		10963: rom = 1'b1;
		10964: rom = 1'b0;
		10965: rom = 1'b1;
		10966: rom = 1'b1;
		10967: rom = 1'b1;
		10968: rom = 1'b1;
		10969: rom = 1'b1;
		10970: rom = 1'b1;
		10971: rom = 1'b1;
		10972: rom = 1'b1;
		10973: rom = 1'b1;
		10974: rom = 1'b1;
		10975: rom = 1'b1;
		10976: rom = 1'b1;
		10977: rom = 1'b1;
		10978: rom = 1'b1;
		10979: rom = 1'b1;
		10980: rom = 1'b1;
		10981: rom = 1'b1;
		10982: rom = 1'b1;
		10983: rom = 1'b1;
		10984: rom = 1'b1;
		10985: rom = 1'b1;
		10986: rom = 1'b1;
		10987: rom = 1'b1;
		10988: rom = 1'b1;
		10989: rom = 1'b1;
		10990: rom = 1'b1;
		10991: rom = 1'b1;
		10992: rom = 1'b0;
		10993: rom = 1'b0;
		10994: rom = 1'b0;
		10995: rom = 1'b0;
		10996: rom = 1'b0;
		10997: rom = 1'b0;
		10998: rom = 1'b0;
		10999: rom = 1'b0;
		11000: rom = 1'b0;
		11001: rom = 1'b0;
		11002: rom = 1'b0;
		11003: rom = 1'b0;
		11004: rom = 1'b0;
		11005: rom = 1'b0;
		11006: rom = 1'b0;
		11007: rom = 1'b0;
		11008: rom = 1'b0;
		11009: rom = 1'b0;
		11010: rom = 1'b0;
		11011: rom = 1'b0;
		11012: rom = 1'b0;
		11013: rom = 1'b0;
		11014: rom = 1'b0;
		11015: rom = 1'b0;
		11016: rom = 1'b0;
		11017: rom = 1'b0;
		11018: rom = 1'b0;
		11019: rom = 1'b0;
		11020: rom = 1'b0;
		11021: rom = 1'b0;
		11022: rom = 1'b0;
		11023: rom = 1'b0;
		11024: rom = 1'b0;
		11025: rom = 1'b0;
		11026: rom = 1'b0;
		11027: rom = 1'b0;
		11028: rom = 1'b0;
		11029: rom = 1'b0;
		11030: rom = 1'b0;
		11031: rom = 1'b0;
		11032: rom = 1'b0;
		11033: rom = 1'b0;
		11034: rom = 1'b0;
		11035: rom = 1'b0;
		11036: rom = 1'b1;
		11037: rom = 1'b1;
		11038: rom = 1'b1;
		11039: rom = 1'b1;
		11040: rom = 1'b1;
		11041: rom = 1'b1;
		11042: rom = 1'b1;
		11043: rom = 1'b1;
		11044: rom = 1'b1;
		11045: rom = 1'b1;
		11046: rom = 1'b1;
		11047: rom = 1'b1;
		11048: rom = 1'b1;
		11049: rom = 1'b1;
		11050: rom = 1'b1;
		11051: rom = 1'b1;
		11052: rom = 1'b0;
		11053: rom = 1'b0;
		11054: rom = 1'b1;
		11055: rom = 1'b1;
		11056: rom = 1'b1;
		11057: rom = 1'b1;
		11058: rom = 1'b1;
		11059: rom = 1'b1;
		11060: rom = 1'b0;
		11061: rom = 1'b1;
		11062: rom = 1'b1;
		11063: rom = 1'b1;
		11064: rom = 1'b1;
		11065: rom = 1'b1;
		11066: rom = 1'b1;
		11067: rom = 1'b1;
		11068: rom = 1'b1;
		11069: rom = 1'b1;
		11070: rom = 1'b1;
		11071: rom = 1'b1;
		11072: rom = 1'b1;
		11073: rom = 1'b1;
		11074: rom = 1'b1;
		11075: rom = 1'b1;
		11076: rom = 1'b1;
		11077: rom = 1'b1;
		11078: rom = 1'b1;
		11079: rom = 1'b1;
		11080: rom = 1'b1;
		11081: rom = 1'b1;
		11082: rom = 1'b1;
		11083: rom = 1'b1;
		11084: rom = 1'b1;
		11085: rom = 1'b1;
		11086: rom = 1'b1;
		11087: rom = 1'b1;
		11088: rom = 1'b1;
		11089: rom = 1'b1;
		11090: rom = 1'b1;
		11091: rom = 1'b0;
		11092: rom = 1'b0;
		11093: rom = 1'b1;
		11094: rom = 1'b1;
		11095: rom = 1'b1;
		11096: rom = 1'b1;
		11097: rom = 1'b1;
		11098: rom = 1'b1;
		11099: rom = 1'b1;
		11100: rom = 1'b1;
		11101: rom = 1'b1;
		11102: rom = 1'b1;
		11103: rom = 1'b1;
		11104: rom = 1'b1;
		11105: rom = 1'b1;
		11106: rom = 1'b1;
		11107: rom = 1'b1;
		11108: rom = 1'b1;
		11109: rom = 1'b1;
		11110: rom = 1'b1;
		11111: rom = 1'b1;
		11112: rom = 1'b1;
		11113: rom = 1'b1;
		11114: rom = 1'b1;
		11115: rom = 1'b1;
		11116: rom = 1'b1;
		11117: rom = 1'b1;
		11118: rom = 1'b1;
		11119: rom = 1'b0;
		11120: rom = 1'b0;
		11121: rom = 1'b0;
		11122: rom = 1'b0;
		11123: rom = 1'b0;
		11124: rom = 1'b0;
		11125: rom = 1'b0;
		11126: rom = 1'b0;
		11127: rom = 1'b0;
		11128: rom = 1'b0;
		11129: rom = 1'b0;
		11130: rom = 1'b0;
		11131: rom = 1'b0;
		11132: rom = 1'b0;
		11133: rom = 1'b0;
		11134: rom = 1'b0;
		11135: rom = 1'b0;
		11136: rom = 1'b0;
		11137: rom = 1'b0;
		11138: rom = 1'b0;
		11139: rom = 1'b0;
		11140: rom = 1'b0;
		11141: rom = 1'b0;
		11142: rom = 1'b0;
		11143: rom = 1'b0;
		11144: rom = 1'b0;
		11145: rom = 1'b0;
		11146: rom = 1'b0;
		11147: rom = 1'b0;
		11148: rom = 1'b0;
		11149: rom = 1'b0;
		11150: rom = 1'b0;
		11151: rom = 1'b0;
		11152: rom = 1'b0;
		11153: rom = 1'b0;
		11154: rom = 1'b0;
		11155: rom = 1'b0;
		11156: rom = 1'b0;
		11157: rom = 1'b0;
		11158: rom = 1'b0;
		11159: rom = 1'b0;
		11160: rom = 1'b0;
		11161: rom = 1'b0;
		11162: rom = 1'b0;
		11163: rom = 1'b1;
		11164: rom = 1'b1;
		11165: rom = 1'b1;
		11166: rom = 1'b1;
		11167: rom = 1'b1;
		11168: rom = 1'b1;
		11169: rom = 1'b1;
		11170: rom = 1'b1;
		11171: rom = 1'b1;
		11172: rom = 1'b1;
		11173: rom = 1'b1;
		11174: rom = 1'b1;
		11175: rom = 1'b1;
		11176: rom = 1'b1;
		11177: rom = 1'b1;
		11178: rom = 1'b1;
		11179: rom = 1'b1;
		11180: rom = 1'b1;
		11181: rom = 1'b1;
		11182: rom = 1'b0;
		11183: rom = 1'b0;
		11184: rom = 1'b1;
		11185: rom = 1'b1;
		11186: rom = 1'b1;
		11187: rom = 1'b1;
		11188: rom = 1'b0;
		11189: rom = 1'b0;
		11190: rom = 1'b1;
		11191: rom = 1'b1;
		11192: rom = 1'b1;
		11193: rom = 1'b1;
		11194: rom = 1'b1;
		11195: rom = 1'b1;
		11196: rom = 1'b1;
		11197: rom = 1'b1;
		11198: rom = 1'b1;
		11199: rom = 1'b1;
		11200: rom = 1'b1;
		11201: rom = 1'b1;
		11202: rom = 1'b1;
		11203: rom = 1'b1;
		11204: rom = 1'b1;
		11205: rom = 1'b1;
		11206: rom = 1'b1;
		11207: rom = 1'b1;
		11208: rom = 1'b1;
		11209: rom = 1'b1;
		11210: rom = 1'b1;
		11211: rom = 1'b1;
		11212: rom = 1'b1;
		11213: rom = 1'b1;
		11214: rom = 1'b1;
		11215: rom = 1'b1;
		11216: rom = 1'b1;
		11217: rom = 1'b1;
		11218: rom = 1'b1;
		11219: rom = 1'b0;
		11220: rom = 1'b1;
		11221: rom = 1'b1;
		11222: rom = 1'b1;
		11223: rom = 1'b1;
		11224: rom = 1'b1;
		11225: rom = 1'b1;
		11226: rom = 1'b1;
		11227: rom = 1'b1;
		11228: rom = 1'b1;
		11229: rom = 1'b1;
		11230: rom = 1'b1;
		11231: rom = 1'b1;
		11232: rom = 1'b1;
		11233: rom = 1'b1;
		11234: rom = 1'b1;
		11235: rom = 1'b1;
		11236: rom = 1'b1;
		11237: rom = 1'b1;
		11238: rom = 1'b1;
		11239: rom = 1'b1;
		11240: rom = 1'b1;
		11241: rom = 1'b1;
		11242: rom = 1'b1;
		11243: rom = 1'b1;
		11244: rom = 1'b1;
		11245: rom = 1'b1;
		11246: rom = 1'b1;
		11247: rom = 1'b0;
		11248: rom = 1'b0;
		11249: rom = 1'b0;
		11250: rom = 1'b0;
		11251: rom = 1'b0;
		11252: rom = 1'b0;
		11253: rom = 1'b0;
		11254: rom = 1'b0;
		11255: rom = 1'b0;
		11256: rom = 1'b0;
		11257: rom = 1'b0;
		11258: rom = 1'b0;
		11259: rom = 1'b0;
		11260: rom = 1'b0;
		11261: rom = 1'b0;
		11262: rom = 1'b0;
		11263: rom = 1'b0;
		11264: rom = 1'b0;
		11265: rom = 1'b0;
		11266: rom = 1'b0;
		11267: rom = 1'b0;
		11268: rom = 1'b0;
		11269: rom = 1'b0;
		11270: rom = 1'b0;
		11271: rom = 1'b0;
		11272: rom = 1'b0;
		11273: rom = 1'b0;
		11274: rom = 1'b0;
		11275: rom = 1'b0;
		11276: rom = 1'b0;
		11277: rom = 1'b0;
		11278: rom = 1'b0;
		11279: rom = 1'b0;
		11280: rom = 1'b0;
		11281: rom = 1'b0;
		11282: rom = 1'b0;
		11283: rom = 1'b0;
		11284: rom = 1'b0;
		11285: rom = 1'b0;
		11286: rom = 1'b0;
		11287: rom = 1'b0;
		11288: rom = 1'b0;
		11289: rom = 1'b0;
		11290: rom = 1'b1;
		11291: rom = 1'b1;
		11292: rom = 1'b1;
		11293: rom = 1'b1;
		11294: rom = 1'b1;
		11295: rom = 1'b1;
		11296: rom = 1'b1;
		11297: rom = 1'b1;
		11298: rom = 1'b1;
		11299: rom = 1'b1;
		11300: rom = 1'b1;
		11301: rom = 1'b1;
		11302: rom = 1'b1;
		11303: rom = 1'b1;
		11304: rom = 1'b1;
		11305: rom = 1'b1;
		11306: rom = 1'b1;
		11307: rom = 1'b1;
		11308: rom = 1'b1;
		11309: rom = 1'b1;
		11310: rom = 1'b1;
		11311: rom = 1'b0;
		11312: rom = 1'b0;
		11313: rom = 1'b1;
		11314: rom = 1'b1;
		11315: rom = 1'b1;
		11316: rom = 1'b1;
		11317: rom = 1'b0;
		11318: rom = 1'b1;
		11319: rom = 1'b1;
		11320: rom = 1'b1;
		11321: rom = 1'b1;
		11322: rom = 1'b1;
		11323: rom = 1'b1;
		11324: rom = 1'b1;
		11325: rom = 1'b1;
		11326: rom = 1'b1;
		11327: rom = 1'b1;
		11328: rom = 1'b1;
		11329: rom = 1'b1;
		11330: rom = 1'b1;
		11331: rom = 1'b1;
		11332: rom = 1'b1;
		11333: rom = 1'b1;
		11334: rom = 1'b1;
		11335: rom = 1'b1;
		11336: rom = 1'b1;
		11337: rom = 1'b1;
		11338: rom = 1'b1;
		11339: rom = 1'b1;
		11340: rom = 1'b1;
		11341: rom = 1'b1;
		11342: rom = 1'b1;
		11343: rom = 1'b1;
		11344: rom = 1'b1;
		11345: rom = 1'b1;
		11346: rom = 1'b0;
		11347: rom = 1'b0;
		11348: rom = 1'b1;
		11349: rom = 1'b1;
		11350: rom = 1'b1;
		11351: rom = 1'b1;
		11352: rom = 1'b1;
		11353: rom = 1'b1;
		11354: rom = 1'b1;
		11355: rom = 1'b1;
		11356: rom = 1'b1;
		11357: rom = 1'b1;
		11358: rom = 1'b1;
		11359: rom = 1'b1;
		11360: rom = 1'b1;
		11361: rom = 1'b1;
		11362: rom = 1'b1;
		11363: rom = 1'b1;
		11364: rom = 1'b1;
		11365: rom = 1'b1;
		11366: rom = 1'b1;
		11367: rom = 1'b1;
		11368: rom = 1'b1;
		11369: rom = 1'b1;
		11370: rom = 1'b1;
		11371: rom = 1'b1;
		11372: rom = 1'b1;
		11373: rom = 1'b1;
		11374: rom = 1'b1;
		11375: rom = 1'b0;
		11376: rom = 1'b0;
		11377: rom = 1'b0;
		11378: rom = 1'b0;
		11379: rom = 1'b0;
		11380: rom = 1'b0;
		11381: rom = 1'b0;
		11382: rom = 1'b0;
		11383: rom = 1'b0;
		11384: rom = 1'b0;
		11385: rom = 1'b0;
		11386: rom = 1'b0;
		11387: rom = 1'b0;
		11388: rom = 1'b0;
		11389: rom = 1'b0;
		11390: rom = 1'b0;
		11391: rom = 1'b0;
		11392: rom = 1'b0;
		11393: rom = 1'b0;
		11394: rom = 1'b0;
		11395: rom = 1'b0;
		11396: rom = 1'b0;
		11397: rom = 1'b0;
		11398: rom = 1'b0;
		11399: rom = 1'b0;
		11400: rom = 1'b0;
		11401: rom = 1'b0;
		11402: rom = 1'b0;
		11403: rom = 1'b0;
		11404: rom = 1'b0;
		11405: rom = 1'b0;
		11406: rom = 1'b0;
		11407: rom = 1'b0;
		11408: rom = 1'b0;
		11409: rom = 1'b0;
		11410: rom = 1'b0;
		11411: rom = 1'b0;
		11412: rom = 1'b0;
		11413: rom = 1'b0;
		11414: rom = 1'b0;
		11415: rom = 1'b0;
		11416: rom = 1'b0;
		11417: rom = 1'b1;
		11418: rom = 1'b1;
		11419: rom = 1'b1;
		11420: rom = 1'b1;
		11421: rom = 1'b1;
		11422: rom = 1'b1;
		11423: rom = 1'b1;
		11424: rom = 1'b1;
		11425: rom = 1'b1;
		11426: rom = 1'b1;
		11427: rom = 1'b1;
		11428: rom = 1'b1;
		11429: rom = 1'b1;
		11430: rom = 1'b1;
		11431: rom = 1'b1;
		11432: rom = 1'b1;
		11433: rom = 1'b1;
		11434: rom = 1'b1;
		11435: rom = 1'b1;
		11436: rom = 1'b1;
		11437: rom = 1'b1;
		11438: rom = 1'b1;
		11439: rom = 1'b1;
		11440: rom = 1'b1;
		11441: rom = 1'b0;
		11442: rom = 1'b0;
		11443: rom = 1'b1;
		11444: rom = 1'b1;
		11445: rom = 1'b0;
		11446: rom = 1'b1;
		11447: rom = 1'b1;
		11448: rom = 1'b1;
		11449: rom = 1'b1;
		11450: rom = 1'b1;
		11451: rom = 1'b1;
		11452: rom = 1'b1;
		11453: rom = 1'b1;
		11454: rom = 1'b1;
		11455: rom = 1'b1;
		11456: rom = 1'b1;
		11457: rom = 1'b1;
		11458: rom = 1'b1;
		11459: rom = 1'b1;
		11460: rom = 1'b1;
		11461: rom = 1'b1;
		11462: rom = 1'b1;
		11463: rom = 1'b1;
		11464: rom = 1'b1;
		11465: rom = 1'b1;
		11466: rom = 1'b1;
		11467: rom = 1'b1;
		11468: rom = 1'b1;
		11469: rom = 1'b1;
		11470: rom = 1'b1;
		11471: rom = 1'b1;
		11472: rom = 1'b1;
		11473: rom = 1'b1;
		11474: rom = 1'b0;
		11475: rom = 1'b0;
		11476: rom = 1'b1;
		11477: rom = 1'b1;
		11478: rom = 1'b1;
		11479: rom = 1'b1;
		11480: rom = 1'b1;
		11481: rom = 1'b1;
		11482: rom = 1'b1;
		11483: rom = 1'b1;
		11484: rom = 1'b1;
		11485: rom = 1'b1;
		11486: rom = 1'b1;
		11487: rom = 1'b1;
		11488: rom = 1'b1;
		11489: rom = 1'b1;
		11490: rom = 1'b1;
		11491: rom = 1'b1;
		11492: rom = 1'b1;
		11493: rom = 1'b1;
		11494: rom = 1'b1;
		11495: rom = 1'b1;
		11496: rom = 1'b1;
		11497: rom = 1'b1;
		11498: rom = 1'b1;
		11499: rom = 1'b1;
		11500: rom = 1'b1;
		11501: rom = 1'b1;
		11502: rom = 1'b0;
		11503: rom = 1'b0;
		11504: rom = 1'b0;
		11505: rom = 1'b0;
		11506: rom = 1'b0;
		11507: rom = 1'b0;
		11508: rom = 1'b0;
		11509: rom = 1'b0;
		11510: rom = 1'b0;
		11511: rom = 1'b0;
		11512: rom = 1'b0;
		11513: rom = 1'b0;
		11514: rom = 1'b0;
		11515: rom = 1'b0;
		11516: rom = 1'b0;
		11517: rom = 1'b0;
		11518: rom = 1'b0;
		11519: rom = 1'b0;
		11520: rom = 1'b0;
		11521: rom = 1'b0;
		11522: rom = 1'b0;
		11523: rom = 1'b0;
		11524: rom = 1'b0;
		11525: rom = 1'b0;
		11526: rom = 1'b0;
		11527: rom = 1'b0;
		11528: rom = 1'b0;
		11529: rom = 1'b0;
		11530: rom = 1'b0;
		11531: rom = 1'b0;
		11532: rom = 1'b0;
		11533: rom = 1'b0;
		11534: rom = 1'b0;
		11535: rom = 1'b0;
		11536: rom = 1'b0;
		11537: rom = 1'b0;
		11538: rom = 1'b0;
		11539: rom = 1'b0;
		11540: rom = 1'b0;
		11541: rom = 1'b0;
		11542: rom = 1'b0;
		11543: rom = 1'b0;
		11544: rom = 1'b0;
		11545: rom = 1'b1;
		11546: rom = 1'b1;
		11547: rom = 1'b1;
		11548: rom = 1'b1;
		11549: rom = 1'b1;
		11550: rom = 1'b1;
		11551: rom = 1'b1;
		11552: rom = 1'b1;
		11553: rom = 1'b1;
		11554: rom = 1'b1;
		11555: rom = 1'b1;
		11556: rom = 1'b1;
		11557: rom = 1'b1;
		11558: rom = 1'b1;
		11559: rom = 1'b1;
		11560: rom = 1'b1;
		11561: rom = 1'b1;
		11562: rom = 1'b1;
		11563: rom = 1'b1;
		11564: rom = 1'b1;
		11565: rom = 1'b1;
		11566: rom = 1'b1;
		11567: rom = 1'b1;
		11568: rom = 1'b1;
		11569: rom = 1'b1;
		11570: rom = 1'b0;
		11571: rom = 1'b0;
		11572: rom = 1'b0;
		11573: rom = 1'b0;
		11574: rom = 1'b1;
		11575: rom = 1'b1;
		11576: rom = 1'b1;
		11577: rom = 1'b1;
		11578: rom = 1'b1;
		11579: rom = 1'b1;
		11580: rom = 1'b1;
		11581: rom = 1'b1;
		11582: rom = 1'b1;
		11583: rom = 1'b1;
		11584: rom = 1'b1;
		11585: rom = 1'b1;
		11586: rom = 1'b1;
		11587: rom = 1'b1;
		11588: rom = 1'b1;
		11589: rom = 1'b1;
		11590: rom = 1'b1;
		11591: rom = 1'b1;
		11592: rom = 1'b1;
		11593: rom = 1'b1;
		11594: rom = 1'b1;
		11595: rom = 1'b1;
		11596: rom = 1'b1;
		11597: rom = 1'b1;
		11598: rom = 1'b1;
		11599: rom = 1'b1;
		11600: rom = 1'b1;
		11601: rom = 1'b1;
		11602: rom = 1'b0;
		11603: rom = 1'b1;
		11604: rom = 1'b1;
		11605: rom = 1'b1;
		11606: rom = 1'b1;
		11607: rom = 1'b1;
		11608: rom = 1'b1;
		11609: rom = 1'b1;
		11610: rom = 1'b1;
		11611: rom = 1'b1;
		11612: rom = 1'b1;
		11613: rom = 1'b1;
		11614: rom = 1'b1;
		11615: rom = 1'b1;
		11616: rom = 1'b1;
		11617: rom = 1'b1;
		11618: rom = 1'b1;
		11619: rom = 1'b1;
		11620: rom = 1'b1;
		11621: rom = 1'b1;
		11622: rom = 1'b1;
		11623: rom = 1'b1;
		11624: rom = 1'b1;
		11625: rom = 1'b1;
		11626: rom = 1'b1;
		11627: rom = 1'b1;
		11628: rom = 1'b1;
		11629: rom = 1'b1;
		11630: rom = 1'b0;
		11631: rom = 1'b0;
		11632: rom = 1'b0;
		11633: rom = 1'b0;
		11634: rom = 1'b0;
		11635: rom = 1'b0;
		11636: rom = 1'b0;
		11637: rom = 1'b0;
		11638: rom = 1'b0;
		11639: rom = 1'b0;
		11640: rom = 1'b0;
		11641: rom = 1'b0;
		11642: rom = 1'b0;
		11643: rom = 1'b0;
		11644: rom = 1'b0;
		11645: rom = 1'b0;
		11646: rom = 1'b0;
		11647: rom = 1'b0;
		11648: rom = 1'b0;
		11649: rom = 1'b0;
		11650: rom = 1'b0;
		11651: rom = 1'b0;
		11652: rom = 1'b0;
		11653: rom = 1'b0;
		11654: rom = 1'b0;
		11655: rom = 1'b0;
		11656: rom = 1'b0;
		11657: rom = 1'b0;
		11658: rom = 1'b0;
		11659: rom = 1'b0;
		11660: rom = 1'b0;
		11661: rom = 1'b0;
		11662: rom = 1'b0;
		11663: rom = 1'b0;
		11664: rom = 1'b0;
		11665: rom = 1'b0;
		11666: rom = 1'b0;
		11667: rom = 1'b0;
		11668: rom = 1'b0;
		11669: rom = 1'b0;
		11670: rom = 1'b0;
		11671: rom = 1'b0;
		11672: rom = 1'b1;
		11673: rom = 1'b1;
		11674: rom = 1'b1;
		11675: rom = 1'b1;
		11676: rom = 1'b1;
		11677: rom = 1'b1;
		11678: rom = 1'b1;
		11679: rom = 1'b1;
		11680: rom = 1'b1;
		11681: rom = 1'b1;
		11682: rom = 1'b1;
		11683: rom = 1'b1;
		11684: rom = 1'b1;
		11685: rom = 1'b1;
		11686: rom = 1'b1;
		11687: rom = 1'b1;
		11688: rom = 1'b1;
		11689: rom = 1'b1;
		11690: rom = 1'b1;
		11691: rom = 1'b1;
		11692: rom = 1'b1;
		11693: rom = 1'b1;
		11694: rom = 1'b1;
		11695: rom = 1'b1;
		11696: rom = 1'b1;
		11697: rom = 1'b1;
		11698: rom = 1'b1;
		11699: rom = 1'b1;
		11700: rom = 1'b0;
		11701: rom = 1'b0;
		11702: rom = 1'b0;
		11703: rom = 1'b1;
		11704: rom = 1'b1;
		11705: rom = 1'b1;
		11706: rom = 1'b1;
		11707: rom = 1'b1;
		11708: rom = 1'b1;
		11709: rom = 1'b1;
		11710: rom = 1'b1;
		11711: rom = 1'b1;
		11712: rom = 1'b1;
		11713: rom = 1'b1;
		11714: rom = 1'b1;
		11715: rom = 1'b1;
		11716: rom = 1'b1;
		11717: rom = 1'b1;
		11718: rom = 1'b1;
		11719: rom = 1'b1;
		11720: rom = 1'b1;
		11721: rom = 1'b1;
		11722: rom = 1'b1;
		11723: rom = 1'b1;
		11724: rom = 1'b1;
		11725: rom = 1'b1;
		11726: rom = 1'b1;
		11727: rom = 1'b1;
		11728: rom = 1'b1;
		11729: rom = 1'b0;
		11730: rom = 1'b0;
		11731: rom = 1'b1;
		11732: rom = 1'b1;
		11733: rom = 1'b1;
		11734: rom = 1'b1;
		11735: rom = 1'b1;
		11736: rom = 1'b1;
		11737: rom = 1'b1;
		11738: rom = 1'b1;
		11739: rom = 1'b1;
		11740: rom = 1'b1;
		11741: rom = 1'b1;
		11742: rom = 1'b1;
		11743: rom = 1'b1;
		11744: rom = 1'b1;
		11745: rom = 1'b1;
		11746: rom = 1'b1;
		11747: rom = 1'b1;
		11748: rom = 1'b1;
		11749: rom = 1'b1;
		11750: rom = 1'b1;
		11751: rom = 1'b1;
		11752: rom = 1'b1;
		11753: rom = 1'b1;
		11754: rom = 1'b1;
		11755: rom = 1'b1;
		11756: rom = 1'b1;
		11757: rom = 1'b0;
		11758: rom = 1'b0;
		11759: rom = 1'b0;
		11760: rom = 1'b0;
		11761: rom = 1'b0;
		11762: rom = 1'b0;
		11763: rom = 1'b0;
		11764: rom = 1'b0;
		11765: rom = 1'b0;
		11766: rom = 1'b0;
		11767: rom = 1'b0;
		11768: rom = 1'b0;
		11769: rom = 1'b0;
		11770: rom = 1'b0;
		11771: rom = 1'b0;
		11772: rom = 1'b0;
		11773: rom = 1'b0;
		11774: rom = 1'b0;
		11775: rom = 1'b0;
		11776: rom = 1'b0;
		11777: rom = 1'b0;
		11778: rom = 1'b0;
		11779: rom = 1'b0;
		11780: rom = 1'b0;
		11781: rom = 1'b0;
		11782: rom = 1'b0;
		11783: rom = 1'b0;
		11784: rom = 1'b0;
		11785: rom = 1'b0;
		11786: rom = 1'b0;
		11787: rom = 1'b0;
		11788: rom = 1'b0;
		11789: rom = 1'b0;
		11790: rom = 1'b0;
		11791: rom = 1'b0;
		11792: rom = 1'b0;
		11793: rom = 1'b0;
		11794: rom = 1'b0;
		11795: rom = 1'b0;
		11796: rom = 1'b0;
		11797: rom = 1'b0;
		11798: rom = 1'b0;
		11799: rom = 1'b1;
		11800: rom = 1'b1;
		11801: rom = 1'b1;
		11802: rom = 1'b1;
		11803: rom = 1'b1;
		11804: rom = 1'b1;
		11805: rom = 1'b1;
		11806: rom = 1'b1;
		11807: rom = 1'b1;
		11808: rom = 1'b1;
		11809: rom = 1'b1;
		11810: rom = 1'b1;
		11811: rom = 1'b1;
		11812: rom = 1'b1;
		11813: rom = 1'b1;
		11814: rom = 1'b1;
		11815: rom = 1'b1;
		11816: rom = 1'b1;
		11817: rom = 1'b1;
		11818: rom = 1'b1;
		11819: rom = 1'b1;
		11820: rom = 1'b1;
		11821: rom = 1'b1;
		11822: rom = 1'b1;
		11823: rom = 1'b1;
		11824: rom = 1'b1;
		11825: rom = 1'b1;
		11826: rom = 1'b1;
		11827: rom = 1'b1;
		11828: rom = 1'b1;
		11829: rom = 1'b1;
		11830: rom = 1'b0;
		11831: rom = 1'b1;
		11832: rom = 1'b1;
		11833: rom = 1'b1;
		11834: rom = 1'b1;
		11835: rom = 1'b1;
		11836: rom = 1'b1;
		11837: rom = 1'b1;
		11838: rom = 1'b1;
		11839: rom = 1'b1;
		11840: rom = 1'b1;
		11841: rom = 1'b1;
		11842: rom = 1'b1;
		11843: rom = 1'b1;
		11844: rom = 1'b1;
		11845: rom = 1'b1;
		11846: rom = 1'b1;
		11847: rom = 1'b1;
		11848: rom = 1'b1;
		11849: rom = 1'b1;
		11850: rom = 1'b1;
		11851: rom = 1'b1;
		11852: rom = 1'b1;
		11853: rom = 1'b1;
		11854: rom = 1'b1;
		11855: rom = 1'b1;
		11856: rom = 1'b1;
		11857: rom = 1'b0;
		11858: rom = 1'b0;
		11859: rom = 1'b1;
		11860: rom = 1'b1;
		11861: rom = 1'b1;
		11862: rom = 1'b1;
		11863: rom = 1'b1;
		11864: rom = 1'b1;
		11865: rom = 1'b1;
		11866: rom = 1'b1;
		11867: rom = 1'b1;
		11868: rom = 1'b1;
		11869: rom = 1'b1;
		11870: rom = 1'b1;
		11871: rom = 1'b1;
		11872: rom = 1'b1;
		11873: rom = 1'b1;
		11874: rom = 1'b1;
		11875: rom = 1'b1;
		11876: rom = 1'b1;
		11877: rom = 1'b1;
		11878: rom = 1'b1;
		11879: rom = 1'b1;
		11880: rom = 1'b1;
		11881: rom = 1'b1;
		11882: rom = 1'b1;
		11883: rom = 1'b1;
		11884: rom = 1'b1;
		11885: rom = 1'b0;
		11886: rom = 1'b0;
		11887: rom = 1'b0;
		11888: rom = 1'b0;
		11889: rom = 1'b0;
		11890: rom = 1'b0;
		11891: rom = 1'b0;
		11892: rom = 1'b0;
		11893: rom = 1'b0;
		11894: rom = 1'b0;
		11895: rom = 1'b0;
		11896: rom = 1'b0;
		11897: rom = 1'b0;
		11898: rom = 1'b0;
		11899: rom = 1'b0;
		11900: rom = 1'b0;
		11901: rom = 1'b0;
		11902: rom = 1'b0;
		11903: rom = 1'b0;
		11904: rom = 1'b0;
		11905: rom = 1'b0;
		11906: rom = 1'b0;
		11907: rom = 1'b0;
		11908: rom = 1'b0;
		11909: rom = 1'b0;
		11910: rom = 1'b0;
		11911: rom = 1'b0;
		11912: rom = 1'b0;
		11913: rom = 1'b0;
		11914: rom = 1'b0;
		11915: rom = 1'b0;
		11916: rom = 1'b0;
		11917: rom = 1'b0;
		11918: rom = 1'b0;
		11919: rom = 1'b0;
		11920: rom = 1'b0;
		11921: rom = 1'b0;
		11922: rom = 1'b0;
		11923: rom = 1'b0;
		11924: rom = 1'b0;
		11925: rom = 1'b0;
		11926: rom = 1'b0;
		11927: rom = 1'b1;
		11928: rom = 1'b1;
		11929: rom = 1'b1;
		11930: rom = 1'b1;
		11931: rom = 1'b1;
		11932: rom = 1'b1;
		11933: rom = 1'b1;
		11934: rom = 1'b1;
		11935: rom = 1'b1;
		11936: rom = 1'b1;
		11937: rom = 1'b1;
		11938: rom = 1'b1;
		11939: rom = 1'b1;
		11940: rom = 1'b1;
		11941: rom = 1'b1;
		11942: rom = 1'b1;
		11943: rom = 1'b1;
		11944: rom = 1'b1;
		11945: rom = 1'b1;
		11946: rom = 1'b1;
		11947: rom = 1'b1;
		11948: rom = 1'b1;
		11949: rom = 1'b1;
		11950: rom = 1'b1;
		11951: rom = 1'b1;
		11952: rom = 1'b1;
		11953: rom = 1'b1;
		11954: rom = 1'b1;
		11955: rom = 1'b1;
		11956: rom = 1'b1;
		11957: rom = 1'b0;
		11958: rom = 1'b0;
		11959: rom = 1'b0;
		11960: rom = 1'b1;
		11961: rom = 1'b1;
		11962: rom = 1'b1;
		11963: rom = 1'b1;
		11964: rom = 1'b1;
		11965: rom = 1'b1;
		11966: rom = 1'b1;
		11967: rom = 1'b1;
		11968: rom = 1'b1;
		11969: rom = 1'b1;
		11970: rom = 1'b1;
		11971: rom = 1'b1;
		11972: rom = 1'b1;
		11973: rom = 1'b1;
		11974: rom = 1'b1;
		11975: rom = 1'b1;
		11976: rom = 1'b1;
		11977: rom = 1'b1;
		11978: rom = 1'b1;
		11979: rom = 1'b1;
		11980: rom = 1'b1;
		11981: rom = 1'b1;
		11982: rom = 1'b1;
		11983: rom = 1'b1;
		11984: rom = 1'b1;
		11985: rom = 1'b0;
		11986: rom = 1'b1;
		11987: rom = 1'b1;
		11988: rom = 1'b1;
		11989: rom = 1'b1;
		11990: rom = 1'b1;
		11991: rom = 1'b1;
		11992: rom = 1'b1;
		11993: rom = 1'b1;
		11994: rom = 1'b1;
		11995: rom = 1'b1;
		11996: rom = 1'b1;
		11997: rom = 1'b1;
		11998: rom = 1'b1;
		11999: rom = 1'b1;
		12000: rom = 1'b1;
		12001: rom = 1'b1;
		12002: rom = 1'b1;
		12003: rom = 1'b1;
		12004: rom = 1'b1;
		12005: rom = 1'b1;
		12006: rom = 1'b1;
		12007: rom = 1'b1;
		12008: rom = 1'b1;
		12009: rom = 1'b1;
		12010: rom = 1'b1;
		12011: rom = 1'b1;
		12012: rom = 1'b1;
		12013: rom = 1'b0;
		12014: rom = 1'b0;
		12015: rom = 1'b0;
		12016: rom = 1'b0;
		12017: rom = 1'b0;
		12018: rom = 1'b0;
		12019: rom = 1'b0;
		12020: rom = 1'b0;
		12021: rom = 1'b0;
		12022: rom = 1'b0;
		12023: rom = 1'b0;
		12024: rom = 1'b0;
		12025: rom = 1'b0;
		12026: rom = 1'b0;
		12027: rom = 1'b0;
		12028: rom = 1'b0;
		12029: rom = 1'b0;
		12030: rom = 1'b0;
		12031: rom = 1'b0;
		12032: rom = 1'b0;
		12033: rom = 1'b0;
		12034: rom = 1'b0;
		12035: rom = 1'b0;
		12036: rom = 1'b0;
		12037: rom = 1'b0;
		12038: rom = 1'b0;
		12039: rom = 1'b0;
		12040: rom = 1'b0;
		12041: rom = 1'b0;
		12042: rom = 1'b0;
		12043: rom = 1'b0;
		12044: rom = 1'b0;
		12045: rom = 1'b0;
		12046: rom = 1'b0;
		12047: rom = 1'b0;
		12048: rom = 1'b0;
		12049: rom = 1'b0;
		12050: rom = 1'b0;
		12051: rom = 1'b0;
		12052: rom = 1'b0;
		12053: rom = 1'b0;
		12054: rom = 1'b1;
		12055: rom = 1'b1;
		12056: rom = 1'b1;
		12057: rom = 1'b1;
		12058: rom = 1'b1;
		12059: rom = 1'b1;
		12060: rom = 1'b1;
		12061: rom = 1'b1;
		12062: rom = 1'b1;
		12063: rom = 1'b1;
		12064: rom = 1'b1;
		12065: rom = 1'b1;
		12066: rom = 1'b1;
		12067: rom = 1'b1;
		12068: rom = 1'b1;
		12069: rom = 1'b1;
		12070: rom = 1'b1;
		12071: rom = 1'b1;
		12072: rom = 1'b1;
		12073: rom = 1'b1;
		12074: rom = 1'b1;
		12075: rom = 1'b1;
		12076: rom = 1'b1;
		12077: rom = 1'b1;
		12078: rom = 1'b1;
		12079: rom = 1'b1;
		12080: rom = 1'b1;
		12081: rom = 1'b1;
		12082: rom = 1'b1;
		12083: rom = 1'b1;
		12084: rom = 1'b0;
		12085: rom = 1'b0;
		12086: rom = 1'b1;
		12087: rom = 1'b0;
		12088: rom = 1'b0;
		12089: rom = 1'b1;
		12090: rom = 1'b1;
		12091: rom = 1'b1;
		12092: rom = 1'b1;
		12093: rom = 1'b1;
		12094: rom = 1'b1;
		12095: rom = 1'b1;
		12096: rom = 1'b1;
		12097: rom = 1'b1;
		12098: rom = 1'b1;
		12099: rom = 1'b1;
		12100: rom = 1'b1;
		12101: rom = 1'b1;
		12102: rom = 1'b1;
		12103: rom = 1'b1;
		12104: rom = 1'b1;
		12105: rom = 1'b1;
		12106: rom = 1'b1;
		12107: rom = 1'b1;
		12108: rom = 1'b1;
		12109: rom = 1'b1;
		12110: rom = 1'b1;
		12111: rom = 1'b1;
		12112: rom = 1'b1;
		12113: rom = 1'b0;
		12114: rom = 1'b1;
		12115: rom = 1'b1;
		12116: rom = 1'b1;
		12117: rom = 1'b1;
		12118: rom = 1'b1;
		12119: rom = 1'b1;
		12120: rom = 1'b1;
		12121: rom = 1'b1;
		12122: rom = 1'b1;
		12123: rom = 1'b1;
		12124: rom = 1'b1;
		12125: rom = 1'b1;
		12126: rom = 1'b1;
		12127: rom = 1'b1;
		12128: rom = 1'b1;
		12129: rom = 1'b1;
		12130: rom = 1'b1;
		12131: rom = 1'b1;
		12132: rom = 1'b1;
		12133: rom = 1'b1;
		12134: rom = 1'b1;
		12135: rom = 1'b1;
		12136: rom = 1'b1;
		12137: rom = 1'b1;
		12138: rom = 1'b1;
		12139: rom = 1'b1;
		12140: rom = 1'b0;
		12141: rom = 1'b0;
		12142: rom = 1'b0;
		12143: rom = 1'b0;
		12144: rom = 1'b0;
		12145: rom = 1'b0;
		12146: rom = 1'b0;
		12147: rom = 1'b0;
		12148: rom = 1'b0;
		12149: rom = 1'b0;
		12150: rom = 1'b0;
		12151: rom = 1'b0;
		12152: rom = 1'b0;
		12153: rom = 1'b0;
		12154: rom = 1'b0;
		12155: rom = 1'b0;
		12156: rom = 1'b0;
		12157: rom = 1'b0;
		12158: rom = 1'b0;
		12159: rom = 1'b0;
		12160: rom = 1'b0;
		12161: rom = 1'b0;
		12162: rom = 1'b0;
		12163: rom = 1'b0;
		12164: rom = 1'b0;
		12165: rom = 1'b0;
		12166: rom = 1'b0;
		12167: rom = 1'b0;
		12168: rom = 1'b0;
		12169: rom = 1'b0;
		12170: rom = 1'b0;
		12171: rom = 1'b0;
		12172: rom = 1'b0;
		12173: rom = 1'b0;
		12174: rom = 1'b0;
		12175: rom = 1'b0;
		12176: rom = 1'b0;
		12177: rom = 1'b0;
		12178: rom = 1'b0;
		12179: rom = 1'b0;
		12180: rom = 1'b0;
		12181: rom = 1'b1;
		12182: rom = 1'b1;
		12183: rom = 1'b1;
		12184: rom = 1'b1;
		12185: rom = 1'b1;
		12186: rom = 1'b1;
		12187: rom = 1'b1;
		12188: rom = 1'b1;
		12189: rom = 1'b1;
		12190: rom = 1'b1;
		12191: rom = 1'b1;
		12192: rom = 1'b1;
		12193: rom = 1'b1;
		12194: rom = 1'b1;
		12195: rom = 1'b1;
		12196: rom = 1'b1;
		12197: rom = 1'b1;
		12198: rom = 1'b1;
		12199: rom = 1'b1;
		12200: rom = 1'b1;
		12201: rom = 1'b1;
		12202: rom = 1'b1;
		12203: rom = 1'b1;
		12204: rom = 1'b1;
		12205: rom = 1'b1;
		12206: rom = 1'b1;
		12207: rom = 1'b1;
		12208: rom = 1'b1;
		12209: rom = 1'b1;
		12210: rom = 1'b1;
		12211: rom = 1'b0;
		12212: rom = 1'b1;
		12213: rom = 1'b1;
		12214: rom = 1'b1;
		12215: rom = 1'b1;
		12216: rom = 1'b0;
		12217: rom = 1'b1;
		12218: rom = 1'b1;
		12219: rom = 1'b1;
		12220: rom = 1'b1;
		12221: rom = 1'b1;
		12222: rom = 1'b1;
		12223: rom = 1'b1;
		12224: rom = 1'b1;
		12225: rom = 1'b1;
		12226: rom = 1'b1;
		12227: rom = 1'b1;
		12228: rom = 1'b1;
		12229: rom = 1'b1;
		12230: rom = 1'b1;
		12231: rom = 1'b1;
		12232: rom = 1'b1;
		12233: rom = 1'b1;
		12234: rom = 1'b1;
		12235: rom = 1'b1;
		12236: rom = 1'b1;
		12237: rom = 1'b1;
		12238: rom = 1'b1;
		12239: rom = 1'b1;
		12240: rom = 1'b1;
		12241: rom = 1'b0;
		12242: rom = 1'b1;
		12243: rom = 1'b1;
		12244: rom = 1'b1;
		12245: rom = 1'b1;
		12246: rom = 1'b1;
		12247: rom = 1'b1;
		12248: rom = 1'b1;
		12249: rom = 1'b1;
		12250: rom = 1'b1;
		12251: rom = 1'b1;
		12252: rom = 1'b1;
		12253: rom = 1'b1;
		12254: rom = 1'b1;
		12255: rom = 1'b1;
		12256: rom = 1'b1;
		12257: rom = 1'b1;
		12258: rom = 1'b1;
		12259: rom = 1'b1;
		12260: rom = 1'b1;
		12261: rom = 1'b1;
		12262: rom = 1'b1;
		12263: rom = 1'b1;
		12264: rom = 1'b1;
		12265: rom = 1'b1;
		12266: rom = 1'b1;
		12267: rom = 1'b0;
		12268: rom = 1'b0;
		12269: rom = 1'b0;
		12270: rom = 1'b0;
		12271: rom = 1'b0;
		12272: rom = 1'b0;
		12273: rom = 1'b0;
		12274: rom = 1'b0;
		12275: rom = 1'b0;
		12276: rom = 1'b0;
		12277: rom = 1'b0;
		12278: rom = 1'b0;
		12279: rom = 1'b0;
		12280: rom = 1'b0;
		12281: rom = 1'b0;
		12282: rom = 1'b0;
		12283: rom = 1'b0;
		12284: rom = 1'b0;
		12285: rom = 1'b0;
		12286: rom = 1'b0;
		12287: rom = 1'b0;
		12288: rom = 1'b0;
		12289: rom = 1'b0;
		12290: rom = 1'b0;
		12291: rom = 1'b0;
		12292: rom = 1'b0;
		12293: rom = 1'b0;
		12294: rom = 1'b0;
		12295: rom = 1'b0;
		12296: rom = 1'b0;
		12297: rom = 1'b0;
		12298: rom = 1'b0;
		12299: rom = 1'b0;
		12300: rom = 1'b0;
		12301: rom = 1'b0;
		12302: rom = 1'b0;
		12303: rom = 1'b0;
		12304: rom = 1'b0;
		12305: rom = 1'b0;
		12306: rom = 1'b0;
		12307: rom = 1'b0;
		12308: rom = 1'b0;
		12309: rom = 1'b1;
		12310: rom = 1'b1;
		12311: rom = 1'b1;
		12312: rom = 1'b1;
		12313: rom = 1'b1;
		12314: rom = 1'b1;
		12315: rom = 1'b1;
		12316: rom = 1'b1;
		12317: rom = 1'b1;
		12318: rom = 1'b1;
		12319: rom = 1'b1;
		12320: rom = 1'b1;
		12321: rom = 1'b1;
		12322: rom = 1'b1;
		12323: rom = 1'b1;
		12324: rom = 1'b1;
		12325: rom = 1'b1;
		12326: rom = 1'b1;
		12327: rom = 1'b1;
		12328: rom = 1'b1;
		12329: rom = 1'b1;
		12330: rom = 1'b1;
		12331: rom = 1'b1;
		12332: rom = 1'b1;
		12333: rom = 1'b1;
		12334: rom = 1'b1;
		12335: rom = 1'b1;
		12336: rom = 1'b1;
		12337: rom = 1'b1;
		12338: rom = 1'b0;
		12339: rom = 1'b1;
		12340: rom = 1'b1;
		12341: rom = 1'b1;
		12342: rom = 1'b1;
		12343: rom = 1'b1;
		12344: rom = 1'b1;
		12345: rom = 1'b0;
		12346: rom = 1'b1;
		12347: rom = 1'b1;
		12348: rom = 1'b1;
		12349: rom = 1'b1;
		12350: rom = 1'b1;
		12351: rom = 1'b1;
		12352: rom = 1'b1;
		12353: rom = 1'b1;
		12354: rom = 1'b1;
		12355: rom = 1'b1;
		12356: rom = 1'b1;
		12357: rom = 1'b1;
		12358: rom = 1'b1;
		12359: rom = 1'b1;
		12360: rom = 1'b1;
		12361: rom = 1'b1;
		12362: rom = 1'b1;
		12363: rom = 1'b1;
		12364: rom = 1'b1;
		12365: rom = 1'b1;
		12366: rom = 1'b1;
		12367: rom = 1'b1;
		12368: rom = 1'b1;
		12369: rom = 1'b0;
		12370: rom = 1'b1;
		12371: rom = 1'b1;
		12372: rom = 1'b1;
		12373: rom = 1'b1;
		12374: rom = 1'b1;
		12375: rom = 1'b1;
		12376: rom = 1'b1;
		12377: rom = 1'b1;
		12378: rom = 1'b1;
		12379: rom = 1'b1;
		12380: rom = 1'b1;
		12381: rom = 1'b1;
		12382: rom = 1'b1;
		12383: rom = 1'b1;
		12384: rom = 1'b1;
		12385: rom = 1'b1;
		12386: rom = 1'b1;
		12387: rom = 1'b1;
		12388: rom = 1'b1;
		12389: rom = 1'b1;
		12390: rom = 1'b1;
		12391: rom = 1'b1;
		12392: rom = 1'b1;
		12393: rom = 1'b1;
		12394: rom = 1'b1;
		12395: rom = 1'b0;
		12396: rom = 1'b0;
		12397: rom = 1'b0;
		12398: rom = 1'b0;
		12399: rom = 1'b0;
		12400: rom = 1'b0;
		12401: rom = 1'b0;
		12402: rom = 1'b0;
		12403: rom = 1'b0;
		12404: rom = 1'b0;
		12405: rom = 1'b0;
		12406: rom = 1'b0;
		12407: rom = 1'b0;
		12408: rom = 1'b0;
		12409: rom = 1'b0;
		12410: rom = 1'b0;
		12411: rom = 1'b0;
		12412: rom = 1'b0;
		12413: rom = 1'b0;
		12414: rom = 1'b0;
		12415: rom = 1'b0;
		12416: rom = 1'b0;
		12417: rom = 1'b0;
		12418: rom = 1'b0;
		12419: rom = 1'b0;
		12420: rom = 1'b0;
		12421: rom = 1'b0;
		12422: rom = 1'b0;
		12423: rom = 1'b0;
		12424: rom = 1'b0;
		12425: rom = 1'b0;
		12426: rom = 1'b0;
		12427: rom = 1'b0;
		12428: rom = 1'b0;
		12429: rom = 1'b0;
		12430: rom = 1'b0;
		12431: rom = 1'b0;
		12432: rom = 1'b0;
		12433: rom = 1'b0;
		12434: rom = 1'b0;
		12435: rom = 1'b0;
		12436: rom = 1'b1;
		12437: rom = 1'b1;
		12438: rom = 1'b1;
		12439: rom = 1'b1;
		12440: rom = 1'b1;
		12441: rom = 1'b1;
		12442: rom = 1'b1;
		12443: rom = 1'b1;
		12444: rom = 1'b1;
		12445: rom = 1'b1;
		12446: rom = 1'b1;
		12447: rom = 1'b1;
		12448: rom = 1'b1;
		12449: rom = 1'b1;
		12450: rom = 1'b1;
		12451: rom = 1'b1;
		12452: rom = 1'b1;
		12453: rom = 1'b1;
		12454: rom = 1'b1;
		12455: rom = 1'b1;
		12456: rom = 1'b1;
		12457: rom = 1'b1;
		12458: rom = 1'b1;
		12459: rom = 1'b1;
		12460: rom = 1'b1;
		12461: rom = 1'b1;
		12462: rom = 1'b1;
		12463: rom = 1'b1;
		12464: rom = 1'b1;
		12465: rom = 1'b0;
		12466: rom = 1'b0;
		12467: rom = 1'b1;
		12468: rom = 1'b1;
		12469: rom = 1'b1;
		12470: rom = 1'b1;
		12471: rom = 1'b1;
		12472: rom = 1'b1;
		12473: rom = 1'b0;
		12474: rom = 1'b0;
		12475: rom = 1'b1;
		12476: rom = 1'b1;
		12477: rom = 1'b1;
		12478: rom = 1'b1;
		12479: rom = 1'b1;
		12480: rom = 1'b1;
		12481: rom = 1'b1;
		12482: rom = 1'b1;
		12483: rom = 1'b1;
		12484: rom = 1'b1;
		12485: rom = 1'b1;
		12486: rom = 1'b1;
		12487: rom = 1'b1;
		12488: rom = 1'b1;
		12489: rom = 1'b1;
		12490: rom = 1'b1;
		12491: rom = 1'b1;
		12492: rom = 1'b1;
		12493: rom = 1'b1;
		12494: rom = 1'b1;
		12495: rom = 1'b1;
		12496: rom = 1'b0;
		12497: rom = 1'b0;
		12498: rom = 1'b1;
		12499: rom = 1'b1;
		12500: rom = 1'b1;
		12501: rom = 1'b1;
		12502: rom = 1'b1;
		12503: rom = 1'b1;
		12504: rom = 1'b1;
		12505: rom = 1'b1;
		12506: rom = 1'b1;
		12507: rom = 1'b1;
		12508: rom = 1'b1;
		12509: rom = 1'b1;
		12510: rom = 1'b1;
		12511: rom = 1'b1;
		12512: rom = 1'b1;
		12513: rom = 1'b1;
		12514: rom = 1'b1;
		12515: rom = 1'b1;
		12516: rom = 1'b1;
		12517: rom = 1'b1;
		12518: rom = 1'b1;
		12519: rom = 1'b1;
		12520: rom = 1'b1;
		12521: rom = 1'b1;
		12522: rom = 1'b0;
		12523: rom = 1'b0;
		12524: rom = 1'b0;
		12525: rom = 1'b0;
		12526: rom = 1'b0;
		12527: rom = 1'b0;
		12528: rom = 1'b0;
		12529: rom = 1'b0;
		12530: rom = 1'b0;
		12531: rom = 1'b0;
		12532: rom = 1'b0;
		12533: rom = 1'b0;
		12534: rom = 1'b0;
		12535: rom = 1'b0;
		12536: rom = 1'b0;
		12537: rom = 1'b0;
		12538: rom = 1'b0;
		12539: rom = 1'b0;
		12540: rom = 1'b0;
		12541: rom = 1'b0;
		12542: rom = 1'b0;
		12543: rom = 1'b0;
		12544: rom = 1'b0;
		12545: rom = 1'b0;
		12546: rom = 1'b0;
		12547: rom = 1'b0;
		12548: rom = 1'b0;
		12549: rom = 1'b0;
		12550: rom = 1'b0;
		12551: rom = 1'b0;
		12552: rom = 1'b0;
		12553: rom = 1'b0;
		12554: rom = 1'b0;
		12555: rom = 1'b0;
		12556: rom = 1'b0;
		12557: rom = 1'b0;
		12558: rom = 1'b0;
		12559: rom = 1'b0;
		12560: rom = 1'b0;
		12561: rom = 1'b0;
		12562: rom = 1'b0;
		12563: rom = 1'b0;
		12564: rom = 1'b1;
		12565: rom = 1'b1;
		12566: rom = 1'b1;
		12567: rom = 1'b1;
		12568: rom = 1'b1;
		12569: rom = 1'b1;
		12570: rom = 1'b1;
		12571: rom = 1'b1;
		12572: rom = 1'b1;
		12573: rom = 1'b1;
		12574: rom = 1'b1;
		12575: rom = 1'b1;
		12576: rom = 1'b1;
		12577: rom = 1'b1;
		12578: rom = 1'b1;
		12579: rom = 1'b1;
		12580: rom = 1'b1;
		12581: rom = 1'b1;
		12582: rom = 1'b1;
		12583: rom = 1'b1;
		12584: rom = 1'b1;
		12585: rom = 1'b1;
		12586: rom = 1'b1;
		12587: rom = 1'b1;
		12588: rom = 1'b1;
		12589: rom = 1'b1;
		12590: rom = 1'b1;
		12591: rom = 1'b1;
		12592: rom = 1'b1;
		12593: rom = 1'b0;
		12594: rom = 1'b1;
		12595: rom = 1'b1;
		12596: rom = 1'b1;
		12597: rom = 1'b1;
		12598: rom = 1'b1;
		12599: rom = 1'b1;
		12600: rom = 1'b1;
		12601: rom = 1'b1;
		12602: rom = 1'b0;
		12603: rom = 1'b0;
		12604: rom = 1'b1;
		12605: rom = 1'b1;
		12606: rom = 1'b1;
		12607: rom = 1'b1;
		12608: rom = 1'b1;
		12609: rom = 1'b1;
		12610: rom = 1'b1;
		12611: rom = 1'b1;
		12612: rom = 1'b1;
		12613: rom = 1'b1;
		12614: rom = 1'b1;
		12615: rom = 1'b1;
		12616: rom = 1'b1;
		12617: rom = 1'b1;
		12618: rom = 1'b1;
		12619: rom = 1'b1;
		12620: rom = 1'b1;
		12621: rom = 1'b1;
		12622: rom = 1'b1;
		12623: rom = 1'b1;
		12624: rom = 1'b0;
		12625: rom = 1'b0;
		12626: rom = 1'b1;
		12627: rom = 1'b1;
		12628: rom = 1'b1;
		12629: rom = 1'b1;
		12630: rom = 1'b1;
		12631: rom = 1'b1;
		12632: rom = 1'b1;
		12633: rom = 1'b1;
		12634: rom = 1'b1;
		12635: rom = 1'b1;
		12636: rom = 1'b1;
		12637: rom = 1'b1;
		12638: rom = 1'b1;
		12639: rom = 1'b1;
		12640: rom = 1'b1;
		12641: rom = 1'b1;
		12642: rom = 1'b1;
		12643: rom = 1'b1;
		12644: rom = 1'b1;
		12645: rom = 1'b1;
		12646: rom = 1'b1;
		12647: rom = 1'b1;
		12648: rom = 1'b1;
		12649: rom = 1'b1;
		12650: rom = 1'b0;
		12651: rom = 1'b0;
		12652: rom = 1'b0;
		12653: rom = 1'b0;
		12654: rom = 1'b0;
		12655: rom = 1'b0;
		12656: rom = 1'b0;
		12657: rom = 1'b0;
		12658: rom = 1'b0;
		12659: rom = 1'b0;
		12660: rom = 1'b0;
		12661: rom = 1'b0;
		12662: rom = 1'b0;
		12663: rom = 1'b0;
		12664: rom = 1'b0;
		12665: rom = 1'b0;
		12666: rom = 1'b0;
		12667: rom = 1'b0;
		12668: rom = 1'b0;
		12669: rom = 1'b0;
		12670: rom = 1'b0;
		12671: rom = 1'b0;
		12672: rom = 1'b0;
		12673: rom = 1'b0;
		12674: rom = 1'b0;
		12675: rom = 1'b0;
		12676: rom = 1'b0;
		12677: rom = 1'b0;
		12678: rom = 1'b0;
		12679: rom = 1'b0;
		12680: rom = 1'b0;
		12681: rom = 1'b0;
		12682: rom = 1'b0;
		12683: rom = 1'b0;
		12684: rom = 1'b0;
		12685: rom = 1'b0;
		12686: rom = 1'b0;
		12687: rom = 1'b0;
		12688: rom = 1'b0;
		12689: rom = 1'b0;
		12690: rom = 1'b0;
		12691: rom = 1'b0;
		12692: rom = 1'b1;
		12693: rom = 1'b1;
		12694: rom = 1'b1;
		12695: rom = 1'b1;
		12696: rom = 1'b1;
		12697: rom = 1'b1;
		12698: rom = 1'b1;
		12699: rom = 1'b1;
		12700: rom = 1'b1;
		12701: rom = 1'b1;
		12702: rom = 1'b1;
		12703: rom = 1'b1;
		12704: rom = 1'b1;
		12705: rom = 1'b1;
		12706: rom = 1'b1;
		12707: rom = 1'b1;
		12708: rom = 1'b1;
		12709: rom = 1'b1;
		12710: rom = 1'b1;
		12711: rom = 1'b1;
		12712: rom = 1'b1;
		12713: rom = 1'b1;
		12714: rom = 1'b1;
		12715: rom = 1'b1;
		12716: rom = 1'b1;
		12717: rom = 1'b1;
		12718: rom = 1'b1;
		12719: rom = 1'b1;
		12720: rom = 1'b0;
		12721: rom = 1'b1;
		12722: rom = 1'b1;
		12723: rom = 1'b1;
		12724: rom = 1'b1;
		12725: rom = 1'b1;
		12726: rom = 1'b1;
		12727: rom = 1'b1;
		12728: rom = 1'b1;
		12729: rom = 1'b1;
		12730: rom = 1'b1;
		12731: rom = 1'b0;
		12732: rom = 1'b0;
		12733: rom = 1'b1;
		12734: rom = 1'b1;
		12735: rom = 1'b1;
		12736: rom = 1'b1;
		12737: rom = 1'b1;
		12738: rom = 1'b1;
		12739: rom = 1'b1;
		12740: rom = 1'b1;
		12741: rom = 1'b1;
		12742: rom = 1'b1;
		12743: rom = 1'b1;
		12744: rom = 1'b1;
		12745: rom = 1'b1;
		12746: rom = 1'b1;
		12747: rom = 1'b1;
		12748: rom = 1'b1;
		12749: rom = 1'b1;
		12750: rom = 1'b1;
		12751: rom = 1'b1;
		12752: rom = 1'b0;
		12753: rom = 1'b0;
		12754: rom = 1'b1;
		12755: rom = 1'b1;
		12756: rom = 1'b1;
		12757: rom = 1'b1;
		12758: rom = 1'b1;
		12759: rom = 1'b1;
		12760: rom = 1'b1;
		12761: rom = 1'b1;
		12762: rom = 1'b1;
		12763: rom = 1'b1;
		12764: rom = 1'b1;
		12765: rom = 1'b1;
		12766: rom = 1'b1;
		12767: rom = 1'b1;
		12768: rom = 1'b1;
		12769: rom = 1'b1;
		12770: rom = 1'b1;
		12771: rom = 1'b1;
		12772: rom = 1'b1;
		12773: rom = 1'b1;
		12774: rom = 1'b1;
		12775: rom = 1'b1;
		12776: rom = 1'b1;
		12777: rom = 1'b0;
		12778: rom = 1'b0;
		12779: rom = 1'b0;
		12780: rom = 1'b0;
		12781: rom = 1'b0;
		12782: rom = 1'b0;
		12783: rom = 1'b0;
		12784: rom = 1'b0;
		12785: rom = 1'b0;
		12786: rom = 1'b0;
		12787: rom = 1'b0;
		12788: rom = 1'b0;
		12789: rom = 1'b0;
		12790: rom = 1'b0;
		12791: rom = 1'b0;
		12792: rom = 1'b0;
		12793: rom = 1'b0;
		12794: rom = 1'b0;
		12795: rom = 1'b0;
		12796: rom = 1'b0;
		12797: rom = 1'b0;
		12798: rom = 1'b0;
		12799: rom = 1'b0;
		12800: rom = 1'b0;
		12801: rom = 1'b0;
		12802: rom = 1'b0;
		12803: rom = 1'b0;
		12804: rom = 1'b0;
		12805: rom = 1'b0;
		12806: rom = 1'b0;
		12807: rom = 1'b0;
		12808: rom = 1'b0;
		12809: rom = 1'b0;
		12810: rom = 1'b0;
		12811: rom = 1'b0;
		12812: rom = 1'b0;
		12813: rom = 1'b0;
		12814: rom = 1'b0;
		12815: rom = 1'b0;
		12816: rom = 1'b0;
		12817: rom = 1'b0;
		12818: rom = 1'b0;
		12819: rom = 1'b1;
		12820: rom = 1'b1;
		12821: rom = 1'b1;
		12822: rom = 1'b1;
		12823: rom = 1'b1;
		12824: rom = 1'b1;
		12825: rom = 1'b1;
		12826: rom = 1'b1;
		12827: rom = 1'b1;
		12828: rom = 1'b1;
		12829: rom = 1'b1;
		12830: rom = 1'b1;
		12831: rom = 1'b1;
		12832: rom = 1'b1;
		12833: rom = 1'b1;
		12834: rom = 1'b1;
		12835: rom = 1'b1;
		12836: rom = 1'b1;
		12837: rom = 1'b1;
		12838: rom = 1'b1;
		12839: rom = 1'b1;
		12840: rom = 1'b1;
		12841: rom = 1'b1;
		12842: rom = 1'b1;
		12843: rom = 1'b1;
		12844: rom = 1'b1;
		12845: rom = 1'b1;
		12846: rom = 1'b1;
		12847: rom = 1'b0;
		12848: rom = 1'b0;
		12849: rom = 1'b1;
		12850: rom = 1'b1;
		12851: rom = 1'b1;
		12852: rom = 1'b1;
		12853: rom = 1'b1;
		12854: rom = 1'b1;
		12855: rom = 1'b1;
		12856: rom = 1'b1;
		12857: rom = 1'b1;
		12858: rom = 1'b1;
		12859: rom = 1'b1;
		12860: rom = 1'b0;
		12861: rom = 1'b0;
		12862: rom = 1'b1;
		12863: rom = 1'b1;
		12864: rom = 1'b1;
		12865: rom = 1'b1;
		12866: rom = 1'b1;
		12867: rom = 1'b1;
		12868: rom = 1'b1;
		12869: rom = 1'b1;
		12870: rom = 1'b1;
		12871: rom = 1'b1;
		12872: rom = 1'b1;
		12873: rom = 1'b1;
		12874: rom = 1'b1;
		12875: rom = 1'b1;
		12876: rom = 1'b1;
		12877: rom = 1'b1;
		12878: rom = 1'b1;
		12879: rom = 1'b1;
		12880: rom = 1'b0;
		12881: rom = 1'b0;
		12882: rom = 1'b1;
		12883: rom = 1'b1;
		12884: rom = 1'b1;
		12885: rom = 1'b1;
		12886: rom = 1'b1;
		12887: rom = 1'b1;
		12888: rom = 1'b1;
		12889: rom = 1'b1;
		12890: rom = 1'b1;
		12891: rom = 1'b1;
		12892: rom = 1'b1;
		12893: rom = 1'b1;
		12894: rom = 1'b1;
		12895: rom = 1'b1;
		12896: rom = 1'b1;
		12897: rom = 1'b1;
		12898: rom = 1'b1;
		12899: rom = 1'b1;
		12900: rom = 1'b1;
		12901: rom = 1'b1;
		12902: rom = 1'b1;
		12903: rom = 1'b1;
		12904: rom = 1'b1;
		12905: rom = 1'b0;
		12906: rom = 1'b0;
		12907: rom = 1'b0;
		12908: rom = 1'b0;
		12909: rom = 1'b0;
		12910: rom = 1'b0;
		12911: rom = 1'b0;
		12912: rom = 1'b0;
		12913: rom = 1'b0;
		12914: rom = 1'b0;
		12915: rom = 1'b0;
		12916: rom = 1'b0;
		12917: rom = 1'b0;
		12918: rom = 1'b0;
		12919: rom = 1'b0;
		12920: rom = 1'b0;
		12921: rom = 1'b0;
		12922: rom = 1'b0;
		12923: rom = 1'b0;
		12924: rom = 1'b0;
		12925: rom = 1'b0;
		12926: rom = 1'b0;
		12927: rom = 1'b0;
		12928: rom = 1'b0;
		12929: rom = 1'b0;
		12930: rom = 1'b0;
		12931: rom = 1'b0;
		12932: rom = 1'b0;
		12933: rom = 1'b0;
		12934: rom = 1'b0;
		12935: rom = 1'b0;
		12936: rom = 1'b0;
		12937: rom = 1'b0;
		12938: rom = 1'b0;
		12939: rom = 1'b0;
		12940: rom = 1'b0;
		12941: rom = 1'b0;
		12942: rom = 1'b0;
		12943: rom = 1'b0;
		12944: rom = 1'b0;
		12945: rom = 1'b0;
		12946: rom = 1'b0;
		12947: rom = 1'b1;
		12948: rom = 1'b1;
		12949: rom = 1'b1;
		12950: rom = 1'b1;
		12951: rom = 1'b1;
		12952: rom = 1'b1;
		12953: rom = 1'b1;
		12954: rom = 1'b1;
		12955: rom = 1'b1;
		12956: rom = 1'b1;
		12957: rom = 1'b1;
		12958: rom = 1'b1;
		12959: rom = 1'b1;
		12960: rom = 1'b1;
		12961: rom = 1'b1;
		12962: rom = 1'b1;
		12963: rom = 1'b1;
		12964: rom = 1'b1;
		12965: rom = 1'b1;
		12966: rom = 1'b1;
		12967: rom = 1'b1;
		12968: rom = 1'b1;
		12969: rom = 1'b1;
		12970: rom = 1'b1;
		12971: rom = 1'b1;
		12972: rom = 1'b1;
		12973: rom = 1'b1;
		12974: rom = 1'b1;
		12975: rom = 1'b0;
		12976: rom = 1'b1;
		12977: rom = 1'b1;
		12978: rom = 1'b1;
		12979: rom = 1'b1;
		12980: rom = 1'b1;
		12981: rom = 1'b1;
		12982: rom = 1'b1;
		12983: rom = 1'b1;
		12984: rom = 1'b1;
		12985: rom = 1'b1;
		12986: rom = 1'b1;
		12987: rom = 1'b1;
		12988: rom = 1'b1;
		12989: rom = 1'b0;
		12990: rom = 1'b0;
		12991: rom = 1'b1;
		12992: rom = 1'b1;
		12993: rom = 1'b1;
		12994: rom = 1'b1;
		12995: rom = 1'b1;
		12996: rom = 1'b1;
		12997: rom = 1'b1;
		12998: rom = 1'b1;
		12999: rom = 1'b1;
		13000: rom = 1'b1;
		13001: rom = 1'b1;
		13002: rom = 1'b1;
		13003: rom = 1'b1;
		13004: rom = 1'b1;
		13005: rom = 1'b1;
		13006: rom = 1'b1;
		13007: rom = 1'b1;
		13008: rom = 1'b0;
		13009: rom = 1'b0;
		13010: rom = 1'b1;
		13011: rom = 1'b1;
		13012: rom = 1'b1;
		13013: rom = 1'b1;
		13014: rom = 1'b1;
		13015: rom = 1'b1;
		13016: rom = 1'b1;
		13017: rom = 1'b1;
		13018: rom = 1'b1;
		13019: rom = 1'b1;
		13020: rom = 1'b1;
		13021: rom = 1'b1;
		13022: rom = 1'b1;
		13023: rom = 1'b1;
		13024: rom = 1'b1;
		13025: rom = 1'b1;
		13026: rom = 1'b1;
		13027: rom = 1'b1;
		13028: rom = 1'b1;
		13029: rom = 1'b1;
		13030: rom = 1'b1;
		13031: rom = 1'b1;
		13032: rom = 1'b0;
		13033: rom = 1'b0;
		13034: rom = 1'b0;
		13035: rom = 1'b0;
		13036: rom = 1'b0;
		13037: rom = 1'b0;
		13038: rom = 1'b0;
		13039: rom = 1'b0;
		13040: rom = 1'b0;
		13041: rom = 1'b0;
		13042: rom = 1'b0;
		13043: rom = 1'b0;
		13044: rom = 1'b0;
		13045: rom = 1'b0;
		13046: rom = 1'b0;
		13047: rom = 1'b0;
		13048: rom = 1'b0;
		13049: rom = 1'b0;
		13050: rom = 1'b0;
		13051: rom = 1'b0;
		13052: rom = 1'b0;
		13053: rom = 1'b0;
		13054: rom = 1'b0;
		13055: rom = 1'b0;
		13056: rom = 1'b0;
		13057: rom = 1'b0;
		13058: rom = 1'b0;
		13059: rom = 1'b0;
		13060: rom = 1'b0;
		13061: rom = 1'b0;
		13062: rom = 1'b0;
		13063: rom = 1'b0;
		13064: rom = 1'b0;
		13065: rom = 1'b0;
		13066: rom = 1'b0;
		13067: rom = 1'b0;
		13068: rom = 1'b0;
		13069: rom = 1'b0;
		13070: rom = 1'b0;
		13071: rom = 1'b0;
		13072: rom = 1'b0;
		13073: rom = 1'b0;
		13074: rom = 1'b1;
		13075: rom = 1'b1;
		13076: rom = 1'b1;
		13077: rom = 1'b1;
		13078: rom = 1'b1;
		13079: rom = 1'b1;
		13080: rom = 1'b1;
		13081: rom = 1'b1;
		13082: rom = 1'b1;
		13083: rom = 1'b1;
		13084: rom = 1'b1;
		13085: rom = 1'b1;
		13086: rom = 1'b1;
		13087: rom = 1'b1;
		13088: rom = 1'b1;
		13089: rom = 1'b1;
		13090: rom = 1'b1;
		13091: rom = 1'b1;
		13092: rom = 1'b1;
		13093: rom = 1'b1;
		13094: rom = 1'b1;
		13095: rom = 1'b1;
		13096: rom = 1'b1;
		13097: rom = 1'b1;
		13098: rom = 1'b1;
		13099: rom = 1'b1;
		13100: rom = 1'b1;
		13101: rom = 1'b1;
		13102: rom = 1'b0;
		13103: rom = 1'b0;
		13104: rom = 1'b1;
		13105: rom = 1'b1;
		13106: rom = 1'b1;
		13107: rom = 1'b1;
		13108: rom = 1'b1;
		13109: rom = 1'b1;
		13110: rom = 1'b1;
		13111: rom = 1'b1;
		13112: rom = 1'b1;
		13113: rom = 1'b1;
		13114: rom = 1'b1;
		13115: rom = 1'b1;
		13116: rom = 1'b1;
		13117: rom = 1'b1;
		13118: rom = 1'b1;
		13119: rom = 1'b0;
		13120: rom = 1'b0;
		13121: rom = 1'b1;
		13122: rom = 1'b1;
		13123: rom = 1'b1;
		13124: rom = 1'b1;
		13125: rom = 1'b1;
		13126: rom = 1'b1;
		13127: rom = 1'b1;
		13128: rom = 1'b1;
		13129: rom = 1'b1;
		13130: rom = 1'b1;
		13131: rom = 1'b1;
		13132: rom = 1'b1;
		13133: rom = 1'b1;
		13134: rom = 1'b1;
		13135: rom = 1'b1;
		13136: rom = 1'b0;
		13137: rom = 1'b0;
		13138: rom = 1'b1;
		13139: rom = 1'b1;
		13140: rom = 1'b1;
		13141: rom = 1'b1;
		13142: rom = 1'b1;
		13143: rom = 1'b1;
		13144: rom = 1'b1;
		13145: rom = 1'b1;
		13146: rom = 1'b1;
		13147: rom = 1'b1;
		13148: rom = 1'b1;
		13149: rom = 1'b1;
		13150: rom = 1'b1;
		13151: rom = 1'b1;
		13152: rom = 1'b1;
		13153: rom = 1'b1;
		13154: rom = 1'b1;
		13155: rom = 1'b1;
		13156: rom = 1'b1;
		13157: rom = 1'b1;
		13158: rom = 1'b1;
		13159: rom = 1'b0;
		13160: rom = 1'b0;
		13161: rom = 1'b0;
		13162: rom = 1'b0;
		13163: rom = 1'b0;
		13164: rom = 1'b0;
		13165: rom = 1'b0;
		13166: rom = 1'b0;
		13167: rom = 1'b0;
		13168: rom = 1'b0;
		13169: rom = 1'b0;
		13170: rom = 1'b0;
		13171: rom = 1'b0;
		13172: rom = 1'b0;
		13173: rom = 1'b0;
		13174: rom = 1'b0;
		13175: rom = 1'b0;
		13176: rom = 1'b0;
		13177: rom = 1'b0;
		13178: rom = 1'b0;
		13179: rom = 1'b0;
		13180: rom = 1'b0;
		13181: rom = 1'b0;
		13182: rom = 1'b0;
		13183: rom = 1'b0;
		13184: rom = 1'b0;
		13185: rom = 1'b0;
		13186: rom = 1'b0;
		13187: rom = 1'b0;
		13188: rom = 1'b0;
		13189: rom = 1'b0;
		13190: rom = 1'b0;
		13191: rom = 1'b0;
		13192: rom = 1'b0;
		13193: rom = 1'b0;
		13194: rom = 1'b0;
		13195: rom = 1'b0;
		13196: rom = 1'b0;
		13197: rom = 1'b0;
		13198: rom = 1'b0;
		13199: rom = 1'b0;
		13200: rom = 1'b0;
		13201: rom = 1'b0;
		13202: rom = 1'b1;
		13203: rom = 1'b1;
		13204: rom = 1'b1;
		13205: rom = 1'b1;
		13206: rom = 1'b1;
		13207: rom = 1'b1;
		13208: rom = 1'b1;
		13209: rom = 1'b1;
		13210: rom = 1'b1;
		13211: rom = 1'b1;
		13212: rom = 1'b1;
		13213: rom = 1'b1;
		13214: rom = 1'b1;
		13215: rom = 1'b1;
		13216: rom = 1'b1;
		13217: rom = 1'b1;
		13218: rom = 1'b1;
		13219: rom = 1'b1;
		13220: rom = 1'b1;
		13221: rom = 1'b1;
		13222: rom = 1'b1;
		13223: rom = 1'b1;
		13224: rom = 1'b1;
		13225: rom = 1'b1;
		13226: rom = 1'b1;
		13227: rom = 1'b1;
		13228: rom = 1'b1;
		13229: rom = 1'b1;
		13230: rom = 1'b0;
		13231: rom = 1'b1;
		13232: rom = 1'b1;
		13233: rom = 1'b1;
		13234: rom = 1'b1;
		13235: rom = 1'b1;
		13236: rom = 1'b1;
		13237: rom = 1'b1;
		13238: rom = 1'b1;
		13239: rom = 1'b1;
		13240: rom = 1'b1;
		13241: rom = 1'b1;
		13242: rom = 1'b1;
		13243: rom = 1'b1;
		13244: rom = 1'b1;
		13245: rom = 1'b1;
		13246: rom = 1'b1;
		13247: rom = 1'b1;
		13248: rom = 1'b0;
		13249: rom = 1'b0;
		13250: rom = 1'b1;
		13251: rom = 1'b1;
		13252: rom = 1'b1;
		13253: rom = 1'b1;
		13254: rom = 1'b1;
		13255: rom = 1'b1;
		13256: rom = 1'b1;
		13257: rom = 1'b1;
		13258: rom = 1'b1;
		13259: rom = 1'b1;
		13260: rom = 1'b1;
		13261: rom = 1'b1;
		13262: rom = 1'b1;
		13263: rom = 1'b1;
		13264: rom = 1'b0;
		13265: rom = 1'b0;
		13266: rom = 1'b1;
		13267: rom = 1'b1;
		13268: rom = 1'b1;
		13269: rom = 1'b1;
		13270: rom = 1'b1;
		13271: rom = 1'b1;
		13272: rom = 1'b1;
		13273: rom = 1'b1;
		13274: rom = 1'b1;
		13275: rom = 1'b1;
		13276: rom = 1'b1;
		13277: rom = 1'b1;
		13278: rom = 1'b1;
		13279: rom = 1'b1;
		13280: rom = 1'b1;
		13281: rom = 1'b1;
		13282: rom = 1'b1;
		13283: rom = 1'b1;
		13284: rom = 1'b1;
		13285: rom = 1'b1;
		13286: rom = 1'b1;
		13287: rom = 1'b0;
		13288: rom = 1'b0;
		13289: rom = 1'b0;
		13290: rom = 1'b0;
		13291: rom = 1'b0;
		13292: rom = 1'b0;
		13293: rom = 1'b0;
		13294: rom = 1'b0;
		13295: rom = 1'b0;
		13296: rom = 1'b0;
		13297: rom = 1'b0;
		13298: rom = 1'b0;
		13299: rom = 1'b0;
		13300: rom = 1'b0;
		13301: rom = 1'b0;
		13302: rom = 1'b0;
		13303: rom = 1'b0;
		13304: rom = 1'b0;
		13305: rom = 1'b0;
		13306: rom = 1'b0;
		13307: rom = 1'b0;
		13308: rom = 1'b0;
		13309: rom = 1'b0;
		13310: rom = 1'b0;
		13311: rom = 1'b0;
		13312: rom = 1'b0;
		13313: rom = 1'b0;
		13314: rom = 1'b0;
		13315: rom = 1'b0;
		13316: rom = 1'b0;
		13317: rom = 1'b0;
		13318: rom = 1'b0;
		13319: rom = 1'b0;
		13320: rom = 1'b0;
		13321: rom = 1'b0;
		13322: rom = 1'b0;
		13323: rom = 1'b0;
		13324: rom = 1'b0;
		13325: rom = 1'b0;
		13326: rom = 1'b0;
		13327: rom = 1'b0;
		13328: rom = 1'b0;
		13329: rom = 1'b0;
		13330: rom = 1'b1;
		13331: rom = 1'b1;
		13332: rom = 1'b1;
		13333: rom = 1'b1;
		13334: rom = 1'b1;
		13335: rom = 1'b1;
		13336: rom = 1'b1;
		13337: rom = 1'b1;
		13338: rom = 1'b1;
		13339: rom = 1'b1;
		13340: rom = 1'b1;
		13341: rom = 1'b1;
		13342: rom = 1'b1;
		13343: rom = 1'b1;
		13344: rom = 1'b1;
		13345: rom = 1'b1;
		13346: rom = 1'b1;
		13347: rom = 1'b1;
		13348: rom = 1'b1;
		13349: rom = 1'b1;
		13350: rom = 1'b1;
		13351: rom = 1'b1;
		13352: rom = 1'b1;
		13353: rom = 1'b1;
		13354: rom = 1'b1;
		13355: rom = 1'b1;
		13356: rom = 1'b1;
		13357: rom = 1'b0;
		13358: rom = 1'b0;
		13359: rom = 1'b1;
		13360: rom = 1'b1;
		13361: rom = 1'b1;
		13362: rom = 1'b1;
		13363: rom = 1'b1;
		13364: rom = 1'b1;
		13365: rom = 1'b1;
		13366: rom = 1'b1;
		13367: rom = 1'b1;
		13368: rom = 1'b1;
		13369: rom = 1'b1;
		13370: rom = 1'b1;
		13371: rom = 1'b1;
		13372: rom = 1'b1;
		13373: rom = 1'b1;
		13374: rom = 1'b1;
		13375: rom = 1'b1;
		13376: rom = 1'b1;
		13377: rom = 1'b1;
		13378: rom = 1'b0;
		13379: rom = 1'b0;
		13380: rom = 1'b0;
		13381: rom = 1'b1;
		13382: rom = 1'b1;
		13383: rom = 1'b1;
		13384: rom = 1'b1;
		13385: rom = 1'b1;
		13386: rom = 1'b1;
		13387: rom = 1'b1;
		13388: rom = 1'b1;
		13389: rom = 1'b1;
		13390: rom = 1'b1;
		13391: rom = 1'b1;
		13392: rom = 1'b0;
		13393: rom = 1'b0;
		13394: rom = 1'b1;
		13395: rom = 1'b1;
		13396: rom = 1'b1;
		13397: rom = 1'b1;
		13398: rom = 1'b1;
		13399: rom = 1'b1;
		13400: rom = 1'b1;
		13401: rom = 1'b1;
		13402: rom = 1'b1;
		13403: rom = 1'b1;
		13404: rom = 1'b1;
		13405: rom = 1'b1;
		13406: rom = 1'b1;
		13407: rom = 1'b1;
		13408: rom = 1'b1;
		13409: rom = 1'b1;
		13410: rom = 1'b1;
		13411: rom = 1'b1;
		13412: rom = 1'b1;
		13413: rom = 1'b1;
		13414: rom = 1'b0;
		13415: rom = 1'b0;
		13416: rom = 1'b0;
		13417: rom = 1'b0;
		13418: rom = 1'b0;
		13419: rom = 1'b0;
		13420: rom = 1'b0;
		13421: rom = 1'b0;
		13422: rom = 1'b0;
		13423: rom = 1'b0;
		13424: rom = 1'b0;
		13425: rom = 1'b0;
		13426: rom = 1'b0;
		13427: rom = 1'b0;
		13428: rom = 1'b0;
		13429: rom = 1'b0;
		13430: rom = 1'b0;
		13431: rom = 1'b0;
		13432: rom = 1'b0;
		13433: rom = 1'b0;
		13434: rom = 1'b0;
		13435: rom = 1'b0;
		13436: rom = 1'b0;
		13437: rom = 1'b0;
		13438: rom = 1'b0;
		13439: rom = 1'b0;
		13440: rom = 1'b0;
		13441: rom = 1'b0;
		13442: rom = 1'b0;
		13443: rom = 1'b0;
		13444: rom = 1'b0;
		13445: rom = 1'b0;
		13446: rom = 1'b0;
		13447: rom = 1'b0;
		13448: rom = 1'b0;
		13449: rom = 1'b0;
		13450: rom = 1'b0;
		13451: rom = 1'b0;
		13452: rom = 1'b0;
		13453: rom = 1'b0;
		13454: rom = 1'b0;
		13455: rom = 1'b0;
		13456: rom = 1'b0;
		13457: rom = 1'b1;
		13458: rom = 1'b1;
		13459: rom = 1'b1;
		13460: rom = 1'b1;
		13461: rom = 1'b1;
		13462: rom = 1'b1;
		13463: rom = 1'b1;
		13464: rom = 1'b1;
		13465: rom = 1'b1;
		13466: rom = 1'b1;
		13467: rom = 1'b1;
		13468: rom = 1'b1;
		13469: rom = 1'b1;
		13470: rom = 1'b1;
		13471: rom = 1'b1;
		13472: rom = 1'b1;
		13473: rom = 1'b1;
		13474: rom = 1'b1;
		13475: rom = 1'b1;
		13476: rom = 1'b1;
		13477: rom = 1'b1;
		13478: rom = 1'b1;
		13479: rom = 1'b1;
		13480: rom = 1'b1;
		13481: rom = 1'b1;
		13482: rom = 1'b1;
		13483: rom = 1'b1;
		13484: rom = 1'b1;
		13485: rom = 1'b0;
		13486: rom = 1'b1;
		13487: rom = 1'b1;
		13488: rom = 1'b1;
		13489: rom = 1'b1;
		13490: rom = 1'b1;
		13491: rom = 1'b1;
		13492: rom = 1'b1;
		13493: rom = 1'b1;
		13494: rom = 1'b1;
		13495: rom = 1'b1;
		13496: rom = 1'b1;
		13497: rom = 1'b1;
		13498: rom = 1'b1;
		13499: rom = 1'b1;
		13500: rom = 1'b1;
		13501: rom = 1'b1;
		13502: rom = 1'b1;
		13503: rom = 1'b1;
		13504: rom = 1'b1;
		13505: rom = 1'b1;
		13506: rom = 1'b1;
		13507: rom = 1'b0;
		13508: rom = 1'b0;
		13509: rom = 1'b0;
		13510: rom = 1'b0;
		13511: rom = 1'b1;
		13512: rom = 1'b1;
		13513: rom = 1'b1;
		13514: rom = 1'b1;
		13515: rom = 1'b1;
		13516: rom = 1'b1;
		13517: rom = 1'b1;
		13518: rom = 1'b1;
		13519: rom = 1'b1;
		13520: rom = 1'b0;
		13521: rom = 1'b0;
		13522: rom = 1'b1;
		13523: rom = 1'b1;
		13524: rom = 1'b1;
		13525: rom = 1'b1;
		13526: rom = 1'b1;
		13527: rom = 1'b1;
		13528: rom = 1'b1;
		13529: rom = 1'b1;
		13530: rom = 1'b1;
		13531: rom = 1'b1;
		13532: rom = 1'b1;
		13533: rom = 1'b1;
		13534: rom = 1'b1;
		13535: rom = 1'b1;
		13536: rom = 1'b1;
		13537: rom = 1'b1;
		13538: rom = 1'b1;
		13539: rom = 1'b1;
		13540: rom = 1'b1;
		13541: rom = 1'b0;
		13542: rom = 1'b0;
		13543: rom = 1'b0;
		13544: rom = 1'b0;
		13545: rom = 1'b0;
		13546: rom = 1'b0;
		13547: rom = 1'b0;
		13548: rom = 1'b0;
		13549: rom = 1'b0;
		13550: rom = 1'b0;
		13551: rom = 1'b0;
		13552: rom = 1'b0;
		13553: rom = 1'b0;
		13554: rom = 1'b0;
		13555: rom = 1'b0;
		13556: rom = 1'b0;
		13557: rom = 1'b0;
		13558: rom = 1'b0;
		13559: rom = 1'b0;
		13560: rom = 1'b0;
		13561: rom = 1'b0;
		13562: rom = 1'b0;
		13563: rom = 1'b0;
		13564: rom = 1'b0;
		13565: rom = 1'b0;
		13566: rom = 1'b0;
		13567: rom = 1'b0;
		13568: rom = 1'b0;
		13569: rom = 1'b0;
		13570: rom = 1'b0;
		13571: rom = 1'b0;
		13572: rom = 1'b0;
		13573: rom = 1'b0;
		13574: rom = 1'b0;
		13575: rom = 1'b0;
		13576: rom = 1'b0;
		13577: rom = 1'b0;
		13578: rom = 1'b0;
		13579: rom = 1'b0;
		13580: rom = 1'b0;
		13581: rom = 1'b0;
		13582: rom = 1'b0;
		13583: rom = 1'b0;
		13584: rom = 1'b0;
		13585: rom = 1'b1;
		13586: rom = 1'b1;
		13587: rom = 1'b1;
		13588: rom = 1'b1;
		13589: rom = 1'b1;
		13590: rom = 1'b1;
		13591: rom = 1'b1;
		13592: rom = 1'b1;
		13593: rom = 1'b1;
		13594: rom = 1'b1;
		13595: rom = 1'b1;
		13596: rom = 1'b1;
		13597: rom = 1'b1;
		13598: rom = 1'b1;
		13599: rom = 1'b1;
		13600: rom = 1'b1;
		13601: rom = 1'b1;
		13602: rom = 1'b1;
		13603: rom = 1'b1;
		13604: rom = 1'b1;
		13605: rom = 1'b1;
		13606: rom = 1'b1;
		13607: rom = 1'b1;
		13608: rom = 1'b1;
		13609: rom = 1'b1;
		13610: rom = 1'b1;
		13611: rom = 1'b1;
		13612: rom = 1'b0;
		13613: rom = 1'b0;
		13614: rom = 1'b1;
		13615: rom = 1'b1;
		13616: rom = 1'b1;
		13617: rom = 1'b1;
		13618: rom = 1'b1;
		13619: rom = 1'b1;
		13620: rom = 1'b1;
		13621: rom = 1'b1;
		13622: rom = 1'b1;
		13623: rom = 1'b1;
		13624: rom = 1'b1;
		13625: rom = 1'b1;
		13626: rom = 1'b1;
		13627: rom = 1'b1;
		13628: rom = 1'b1;
		13629: rom = 1'b1;
		13630: rom = 1'b1;
		13631: rom = 1'b1;
		13632: rom = 1'b1;
		13633: rom = 1'b1;
		13634: rom = 1'b1;
		13635: rom = 1'b1;
		13636: rom = 1'b1;
		13637: rom = 1'b1;
		13638: rom = 1'b0;
		13639: rom = 1'b0;
		13640: rom = 1'b0;
		13641: rom = 1'b0;
		13642: rom = 1'b0;
		13643: rom = 1'b1;
		13644: rom = 1'b1;
		13645: rom = 1'b1;
		13646: rom = 1'b1;
		13647: rom = 1'b1;
		13648: rom = 1'b0;
		13649: rom = 1'b0;
		13650: rom = 1'b1;
		13651: rom = 1'b1;
		13652: rom = 1'b1;
		13653: rom = 1'b1;
		13654: rom = 1'b1;
		13655: rom = 1'b1;
		13656: rom = 1'b1;
		13657: rom = 1'b1;
		13658: rom = 1'b1;
		13659: rom = 1'b1;
		13660: rom = 1'b1;
		13661: rom = 1'b1;
		13662: rom = 1'b1;
		13663: rom = 1'b1;
		13664: rom = 1'b1;
		13665: rom = 1'b1;
		13666: rom = 1'b1;
		13667: rom = 1'b1;
		13668: rom = 1'b1;
		13669: rom = 1'b0;
		13670: rom = 1'b0;
		13671: rom = 1'b0;
		13672: rom = 1'b0;
		13673: rom = 1'b0;
		13674: rom = 1'b0;
		13675: rom = 1'b0;
		13676: rom = 1'b0;
		13677: rom = 1'b0;
		13678: rom = 1'b0;
		13679: rom = 1'b0;
		13680: rom = 1'b0;
		13681: rom = 1'b0;
		13682: rom = 1'b0;
		13683: rom = 1'b0;
		13684: rom = 1'b0;
		13685: rom = 1'b0;
		13686: rom = 1'b0;
		13687: rom = 1'b0;
		13688: rom = 1'b0;
		13689: rom = 1'b0;
		13690: rom = 1'b0;
		13691: rom = 1'b0;
		13692: rom = 1'b0;
		13693: rom = 1'b0;
		13694: rom = 1'b0;
		13695: rom = 1'b0;
		13696: rom = 1'b0;
		13697: rom = 1'b0;
		13698: rom = 1'b0;
		13699: rom = 1'b0;
		13700: rom = 1'b0;
		13701: rom = 1'b0;
		13702: rom = 1'b0;
		13703: rom = 1'b0;
		13704: rom = 1'b0;
		13705: rom = 1'b0;
		13706: rom = 1'b0;
		13707: rom = 1'b0;
		13708: rom = 1'b0;
		13709: rom = 1'b0;
		13710: rom = 1'b0;
		13711: rom = 1'b0;
		13712: rom = 1'b1;
		13713: rom = 1'b1;
		13714: rom = 1'b1;
		13715: rom = 1'b1;
		13716: rom = 1'b1;
		13717: rom = 1'b1;
		13718: rom = 1'b1;
		13719: rom = 1'b1;
		13720: rom = 1'b1;
		13721: rom = 1'b1;
		13722: rom = 1'b1;
		13723: rom = 1'b1;
		13724: rom = 1'b1;
		13725: rom = 1'b1;
		13726: rom = 1'b1;
		13727: rom = 1'b1;
		13728: rom = 1'b1;
		13729: rom = 1'b1;
		13730: rom = 1'b1;
		13731: rom = 1'b1;
		13732: rom = 1'b1;
		13733: rom = 1'b1;
		13734: rom = 1'b1;
		13735: rom = 1'b1;
		13736: rom = 1'b1;
		13737: rom = 1'b1;
		13738: rom = 1'b1;
		13739: rom = 1'b1;
		13740: rom = 1'b0;
		13741: rom = 1'b1;
		13742: rom = 1'b1;
		13743: rom = 1'b1;
		13744: rom = 1'b1;
		13745: rom = 1'b1;
		13746: rom = 1'b1;
		13747: rom = 1'b1;
		13748: rom = 1'b1;
		13749: rom = 1'b1;
		13750: rom = 1'b1;
		13751: rom = 1'b1;
		13752: rom = 1'b1;
		13753: rom = 1'b1;
		13754: rom = 1'b1;
		13755: rom = 1'b1;
		13756: rom = 1'b1;
		13757: rom = 1'b1;
		13758: rom = 1'b1;
		13759: rom = 1'b1;
		13760: rom = 1'b1;
		13761: rom = 1'b1;
		13762: rom = 1'b1;
		13763: rom = 1'b1;
		13764: rom = 1'b1;
		13765: rom = 1'b1;
		13766: rom = 1'b1;
		13767: rom = 1'b1;
		13768: rom = 1'b1;
		13769: rom = 1'b1;
		13770: rom = 1'b0;
		13771: rom = 1'b0;
		13772: rom = 1'b0;
		13773: rom = 1'b0;
		13774: rom = 1'b0;
		13775: rom = 1'b0;
		13776: rom = 1'b0;
		13777: rom = 1'b1;
		13778: rom = 1'b1;
		13779: rom = 1'b1;
		13780: rom = 1'b1;
		13781: rom = 1'b1;
		13782: rom = 1'b1;
		13783: rom = 1'b1;
		13784: rom = 1'b1;
		13785: rom = 1'b1;
		13786: rom = 1'b1;
		13787: rom = 1'b1;
		13788: rom = 1'b1;
		13789: rom = 1'b1;
		13790: rom = 1'b1;
		13791: rom = 1'b1;
		13792: rom = 1'b1;
		13793: rom = 1'b1;
		13794: rom = 1'b1;
		13795: rom = 1'b1;
		13796: rom = 1'b0;
		13797: rom = 1'b0;
		13798: rom = 1'b0;
		13799: rom = 1'b0;
		13800: rom = 1'b0;
		13801: rom = 1'b0;
		13802: rom = 1'b0;
		13803: rom = 1'b0;
		13804: rom = 1'b0;
		13805: rom = 1'b0;
		13806: rom = 1'b0;
		13807: rom = 1'b0;
		13808: rom = 1'b0;
		13809: rom = 1'b0;
		13810: rom = 1'b0;
		13811: rom = 1'b0;
		13812: rom = 1'b0;
		13813: rom = 1'b0;
		13814: rom = 1'b0;
		13815: rom = 1'b0;
		13816: rom = 1'b0;
		13817: rom = 1'b0;
		13818: rom = 1'b0;
		13819: rom = 1'b0;
		13820: rom = 1'b0;
		13821: rom = 1'b0;
		13822: rom = 1'b0;
		13823: rom = 1'b0;
		13824: rom = 1'b0;
		13825: rom = 1'b0;
		13826: rom = 1'b0;
		13827: rom = 1'b0;
		13828: rom = 1'b0;
		13829: rom = 1'b0;
		13830: rom = 1'b0;
		13831: rom = 1'b0;
		13832: rom = 1'b0;
		13833: rom = 1'b0;
		13834: rom = 1'b0;
		13835: rom = 1'b0;
		13836: rom = 1'b0;
		13837: rom = 1'b0;
		13838: rom = 1'b0;
		13839: rom = 1'b0;
		13840: rom = 1'b1;
		13841: rom = 1'b1;
		13842: rom = 1'b1;
		13843: rom = 1'b1;
		13844: rom = 1'b1;
		13845: rom = 1'b1;
		13846: rom = 1'b1;
		13847: rom = 1'b1;
		13848: rom = 1'b1;
		13849: rom = 1'b1;
		13850: rom = 1'b1;
		13851: rom = 1'b1;
		13852: rom = 1'b1;
		13853: rom = 1'b1;
		13854: rom = 1'b1;
		13855: rom = 1'b1;
		13856: rom = 1'b1;
		13857: rom = 1'b1;
		13858: rom = 1'b1;
		13859: rom = 1'b1;
		13860: rom = 1'b1;
		13861: rom = 1'b1;
		13862: rom = 1'b1;
		13863: rom = 1'b1;
		13864: rom = 1'b1;
		13865: rom = 1'b1;
		13866: rom = 1'b1;
		13867: rom = 1'b1;
		13868: rom = 1'b0;
		13869: rom = 1'b1;
		13870: rom = 1'b1;
		13871: rom = 1'b1;
		13872: rom = 1'b1;
		13873: rom = 1'b1;
		13874: rom = 1'b1;
		13875: rom = 1'b1;
		13876: rom = 1'b1;
		13877: rom = 1'b1;
		13878: rom = 1'b1;
		13879: rom = 1'b1;
		13880: rom = 1'b1;
		13881: rom = 1'b1;
		13882: rom = 1'b1;
		13883: rom = 1'b1;
		13884: rom = 1'b1;
		13885: rom = 1'b1;
		13886: rom = 1'b1;
		13887: rom = 1'b1;
		13888: rom = 1'b1;
		13889: rom = 1'b1;
		13890: rom = 1'b1;
		13891: rom = 1'b1;
		13892: rom = 1'b1;
		13893: rom = 1'b1;
		13894: rom = 1'b1;
		13895: rom = 1'b1;
		13896: rom = 1'b1;
		13897: rom = 1'b1;
		13898: rom = 1'b1;
		13899: rom = 1'b1;
		13900: rom = 1'b1;
		13901: rom = 1'b1;
		13902: rom = 1'b1;
		13903: rom = 1'b1;
		13904: rom = 1'b0;
		13905: rom = 1'b1;
		13906: rom = 1'b1;
		13907: rom = 1'b1;
		13908: rom = 1'b1;
		13909: rom = 1'b1;
		13910: rom = 1'b1;
		13911: rom = 1'b1;
		13912: rom = 1'b1;
		13913: rom = 1'b1;
		13914: rom = 1'b1;
		13915: rom = 1'b1;
		13916: rom = 1'b1;
		13917: rom = 1'b1;
		13918: rom = 1'b1;
		13919: rom = 1'b1;
		13920: rom = 1'b1;
		13921: rom = 1'b1;
		13922: rom = 1'b1;
		13923: rom = 1'b0;
		13924: rom = 1'b0;
		13925: rom = 1'b0;
		13926: rom = 1'b0;
		13927: rom = 1'b0;
		13928: rom = 1'b0;
		13929: rom = 1'b0;
		13930: rom = 1'b0;
		13931: rom = 1'b0;
		13932: rom = 1'b0;
		13933: rom = 1'b0;
		13934: rom = 1'b0;
		13935: rom = 1'b0;
		13936: rom = 1'b0;
		13937: rom = 1'b0;
		13938: rom = 1'b0;
		13939: rom = 1'b0;
		13940: rom = 1'b0;
		13941: rom = 1'b0;
		13942: rom = 1'b0;
		13943: rom = 1'b0;
		13944: rom = 1'b0;
		13945: rom = 1'b0;
		13946: rom = 1'b0;
		13947: rom = 1'b0;
		13948: rom = 1'b0;
		13949: rom = 1'b0;
		13950: rom = 1'b0;
		13951: rom = 1'b0;
		13952: rom = 1'b0;
		13953: rom = 1'b0;
		13954: rom = 1'b0;
		13955: rom = 1'b0;
		13956: rom = 1'b0;
		13957: rom = 1'b0;
		13958: rom = 1'b0;
		13959: rom = 1'b0;
		13960: rom = 1'b0;
		13961: rom = 1'b0;
		13962: rom = 1'b0;
		13963: rom = 1'b0;
		13964: rom = 1'b0;
		13965: rom = 1'b0;
		13966: rom = 1'b0;
		13967: rom = 1'b1;
		13968: rom = 1'b1;
		13969: rom = 1'b1;
		13970: rom = 1'b1;
		13971: rom = 1'b1;
		13972: rom = 1'b1;
		13973: rom = 1'b1;
		13974: rom = 1'b1;
		13975: rom = 1'b1;
		13976: rom = 1'b1;
		13977: rom = 1'b1;
		13978: rom = 1'b1;
		13979: rom = 1'b1;
		13980: rom = 1'b1;
		13981: rom = 1'b1;
		13982: rom = 1'b1;
		13983: rom = 1'b1;
		13984: rom = 1'b1;
		13985: rom = 1'b1;
		13986: rom = 1'b1;
		13987: rom = 1'b1;
		13988: rom = 1'b1;
		13989: rom = 1'b1;
		13990: rom = 1'b1;
		13991: rom = 1'b1;
		13992: rom = 1'b1;
		13993: rom = 1'b1;
		13994: rom = 1'b1;
		13995: rom = 1'b0;
		13996: rom = 1'b0;
		13997: rom = 1'b1;
		13998: rom = 1'b1;
		13999: rom = 1'b1;
		14000: rom = 1'b1;
		14001: rom = 1'b1;
		14002: rom = 1'b1;
		14003: rom = 1'b1;
		14004: rom = 1'b1;
		14005: rom = 1'b1;
		14006: rom = 1'b1;
		14007: rom = 1'b1;
		14008: rom = 1'b1;
		14009: rom = 1'b1;
		14010: rom = 1'b1;
		14011: rom = 1'b1;
		14012: rom = 1'b1;
		14013: rom = 1'b1;
		14014: rom = 1'b1;
		14015: rom = 1'b1;
		14016: rom = 1'b1;
		14017: rom = 1'b1;
		14018: rom = 1'b1;
		14019: rom = 1'b1;
		14020: rom = 1'b1;
		14021: rom = 1'b1;
		14022: rom = 1'b1;
		14023: rom = 1'b1;
		14024: rom = 1'b1;
		14025: rom = 1'b1;
		14026: rom = 1'b1;
		14027: rom = 1'b1;
		14028: rom = 1'b1;
		14029: rom = 1'b1;
		14030: rom = 1'b1;
		14031: rom = 1'b1;
		14032: rom = 1'b0;
		14033: rom = 1'b1;
		14034: rom = 1'b1;
		14035: rom = 1'b1;
		14036: rom = 1'b1;
		14037: rom = 1'b1;
		14038: rom = 1'b1;
		14039: rom = 1'b1;
		14040: rom = 1'b1;
		14041: rom = 1'b1;
		14042: rom = 1'b1;
		14043: rom = 1'b1;
		14044: rom = 1'b1;
		14045: rom = 1'b1;
		14046: rom = 1'b1;
		14047: rom = 1'b1;
		14048: rom = 1'b1;
		14049: rom = 1'b1;
		14050: rom = 1'b0;
		14051: rom = 1'b0;
		14052: rom = 1'b0;
		14053: rom = 1'b0;
		14054: rom = 1'b0;
		14055: rom = 1'b0;
		14056: rom = 1'b0;
		14057: rom = 1'b0;
		14058: rom = 1'b0;
		14059: rom = 1'b0;
		14060: rom = 1'b0;
		14061: rom = 1'b0;
		14062: rom = 1'b0;
		14063: rom = 1'b0;
		14064: rom = 1'b0;
		14065: rom = 1'b0;
		14066: rom = 1'b0;
		14067: rom = 1'b0;
		14068: rom = 1'b0;
		14069: rom = 1'b0;
		14070: rom = 1'b0;
		14071: rom = 1'b0;
		14072: rom = 1'b0;
		14073: rom = 1'b0;
		14074: rom = 1'b0;
		14075: rom = 1'b0;
		14076: rom = 1'b0;
		14077: rom = 1'b0;
		14078: rom = 1'b0;
		14079: rom = 1'b0;
		14080: rom = 1'b0;
		14081: rom = 1'b0;
		14082: rom = 1'b0;
		14083: rom = 1'b0;
		14084: rom = 1'b0;
		14085: rom = 1'b0;
		14086: rom = 1'b0;
		14087: rom = 1'b0;
		14088: rom = 1'b0;
		14089: rom = 1'b0;
		14090: rom = 1'b0;
		14091: rom = 1'b0;
		14092: rom = 1'b0;
		14093: rom = 1'b0;
		14094: rom = 1'b0;
		14095: rom = 1'b1;
		14096: rom = 1'b1;
		14097: rom = 1'b1;
		14098: rom = 1'b1;
		14099: rom = 1'b1;
		14100: rom = 1'b1;
		14101: rom = 1'b1;
		14102: rom = 1'b1;
		14103: rom = 1'b1;
		14104: rom = 1'b1;
		14105: rom = 1'b1;
		14106: rom = 1'b1;
		14107: rom = 1'b1;
		14108: rom = 1'b1;
		14109: rom = 1'b1;
		14110: rom = 1'b1;
		14111: rom = 1'b1;
		14112: rom = 1'b1;
		14113: rom = 1'b1;
		14114: rom = 1'b1;
		14115: rom = 1'b1;
		14116: rom = 1'b1;
		14117: rom = 1'b1;
		14118: rom = 1'b1;
		14119: rom = 1'b1;
		14120: rom = 1'b1;
		14121: rom = 1'b1;
		14122: rom = 1'b1;
		14123: rom = 1'b0;
		14124: rom = 1'b1;
		14125: rom = 1'b1;
		14126: rom = 1'b1;
		14127: rom = 1'b1;
		14128: rom = 1'b1;
		14129: rom = 1'b1;
		14130: rom = 1'b1;
		14131: rom = 1'b1;
		14132: rom = 1'b1;
		14133: rom = 1'b1;
		14134: rom = 1'b1;
		14135: rom = 1'b1;
		14136: rom = 1'b1;
		14137: rom = 1'b1;
		14138: rom = 1'b1;
		14139: rom = 1'b1;
		14140: rom = 1'b1;
		14141: rom = 1'b1;
		14142: rom = 1'b1;
		14143: rom = 1'b1;
		14144: rom = 1'b1;
		14145: rom = 1'b1;
		14146: rom = 1'b1;
		14147: rom = 1'b1;
		14148: rom = 1'b1;
		14149: rom = 1'b1;
		14150: rom = 1'b1;
		14151: rom = 1'b1;
		14152: rom = 1'b1;
		14153: rom = 1'b1;
		14154: rom = 1'b1;
		14155: rom = 1'b1;
		14156: rom = 1'b1;
		14157: rom = 1'b1;
		14158: rom = 1'b1;
		14159: rom = 1'b1;
		14160: rom = 1'b0;
		14161: rom = 1'b1;
		14162: rom = 1'b1;
		14163: rom = 1'b1;
		14164: rom = 1'b1;
		14165: rom = 1'b1;
		14166: rom = 1'b1;
		14167: rom = 1'b1;
		14168: rom = 1'b1;
		14169: rom = 1'b1;
		14170: rom = 1'b1;
		14171: rom = 1'b1;
		14172: rom = 1'b1;
		14173: rom = 1'b1;
		14174: rom = 1'b1;
		14175: rom = 1'b1;
		14176: rom = 1'b1;
		14177: rom = 1'b0;
		14178: rom = 1'b0;
		14179: rom = 1'b0;
		14180: rom = 1'b0;
		14181: rom = 1'b0;
		14182: rom = 1'b0;
		14183: rom = 1'b0;
		14184: rom = 1'b0;
		14185: rom = 1'b0;
		14186: rom = 1'b0;
		14187: rom = 1'b0;
		14188: rom = 1'b0;
		14189: rom = 1'b0;
		14190: rom = 1'b0;
		14191: rom = 1'b0;
		14192: rom = 1'b0;
		14193: rom = 1'b0;
		14194: rom = 1'b0;
		14195: rom = 1'b0;
		14196: rom = 1'b0;
		14197: rom = 1'b0;
		14198: rom = 1'b0;
		14199: rom = 1'b0;
		14200: rom = 1'b0;
		14201: rom = 1'b0;
		14202: rom = 1'b0;
		14203: rom = 1'b0;
		14204: rom = 1'b0;
		14205: rom = 1'b0;
		14206: rom = 1'b0;
		14207: rom = 1'b0;
		14208: rom = 1'b0;
		14209: rom = 1'b0;
		14210: rom = 1'b0;
		14211: rom = 1'b0;
		14212: rom = 1'b0;
		14213: rom = 1'b0;
		14214: rom = 1'b0;
		14215: rom = 1'b0;
		14216: rom = 1'b0;
		14217: rom = 1'b0;
		14218: rom = 1'b0;
		14219: rom = 1'b0;
		14220: rom = 1'b0;
		14221: rom = 1'b0;
		14222: rom = 1'b1;
		14223: rom = 1'b1;
		14224: rom = 1'b1;
		14225: rom = 1'b1;
		14226: rom = 1'b1;
		14227: rom = 1'b1;
		14228: rom = 1'b1;
		14229: rom = 1'b1;
		14230: rom = 1'b1;
		14231: rom = 1'b1;
		14232: rom = 1'b1;
		14233: rom = 1'b1;
		14234: rom = 1'b1;
		14235: rom = 1'b1;
		14236: rom = 1'b1;
		14237: rom = 1'b1;
		14238: rom = 1'b1;
		14239: rom = 1'b1;
		14240: rom = 1'b1;
		14241: rom = 1'b1;
		14242: rom = 1'b1;
		14243: rom = 1'b1;
		14244: rom = 1'b1;
		14245: rom = 1'b1;
		14246: rom = 1'b1;
		14247: rom = 1'b1;
		14248: rom = 1'b1;
		14249: rom = 1'b1;
		14250: rom = 1'b1;
		14251: rom = 1'b0;
		14252: rom = 1'b1;
		14253: rom = 1'b1;
		14254: rom = 1'b1;
		14255: rom = 1'b1;
		14256: rom = 1'b1;
		14257: rom = 1'b1;
		14258: rom = 1'b1;
		14259: rom = 1'b1;
		14260: rom = 1'b1;
		14261: rom = 1'b1;
		14262: rom = 1'b1;
		14263: rom = 1'b1;
		14264: rom = 1'b1;
		14265: rom = 1'b1;
		14266: rom = 1'b1;
		14267: rom = 1'b1;
		14268: rom = 1'b1;
		14269: rom = 1'b1;
		14270: rom = 1'b1;
		14271: rom = 1'b1;
		14272: rom = 1'b1;
		14273: rom = 1'b1;
		14274: rom = 1'b1;
		14275: rom = 1'b1;
		14276: rom = 1'b1;
		14277: rom = 1'b1;
		14278: rom = 1'b1;
		14279: rom = 1'b1;
		14280: rom = 1'b1;
		14281: rom = 1'b1;
		14282: rom = 1'b1;
		14283: rom = 1'b1;
		14284: rom = 1'b1;
		14285: rom = 1'b1;
		14286: rom = 1'b1;
		14287: rom = 1'b1;
		14288: rom = 1'b0;
		14289: rom = 1'b1;
		14290: rom = 1'b1;
		14291: rom = 1'b1;
		14292: rom = 1'b1;
		14293: rom = 1'b1;
		14294: rom = 1'b1;
		14295: rom = 1'b1;
		14296: rom = 1'b1;
		14297: rom = 1'b1;
		14298: rom = 1'b1;
		14299: rom = 1'b1;
		14300: rom = 1'b1;
		14301: rom = 1'b1;
		14302: rom = 1'b1;
		14303: rom = 1'b1;
		14304: rom = 1'b0;
		14305: rom = 1'b0;
		14306: rom = 1'b0;
		14307: rom = 1'b0;
		14308: rom = 1'b0;
		14309: rom = 1'b0;
		14310: rom = 1'b0;
		14311: rom = 1'b0;
		14312: rom = 1'b0;
		14313: rom = 1'b0;
		14314: rom = 1'b0;
		14315: rom = 1'b0;
		14316: rom = 1'b0;
		14317: rom = 1'b0;
		14318: rom = 1'b0;
		14319: rom = 1'b0;
		14320: rom = 1'b0;
		14321: rom = 1'b0;
		14322: rom = 1'b0;
		14323: rom = 1'b0;
		14324: rom = 1'b0;
		14325: rom = 1'b0;
		14326: rom = 1'b0;
		14327: rom = 1'b0;
		14328: rom = 1'b0;
		14329: rom = 1'b0;
		14330: rom = 1'b0;
		14331: rom = 1'b0;
		14332: rom = 1'b0;
		14333: rom = 1'b0;
		14334: rom = 1'b0;
		14335: rom = 1'b0;
		14336: rom = 1'b0;
		14337: rom = 1'b0;
		14338: rom = 1'b0;
		14339: rom = 1'b0;
		14340: rom = 1'b0;
		14341: rom = 1'b0;
		14342: rom = 1'b0;
		14343: rom = 1'b0;
		14344: rom = 1'b0;
		14345: rom = 1'b0;
		14346: rom = 1'b0;
		14347: rom = 1'b0;
		14348: rom = 1'b0;
		14349: rom = 1'b0;
		14350: rom = 1'b1;
		14351: rom = 1'b1;
		14352: rom = 1'b1;
		14353: rom = 1'b1;
		14354: rom = 1'b1;
		14355: rom = 1'b1;
		14356: rom = 1'b1;
		14357: rom = 1'b1;
		14358: rom = 1'b1;
		14359: rom = 1'b1;
		14360: rom = 1'b1;
		14361: rom = 1'b1;
		14362: rom = 1'b1;
		14363: rom = 1'b1;
		14364: rom = 1'b1;
		14365: rom = 1'b1;
		14366: rom = 1'b1;
		14367: rom = 1'b1;
		14368: rom = 1'b1;
		14369: rom = 1'b1;
		14370: rom = 1'b1;
		14371: rom = 1'b1;
		14372: rom = 1'b1;
		14373: rom = 1'b1;
		14374: rom = 1'b1;
		14375: rom = 1'b1;
		14376: rom = 1'b1;
		14377: rom = 1'b1;
		14378: rom = 1'b0;
		14379: rom = 1'b0;
		14380: rom = 1'b1;
		14381: rom = 1'b1;
		14382: rom = 1'b1;
		14383: rom = 1'b1;
		14384: rom = 1'b1;
		14385: rom = 1'b1;
		14386: rom = 1'b1;
		14387: rom = 1'b1;
		14388: rom = 1'b1;
		14389: rom = 1'b1;
		14390: rom = 1'b1;
		14391: rom = 1'b1;
		14392: rom = 1'b1;
		14393: rom = 1'b1;
		14394: rom = 1'b1;
		14395: rom = 1'b1;
		14396: rom = 1'b1;
		14397: rom = 1'b1;
		14398: rom = 1'b1;
		14399: rom = 1'b1;
		14400: rom = 1'b1;
		14401: rom = 1'b1;
		14402: rom = 1'b1;
		14403: rom = 1'b1;
		14404: rom = 1'b1;
		14405: rom = 1'b1;
		14406: rom = 1'b1;
		14407: rom = 1'b1;
		14408: rom = 1'b1;
		14409: rom = 1'b1;
		14410: rom = 1'b1;
		14411: rom = 1'b1;
		14412: rom = 1'b1;
		14413: rom = 1'b1;
		14414: rom = 1'b1;
		14415: rom = 1'b1;
		14416: rom = 1'b0;
		14417: rom = 1'b1;
		14418: rom = 1'b1;
		14419: rom = 1'b1;
		14420: rom = 1'b1;
		14421: rom = 1'b1;
		14422: rom = 1'b1;
		14423: rom = 1'b1;
		14424: rom = 1'b1;
		14425: rom = 1'b1;
		14426: rom = 1'b1;
		14427: rom = 1'b1;
		14428: rom = 1'b1;
		14429: rom = 1'b1;
		14430: rom = 1'b1;
		14431: rom = 1'b0;
		14432: rom = 1'b0;
		14433: rom = 1'b0;
		14434: rom = 1'b0;
		14435: rom = 1'b0;
		14436: rom = 1'b0;
		14437: rom = 1'b0;
		14438: rom = 1'b0;
		14439: rom = 1'b0;
		14440: rom = 1'b0;
		14441: rom = 1'b0;
		14442: rom = 1'b0;
		14443: rom = 1'b0;
		14444: rom = 1'b0;
		14445: rom = 1'b0;
		14446: rom = 1'b0;
		14447: rom = 1'b0;
		14448: rom = 1'b0;
		14449: rom = 1'b0;
		14450: rom = 1'b0;
		14451: rom = 1'b0;
		14452: rom = 1'b0;
		14453: rom = 1'b0;
		14454: rom = 1'b0;
		14455: rom = 1'b0;
		14456: rom = 1'b0;
		14457: rom = 1'b0;
		14458: rom = 1'b0;
		14459: rom = 1'b0;
		14460: rom = 1'b0;
		14461: rom = 1'b0;
		14462: rom = 1'b0;
		14463: rom = 1'b0;
		14464: rom = 1'b0;
		14465: rom = 1'b0;
		14466: rom = 1'b0;
		14467: rom = 1'b0;
		14468: rom = 1'b0;
		14469: rom = 1'b0;
		14470: rom = 1'b0;
		14471: rom = 1'b0;
		14472: rom = 1'b0;
		14473: rom = 1'b0;
		14474: rom = 1'b0;
		14475: rom = 1'b0;
		14476: rom = 1'b0;
		14477: rom = 1'b1;
		14478: rom = 1'b1;
		14479: rom = 1'b1;
		14480: rom = 1'b1;
		14481: rom = 1'b1;
		14482: rom = 1'b1;
		14483: rom = 1'b1;
		14484: rom = 1'b1;
		14485: rom = 1'b1;
		14486: rom = 1'b1;
		14487: rom = 1'b1;
		14488: rom = 1'b1;
		14489: rom = 1'b1;
		14490: rom = 1'b1;
		14491: rom = 1'b1;
		14492: rom = 1'b1;
		14493: rom = 1'b1;
		14494: rom = 1'b1;
		14495: rom = 1'b1;
		14496: rom = 1'b1;
		14497: rom = 1'b1;
		14498: rom = 1'b1;
		14499: rom = 1'b1;
		14500: rom = 1'b1;
		14501: rom = 1'b1;
		14502: rom = 1'b1;
		14503: rom = 1'b1;
		14504: rom = 1'b1;
		14505: rom = 1'b1;
		14506: rom = 1'b0;
		14507: rom = 1'b0;
		14508: rom = 1'b1;
		14509: rom = 1'b1;
		14510: rom = 1'b1;
		14511: rom = 1'b1;
		14512: rom = 1'b1;
		14513: rom = 1'b1;
		14514: rom = 1'b1;
		14515: rom = 1'b1;
		14516: rom = 1'b1;
		14517: rom = 1'b1;
		14518: rom = 1'b1;
		14519: rom = 1'b1;
		14520: rom = 1'b1;
		14521: rom = 1'b1;
		14522: rom = 1'b1;
		14523: rom = 1'b1;
		14524: rom = 1'b1;
		14525: rom = 1'b1;
		14526: rom = 1'b1;
		14527: rom = 1'b1;
		14528: rom = 1'b1;
		14529: rom = 1'b1;
		14530: rom = 1'b1;
		14531: rom = 1'b1;
		14532: rom = 1'b1;
		14533: rom = 1'b1;
		14534: rom = 1'b1;
		14535: rom = 1'b1;
		14536: rom = 1'b1;
		14537: rom = 1'b1;
		14538: rom = 1'b1;
		14539: rom = 1'b1;
		14540: rom = 1'b1;
		14541: rom = 1'b1;
		14542: rom = 1'b1;
		14543: rom = 1'b1;
		14544: rom = 1'b0;
		14545: rom = 1'b1;
		14546: rom = 1'b1;
		14547: rom = 1'b1;
		14548: rom = 1'b1;
		14549: rom = 1'b1;
		14550: rom = 1'b1;
		14551: rom = 1'b1;
		14552: rom = 1'b1;
		14553: rom = 1'b1;
		14554: rom = 1'b1;
		14555: rom = 1'b1;
		14556: rom = 1'b1;
		14557: rom = 1'b1;
		14558: rom = 1'b0;
		14559: rom = 1'b0;
		14560: rom = 1'b0;
		14561: rom = 1'b0;
		14562: rom = 1'b0;
		14563: rom = 1'b0;
		14564: rom = 1'b0;
		14565: rom = 1'b0;
		14566: rom = 1'b0;
		14567: rom = 1'b0;
		14568: rom = 1'b0;
		14569: rom = 1'b0;
		14570: rom = 1'b0;
		14571: rom = 1'b0;
		14572: rom = 1'b0;
		14573: rom = 1'b0;
		14574: rom = 1'b0;
		14575: rom = 1'b0;
		14576: rom = 1'b0;
		14577: rom = 1'b0;
		14578: rom = 1'b0;
		14579: rom = 1'b0;
		14580: rom = 1'b0;
		14581: rom = 1'b0;
		14582: rom = 1'b0;
		14583: rom = 1'b0;
		14584: rom = 1'b0;
		14585: rom = 1'b0;
		14586: rom = 1'b0;
		14587: rom = 1'b0;
		14588: rom = 1'b0;
		14589: rom = 1'b0;
		14590: rom = 1'b0;
		14591: rom = 1'b0;
		14592: rom = 1'b0;
		14593: rom = 1'b0;
		14594: rom = 1'b0;
		14595: rom = 1'b0;
		14596: rom = 1'b0;
		14597: rom = 1'b0;
		14598: rom = 1'b0;
		14599: rom = 1'b0;
		14600: rom = 1'b0;
		14601: rom = 1'b0;
		14602: rom = 1'b0;
		14603: rom = 1'b0;
		14604: rom = 1'b1;
		14605: rom = 1'b1;
		14606: rom = 1'b1;
		14607: rom = 1'b1;
		14608: rom = 1'b1;
		14609: rom = 1'b1;
		14610: rom = 1'b1;
		14611: rom = 1'b1;
		14612: rom = 1'b1;
		14613: rom = 1'b1;
		14614: rom = 1'b1;
		14615: rom = 1'b1;
		14616: rom = 1'b1;
		14617: rom = 1'b1;
		14618: rom = 1'b1;
		14619: rom = 1'b1;
		14620: rom = 1'b1;
		14621: rom = 1'b1;
		14622: rom = 1'b1;
		14623: rom = 1'b1;
		14624: rom = 1'b1;
		14625: rom = 1'b1;
		14626: rom = 1'b1;
		14627: rom = 1'b1;
		14628: rom = 1'b1;
		14629: rom = 1'b1;
		14630: rom = 1'b1;
		14631: rom = 1'b1;
		14632: rom = 1'b1;
		14633: rom = 1'b1;
		14634: rom = 1'b0;
		14635: rom = 1'b1;
		14636: rom = 1'b1;
		14637: rom = 1'b1;
		14638: rom = 1'b1;
		14639: rom = 1'b1;
		14640: rom = 1'b1;
		14641: rom = 1'b1;
		14642: rom = 1'b1;
		14643: rom = 1'b1;
		14644: rom = 1'b1;
		14645: rom = 1'b1;
		14646: rom = 1'b1;
		14647: rom = 1'b1;
		14648: rom = 1'b1;
		14649: rom = 1'b1;
		14650: rom = 1'b1;
		14651: rom = 1'b1;
		14652: rom = 1'b1;
		14653: rom = 1'b1;
		14654: rom = 1'b1;
		14655: rom = 1'b1;
		14656: rom = 1'b1;
		14657: rom = 1'b1;
		14658: rom = 1'b1;
		14659: rom = 1'b1;
		14660: rom = 1'b1;
		14661: rom = 1'b1;
		14662: rom = 1'b1;
		14663: rom = 1'b1;
		14664: rom = 1'b1;
		14665: rom = 1'b1;
		14666: rom = 1'b1;
		14667: rom = 1'b1;
		14668: rom = 1'b1;
		14669: rom = 1'b1;
		14670: rom = 1'b1;
		14671: rom = 1'b1;
		14672: rom = 1'b0;
		14673: rom = 1'b1;
		14674: rom = 1'b1;
		14675: rom = 1'b1;
		14676: rom = 1'b1;
		14677: rom = 1'b1;
		14678: rom = 1'b1;
		14679: rom = 1'b1;
		14680: rom = 1'b1;
		14681: rom = 1'b1;
		14682: rom = 1'b1;
		14683: rom = 1'b1;
		14684: rom = 1'b1;
		14685: rom = 1'b0;
		14686: rom = 1'b0;
		14687: rom = 1'b0;
		14688: rom = 1'b0;
		14689: rom = 1'b0;
		14690: rom = 1'b0;
		14691: rom = 1'b0;
		14692: rom = 1'b0;
		14693: rom = 1'b0;
		14694: rom = 1'b0;
		14695: rom = 1'b0;
		14696: rom = 1'b0;
		14697: rom = 1'b0;
		14698: rom = 1'b0;
		14699: rom = 1'b0;
		14700: rom = 1'b0;
		14701: rom = 1'b0;
		14702: rom = 1'b0;
		14703: rom = 1'b0;
		14704: rom = 1'b0;
		14705: rom = 1'b0;
		14706: rom = 1'b0;
		14707: rom = 1'b0;
		14708: rom = 1'b0;
		14709: rom = 1'b0;
		14710: rom = 1'b0;
		14711: rom = 1'b0;
		14712: rom = 1'b0;
		14713: rom = 1'b0;
		14714: rom = 1'b0;
		14715: rom = 1'b0;
		14716: rom = 1'b0;
		14717: rom = 1'b0;
		14718: rom = 1'b0;
		14719: rom = 1'b0;
		14720: rom = 1'b0;
		14721: rom = 1'b0;
		14722: rom = 1'b0;
		14723: rom = 1'b0;
		14724: rom = 1'b0;
		14725: rom = 1'b0;
		14726: rom = 1'b0;
		14727: rom = 1'b0;
		14728: rom = 1'b0;
		14729: rom = 1'b0;
		14730: rom = 1'b0;
		14731: rom = 1'b1;
		14732: rom = 1'b1;
		14733: rom = 1'b1;
		14734: rom = 1'b1;
		14735: rom = 1'b1;
		14736: rom = 1'b1;
		14737: rom = 1'b1;
		14738: rom = 1'b1;
		14739: rom = 1'b1;
		14740: rom = 1'b1;
		14741: rom = 1'b1;
		14742: rom = 1'b1;
		14743: rom = 1'b1;
		14744: rom = 1'b1;
		14745: rom = 1'b1;
		14746: rom = 1'b1;
		14747: rom = 1'b1;
		14748: rom = 1'b1;
		14749: rom = 1'b1;
		14750: rom = 1'b1;
		14751: rom = 1'b1;
		14752: rom = 1'b1;
		14753: rom = 1'b1;
		14754: rom = 1'b1;
		14755: rom = 1'b1;
		14756: rom = 1'b1;
		14757: rom = 1'b1;
		14758: rom = 1'b1;
		14759: rom = 1'b1;
		14760: rom = 1'b1;
		14761: rom = 1'b1;
		14762: rom = 1'b0;
		14763: rom = 1'b1;
		14764: rom = 1'b1;
		14765: rom = 1'b1;
		14766: rom = 1'b1;
		14767: rom = 1'b1;
		14768: rom = 1'b1;
		14769: rom = 1'b1;
		14770: rom = 1'b1;
		14771: rom = 1'b1;
		14772: rom = 1'b1;
		14773: rom = 1'b1;
		14774: rom = 1'b1;
		14775: rom = 1'b1;
		14776: rom = 1'b1;
		14777: rom = 1'b1;
		14778: rom = 1'b1;
		14779: rom = 1'b1;
		14780: rom = 1'b1;
		14781: rom = 1'b1;
		14782: rom = 1'b1;
		14783: rom = 1'b1;
		14784: rom = 1'b1;
		14785: rom = 1'b1;
		14786: rom = 1'b1;
		14787: rom = 1'b1;
		14788: rom = 1'b1;
		14789: rom = 1'b1;
		14790: rom = 1'b1;
		14791: rom = 1'b1;
		14792: rom = 1'b1;
		14793: rom = 1'b1;
		14794: rom = 1'b1;
		14795: rom = 1'b1;
		14796: rom = 1'b1;
		14797: rom = 1'b1;
		14798: rom = 1'b1;
		14799: rom = 1'b1;
		14800: rom = 1'b0;
		14801: rom = 1'b1;
		14802: rom = 1'b1;
		14803: rom = 1'b1;
		14804: rom = 1'b1;
		14805: rom = 1'b1;
		14806: rom = 1'b1;
		14807: rom = 1'b1;
		14808: rom = 1'b1;
		14809: rom = 1'b1;
		14810: rom = 1'b1;
		14811: rom = 1'b1;
		14812: rom = 1'b0;
		14813: rom = 1'b0;
		14814: rom = 1'b0;
		14815: rom = 1'b0;
		14816: rom = 1'b0;
		14817: rom = 1'b0;
		14818: rom = 1'b0;
		14819: rom = 1'b0;
		14820: rom = 1'b0;
		14821: rom = 1'b0;
		14822: rom = 1'b0;
		14823: rom = 1'b0;
		14824: rom = 1'b0;
		14825: rom = 1'b0;
		14826: rom = 1'b0;
		14827: rom = 1'b0;
		14828: rom = 1'b0;
		14829: rom = 1'b0;
		14830: rom = 1'b0;
		14831: rom = 1'b0;
		14832: rom = 1'b0;
		14833: rom = 1'b0;
		14834: rom = 1'b0;
		14835: rom = 1'b0;
		14836: rom = 1'b0;
		14837: rom = 1'b0;
		14838: rom = 1'b0;
		14839: rom = 1'b0;
		14840: rom = 1'b0;
		14841: rom = 1'b0;
		14842: rom = 1'b0;
		14843: rom = 1'b0;
		14844: rom = 1'b0;
		14845: rom = 1'b0;
		14846: rom = 1'b0;
		14847: rom = 1'b0;
		14848: rom = 1'b0;
		14849: rom = 1'b0;
		14850: rom = 1'b0;
		14851: rom = 1'b0;
		14852: rom = 1'b0;
		14853: rom = 1'b0;
		14854: rom = 1'b0;
		14855: rom = 1'b0;
		14856: rom = 1'b0;
		14857: rom = 1'b0;
		14858: rom = 1'b1;
		14859: rom = 1'b1;
		14860: rom = 1'b1;
		14861: rom = 1'b1;
		14862: rom = 1'b1;
		14863: rom = 1'b1;
		14864: rom = 1'b1;
		14865: rom = 1'b1;
		14866: rom = 1'b1;
		14867: rom = 1'b1;
		14868: rom = 1'b1;
		14869: rom = 1'b1;
		14870: rom = 1'b1;
		14871: rom = 1'b1;
		14872: rom = 1'b1;
		14873: rom = 1'b1;
		14874: rom = 1'b1;
		14875: rom = 1'b1;
		14876: rom = 1'b1;
		14877: rom = 1'b1;
		14878: rom = 1'b1;
		14879: rom = 1'b1;
		14880: rom = 1'b1;
		14881: rom = 1'b1;
		14882: rom = 1'b1;
		14883: rom = 1'b1;
		14884: rom = 1'b1;
		14885: rom = 1'b1;
		14886: rom = 1'b1;
		14887: rom = 1'b1;
		14888: rom = 1'b1;
		14889: rom = 1'b0;
		14890: rom = 1'b0;
		14891: rom = 1'b1;
		14892: rom = 1'b1;
		14893: rom = 1'b1;
		14894: rom = 1'b1;
		14895: rom = 1'b1;
		14896: rom = 1'b1;
		14897: rom = 1'b1;
		14898: rom = 1'b1;
		14899: rom = 1'b1;
		14900: rom = 1'b1;
		14901: rom = 1'b1;
		14902: rom = 1'b1;
		14903: rom = 1'b1;
		14904: rom = 1'b1;
		14905: rom = 1'b1;
		14906: rom = 1'b1;
		14907: rom = 1'b1;
		14908: rom = 1'b1;
		14909: rom = 1'b1;
		14910: rom = 1'b1;
		14911: rom = 1'b1;
		14912: rom = 1'b1;
		14913: rom = 1'b1;
		14914: rom = 1'b1;
		14915: rom = 1'b1;
		14916: rom = 1'b1;
		14917: rom = 1'b1;
		14918: rom = 1'b1;
		14919: rom = 1'b1;
		14920: rom = 1'b1;
		14921: rom = 1'b1;
		14922: rom = 1'b1;
		14923: rom = 1'b1;
		14924: rom = 1'b1;
		14925: rom = 1'b1;
		14926: rom = 1'b1;
		14927: rom = 1'b0;
		14928: rom = 1'b0;
		14929: rom = 1'b1;
		14930: rom = 1'b1;
		14931: rom = 1'b1;
		14932: rom = 1'b1;
		14933: rom = 1'b1;
		14934: rom = 1'b1;
		14935: rom = 1'b1;
		14936: rom = 1'b1;
		14937: rom = 1'b1;
		14938: rom = 1'b0;
		14939: rom = 1'b0;
		14940: rom = 1'b0;
		14941: rom = 1'b0;
		14942: rom = 1'b0;
		14943: rom = 1'b0;
		14944: rom = 1'b0;
		14945: rom = 1'b0;
		14946: rom = 1'b0;
		14947: rom = 1'b0;
		14948: rom = 1'b0;
		14949: rom = 1'b0;
		14950: rom = 1'b0;
		14951: rom = 1'b0;
		14952: rom = 1'b0;
		14953: rom = 1'b0;
		14954: rom = 1'b0;
		14955: rom = 1'b0;
		14956: rom = 1'b0;
		14957: rom = 1'b0;
		14958: rom = 1'b0;
		14959: rom = 1'b0;
		14960: rom = 1'b0;
		14961: rom = 1'b0;
		14962: rom = 1'b0;
		14963: rom = 1'b0;
		14964: rom = 1'b0;
		14965: rom = 1'b0;
		14966: rom = 1'b0;
		14967: rom = 1'b0;
		14968: rom = 1'b0;
		14969: rom = 1'b0;
		14970: rom = 1'b0;
		14971: rom = 1'b0;
		14972: rom = 1'b0;
		14973: rom = 1'b0;
		14974: rom = 1'b0;
		14975: rom = 1'b0;
		14976: rom = 1'b0;
		14977: rom = 1'b0;
		14978: rom = 1'b0;
		14979: rom = 1'b0;
		14980: rom = 1'b0;
		14981: rom = 1'b0;
		14982: rom = 1'b0;
		14983: rom = 1'b0;
		14984: rom = 1'b0;
		14985: rom = 1'b1;
		14986: rom = 1'b1;
		14987: rom = 1'b1;
		14988: rom = 1'b1;
		14989: rom = 1'b1;
		14990: rom = 1'b1;
		14991: rom = 1'b1;
		14992: rom = 1'b1;
		14993: rom = 1'b1;
		14994: rom = 1'b1;
		14995: rom = 1'b1;
		14996: rom = 1'b1;
		14997: rom = 1'b1;
		14998: rom = 1'b1;
		14999: rom = 1'b1;
		15000: rom = 1'b1;
		15001: rom = 1'b1;
		15002: rom = 1'b1;
		15003: rom = 1'b1;
		15004: rom = 1'b1;
		15005: rom = 1'b1;
		15006: rom = 1'b1;
		15007: rom = 1'b1;
		15008: rom = 1'b1;
		15009: rom = 1'b1;
		15010: rom = 1'b1;
		15011: rom = 1'b1;
		15012: rom = 1'b1;
		15013: rom = 1'b1;
		15014: rom = 1'b1;
		15015: rom = 1'b1;
		15016: rom = 1'b1;
		15017: rom = 1'b0;
		15018: rom = 1'b0;
		15019: rom = 1'b1;
		15020: rom = 1'b1;
		15021: rom = 1'b1;
		15022: rom = 1'b1;
		15023: rom = 1'b1;
		15024: rom = 1'b1;
		15025: rom = 1'b1;
		15026: rom = 1'b1;
		15027: rom = 1'b1;
		15028: rom = 1'b1;
		15029: rom = 1'b1;
		15030: rom = 1'b1;
		15031: rom = 1'b1;
		15032: rom = 1'b1;
		15033: rom = 1'b1;
		15034: rom = 1'b1;
		15035: rom = 1'b1;
		15036: rom = 1'b1;
		15037: rom = 1'b1;
		15038: rom = 1'b1;
		15039: rom = 1'b1;
		15040: rom = 1'b1;
		15041: rom = 1'b1;
		15042: rom = 1'b1;
		15043: rom = 1'b1;
		15044: rom = 1'b1;
		15045: rom = 1'b1;
		15046: rom = 1'b1;
		15047: rom = 1'b1;
		15048: rom = 1'b1;
		15049: rom = 1'b1;
		15050: rom = 1'b1;
		15051: rom = 1'b1;
		15052: rom = 1'b1;
		15053: rom = 1'b1;
		15054: rom = 1'b0;
		15055: rom = 1'b0;
		15056: rom = 1'b1;
		15057: rom = 1'b1;
		15058: rom = 1'b1;
		15059: rom = 1'b1;
		15060: rom = 1'b1;
		15061: rom = 1'b1;
		15062: rom = 1'b1;
		15063: rom = 1'b1;
		15064: rom = 1'b1;
		15065: rom = 1'b0;
		15066: rom = 1'b0;
		15067: rom = 1'b0;
		15068: rom = 1'b0;
		15069: rom = 1'b0;
		15070: rom = 1'b0;
		15071: rom = 1'b0;
		15072: rom = 1'b0;
		15073: rom = 1'b0;
		15074: rom = 1'b0;
		15075: rom = 1'b0;
		15076: rom = 1'b0;
		15077: rom = 1'b0;
		15078: rom = 1'b0;
		15079: rom = 1'b0;
		15080: rom = 1'b0;
		15081: rom = 1'b0;
		15082: rom = 1'b0;
		15083: rom = 1'b0;
		15084: rom = 1'b0;
		15085: rom = 1'b0;
		15086: rom = 1'b0;
		15087: rom = 1'b0;
		15088: rom = 1'b0;
		15089: rom = 1'b0;
		15090: rom = 1'b0;
		15091: rom = 1'b0;
		15092: rom = 1'b0;
		15093: rom = 1'b0;
		15094: rom = 1'b0;
		15095: rom = 1'b0;
		15096: rom = 1'b0;
		15097: rom = 1'b0;
		15098: rom = 1'b0;
		15099: rom = 1'b0;
		15100: rom = 1'b0;
		15101: rom = 1'b0;
		15102: rom = 1'b0;
		15103: rom = 1'b0;
		15104: rom = 1'b0;
		15105: rom = 1'b0;
		15106: rom = 1'b0;
		15107: rom = 1'b0;
		15108: rom = 1'b0;
		15109: rom = 1'b0;
		15110: rom = 1'b0;
		15111: rom = 1'b0;
		15112: rom = 1'b1;
		15113: rom = 1'b1;
		15114: rom = 1'b1;
		15115: rom = 1'b1;
		15116: rom = 1'b1;
		15117: rom = 1'b1;
		15118: rom = 1'b1;
		15119: rom = 1'b1;
		15120: rom = 1'b1;
		15121: rom = 1'b1;
		15122: rom = 1'b1;
		15123: rom = 1'b1;
		15124: rom = 1'b1;
		15125: rom = 1'b1;
		15126: rom = 1'b1;
		15127: rom = 1'b1;
		15128: rom = 1'b1;
		15129: rom = 1'b1;
		15130: rom = 1'b1;
		15131: rom = 1'b1;
		15132: rom = 1'b1;
		15133: rom = 1'b1;
		15134: rom = 1'b1;
		15135: rom = 1'b1;
		15136: rom = 1'b1;
		15137: rom = 1'b1;
		15138: rom = 1'b1;
		15139: rom = 1'b1;
		15140: rom = 1'b1;
		15141: rom = 1'b1;
		15142: rom = 1'b1;
		15143: rom = 1'b1;
		15144: rom = 1'b1;
		15145: rom = 1'b0;
		15146: rom = 1'b1;
		15147: rom = 1'b1;
		15148: rom = 1'b1;
		15149: rom = 1'b1;
		15150: rom = 1'b1;
		15151: rom = 1'b1;
		15152: rom = 1'b1;
		15153: rom = 1'b1;
		15154: rom = 1'b1;
		15155: rom = 1'b1;
		15156: rom = 1'b1;
		15157: rom = 1'b1;
		15158: rom = 1'b1;
		15159: rom = 1'b1;
		15160: rom = 1'b1;
		15161: rom = 1'b1;
		15162: rom = 1'b1;
		15163: rom = 1'b1;
		15164: rom = 1'b1;
		15165: rom = 1'b1;
		15166: rom = 1'b1;
		15167: rom = 1'b1;
		15168: rom = 1'b1;
		15169: rom = 1'b1;
		15170: rom = 1'b1;
		15171: rom = 1'b1;
		15172: rom = 1'b1;
		15173: rom = 1'b1;
		15174: rom = 1'b1;
		15175: rom = 1'b1;
		15176: rom = 1'b1;
		15177: rom = 1'b1;
		15178: rom = 1'b1;
		15179: rom = 1'b1;
		15180: rom = 1'b0;
		15181: rom = 1'b0;
		15182: rom = 1'b0;
		15183: rom = 1'b0;
		15184: rom = 1'b1;
		15185: rom = 1'b1;
		15186: rom = 1'b1;
		15187: rom = 1'b1;
		15188: rom = 1'b1;
		15189: rom = 1'b1;
		15190: rom = 1'b1;
		15191: rom = 1'b0;
		15192: rom = 1'b0;
		15193: rom = 1'b0;
		15194: rom = 1'b0;
		15195: rom = 1'b0;
		15196: rom = 1'b0;
		15197: rom = 1'b0;
		15198: rom = 1'b0;
		15199: rom = 1'b0;
		15200: rom = 1'b0;
		15201: rom = 1'b0;
		15202: rom = 1'b0;
		15203: rom = 1'b0;
		15204: rom = 1'b0;
		15205: rom = 1'b0;
		15206: rom = 1'b0;
		15207: rom = 1'b0;
		15208: rom = 1'b0;
		15209: rom = 1'b0;
		15210: rom = 1'b0;
		15211: rom = 1'b0;
		15212: rom = 1'b0;
		15213: rom = 1'b0;
		15214: rom = 1'b0;
		15215: rom = 1'b0;
		15216: rom = 1'b0;
		15217: rom = 1'b0;
		15218: rom = 1'b0;
		15219: rom = 1'b0;
		15220: rom = 1'b0;
		15221: rom = 1'b0;
		15222: rom = 1'b0;
		15223: rom = 1'b0;
		15224: rom = 1'b0;
		15225: rom = 1'b0;
		15226: rom = 1'b0;
		15227: rom = 1'b0;
		15228: rom = 1'b0;
		15229: rom = 1'b0;
		15230: rom = 1'b0;
		15231: rom = 1'b0;
		15232: rom = 1'b0;
		15233: rom = 1'b0;
		15234: rom = 1'b0;
		15235: rom = 1'b0;
		15236: rom = 1'b0;
		15237: rom = 1'b0;
		15238: rom = 1'b1;
		15239: rom = 1'b1;
		15240: rom = 1'b1;
		15241: rom = 1'b1;
		15242: rom = 1'b1;
		15243: rom = 1'b1;
		15244: rom = 1'b1;
		15245: rom = 1'b1;
		15246: rom = 1'b1;
		15247: rom = 1'b1;
		15248: rom = 1'b1;
		15249: rom = 1'b1;
		15250: rom = 1'b1;
		15251: rom = 1'b1;
		15252: rom = 1'b1;
		15253: rom = 1'b1;
		15254: rom = 1'b1;
		15255: rom = 1'b1;
		15256: rom = 1'b1;
		15257: rom = 1'b1;
		15258: rom = 1'b1;
		15259: rom = 1'b1;
		15260: rom = 1'b1;
		15261: rom = 1'b1;
		15262: rom = 1'b1;
		15263: rom = 1'b1;
		15264: rom = 1'b1;
		15265: rom = 1'b1;
		15266: rom = 1'b1;
		15267: rom = 1'b1;
		15268: rom = 1'b1;
		15269: rom = 1'b1;
		15270: rom = 1'b1;
		15271: rom = 1'b1;
		15272: rom = 1'b0;
		15273: rom = 1'b0;
		15274: rom = 1'b1;
		15275: rom = 1'b1;
		15276: rom = 1'b1;
		15277: rom = 1'b1;
		15278: rom = 1'b1;
		15279: rom = 1'b1;
		15280: rom = 1'b1;
		15281: rom = 1'b1;
		15282: rom = 1'b1;
		15283: rom = 1'b1;
		15284: rom = 1'b1;
		15285: rom = 1'b1;
		15286: rom = 1'b1;
		15287: rom = 1'b1;
		15288: rom = 1'b1;
		15289: rom = 1'b1;
		15290: rom = 1'b1;
		15291: rom = 1'b1;
		15292: rom = 1'b1;
		15293: rom = 1'b1;
		15294: rom = 1'b1;
		15295: rom = 1'b1;
		15296: rom = 1'b1;
		15297: rom = 1'b1;
		15298: rom = 1'b1;
		15299: rom = 1'b1;
		15300: rom = 1'b1;
		15301: rom = 1'b1;
		15302: rom = 1'b1;
		15303: rom = 1'b1;
		15304: rom = 1'b1;
		15305: rom = 1'b1;
		15306: rom = 1'b0;
		15307: rom = 1'b0;
		15308: rom = 1'b0;
		15309: rom = 1'b0;
		15310: rom = 1'b0;
		15311: rom = 1'b0;
		15312: rom = 1'b1;
		15313: rom = 1'b1;
		15314: rom = 1'b1;
		15315: rom = 1'b1;
		15316: rom = 1'b1;
		15317: rom = 1'b0;
		15318: rom = 1'b0;
		15319: rom = 1'b0;
		15320: rom = 1'b0;
		15321: rom = 1'b0;
		15322: rom = 1'b0;
		15323: rom = 1'b0;
		15324: rom = 1'b0;
		15325: rom = 1'b0;
		15326: rom = 1'b0;
		15327: rom = 1'b0;
		15328: rom = 1'b0;
		15329: rom = 1'b0;
		15330: rom = 1'b0;
		15331: rom = 1'b0;
		15332: rom = 1'b0;
		15333: rom = 1'b0;
		15334: rom = 1'b0;
		15335: rom = 1'b0;
		15336: rom = 1'b0;
		15337: rom = 1'b0;
		15338: rom = 1'b0;
		15339: rom = 1'b0;
		15340: rom = 1'b0;
		15341: rom = 1'b0;
		15342: rom = 1'b0;
		15343: rom = 1'b0;
		15344: rom = 1'b0;
		15345: rom = 1'b0;
		15346: rom = 1'b0;
		15347: rom = 1'b0;
		15348: rom = 1'b0;
		15349: rom = 1'b0;
		15350: rom = 1'b0;
		15351: rom = 1'b0;
		15352: rom = 1'b0;
		15353: rom = 1'b0;
		15354: rom = 1'b0;
		15355: rom = 1'b0;
		15356: rom = 1'b0;
		15357: rom = 1'b0;
		15358: rom = 1'b0;
		15359: rom = 1'b0;
		15360: rom = 1'b0;
		15361: rom = 1'b0;
		15362: rom = 1'b0;
		15363: rom = 1'b0;
		15364: rom = 1'b0;
		15365: rom = 1'b0;
		15366: rom = 1'b0;
		15367: rom = 1'b1;
		15368: rom = 1'b1;
		15369: rom = 1'b1;
		15370: rom = 1'b1;
		15371: rom = 1'b1;
		15372: rom = 1'b1;
		15373: rom = 1'b1;
		15374: rom = 1'b1;
		15375: rom = 1'b1;
		15376: rom = 1'b1;
		15377: rom = 1'b1;
		15378: rom = 1'b1;
		15379: rom = 1'b1;
		15380: rom = 1'b1;
		15381: rom = 1'b1;
		15382: rom = 1'b1;
		15383: rom = 1'b1;
		15384: rom = 1'b1;
		15385: rom = 1'b1;
		15386: rom = 1'b1;
		15387: rom = 1'b1;
		15388: rom = 1'b1;
		15389: rom = 1'b1;
		15390: rom = 1'b1;
		15391: rom = 1'b1;
		15392: rom = 1'b1;
		15393: rom = 1'b1;
		15394: rom = 1'b1;
		15395: rom = 1'b1;
		15396: rom = 1'b1;
		15397: rom = 1'b0;
		15398: rom = 1'b0;
		15399: rom = 1'b0;
		15400: rom = 1'b0;
		15401: rom = 1'b0;
		15402: rom = 1'b1;
		15403: rom = 1'b1;
		15404: rom = 1'b1;
		15405: rom = 1'b1;
		15406: rom = 1'b1;
		15407: rom = 1'b1;
		15408: rom = 1'b1;
		15409: rom = 1'b1;
		15410: rom = 1'b1;
		15411: rom = 1'b1;
		15412: rom = 1'b1;
		15413: rom = 1'b1;
		15414: rom = 1'b1;
		15415: rom = 1'b1;
		15416: rom = 1'b1;
		15417: rom = 1'b1;
		15418: rom = 1'b1;
		15419: rom = 1'b1;
		15420: rom = 1'b1;
		15421: rom = 1'b1;
		15422: rom = 1'b1;
		15423: rom = 1'b1;
		15424: rom = 1'b1;
		15425: rom = 1'b1;
		15426: rom = 1'b1;
		15427: rom = 1'b1;
		15428: rom = 1'b1;
		15429: rom = 1'b1;
		15430: rom = 1'b1;
		15431: rom = 1'b1;
		15432: rom = 1'b0;
		15433: rom = 1'b0;
		15434: rom = 1'b0;
		15435: rom = 1'b0;
		15436: rom = 1'b0;
		15437: rom = 1'b0;
		15438: rom = 1'b0;
		15439: rom = 1'b0;
		15440: rom = 1'b1;
		15441: rom = 1'b1;
		15442: rom = 1'b1;
		15443: rom = 1'b0;
		15444: rom = 1'b0;
		15445: rom = 1'b0;
		15446: rom = 1'b0;
		15447: rom = 1'b0;
		15448: rom = 1'b0;
		15449: rom = 1'b0;
		15450: rom = 1'b0;
		15451: rom = 1'b0;
		15452: rom = 1'b0;
		15453: rom = 1'b0;
		15454: rom = 1'b0;
		15455: rom = 1'b0;
		15456: rom = 1'b0;
		15457: rom = 1'b0;
		15458: rom = 1'b0;
		15459: rom = 1'b0;
		15460: rom = 1'b0;
		15461: rom = 1'b0;
		15462: rom = 1'b0;
		15463: rom = 1'b0;
		15464: rom = 1'b0;
		15465: rom = 1'b0;
		15466: rom = 1'b0;
		15467: rom = 1'b0;
		15468: rom = 1'b0;
		15469: rom = 1'b0;
		15470: rom = 1'b0;
		15471: rom = 1'b0;
		15472: rom = 1'b0;
		15473: rom = 1'b0;
		15474: rom = 1'b0;
		15475: rom = 1'b0;
		15476: rom = 1'b0;
		15477: rom = 1'b0;
		15478: rom = 1'b0;
		15479: rom = 1'b0;
		15480: rom = 1'b0;
		15481: rom = 1'b0;
		15482: rom = 1'b0;
		15483: rom = 1'b0;
		15484: rom = 1'b0;
		15485: rom = 1'b0;
		15486: rom = 1'b0;
		15487: rom = 1'b0;
		15488: rom = 1'b0;
		15489: rom = 1'b0;
		15490: rom = 1'b0;
		15491: rom = 1'b0;
		15492: rom = 1'b0;
		15493: rom = 1'b0;
		15494: rom = 1'b0;
		15495: rom = 1'b0;
		15496: rom = 1'b0;
		15497: rom = 1'b0;
		15498: rom = 1'b0;
		15499: rom = 1'b0;
		15500: rom = 1'b0;
		15501: rom = 1'b0;
		15502: rom = 1'b1;
		15503: rom = 1'b1;
		15504: rom = 1'b1;
		15505: rom = 1'b1;
		15506: rom = 1'b1;
		15507: rom = 1'b1;
		15508: rom = 1'b1;
		15509: rom = 1'b1;
		15510: rom = 1'b1;
		15511: rom = 1'b1;
		15512: rom = 1'b1;
		15513: rom = 1'b1;
		15514: rom = 1'b1;
		15515: rom = 1'b1;
		15516: rom = 1'b1;
		15517: rom = 1'b1;
		15518: rom = 1'b1;
		15519: rom = 1'b0;
		15520: rom = 1'b0;
		15521: rom = 1'b0;
		15522: rom = 1'b0;
		15523: rom = 1'b0;
		15524: rom = 1'b0;
		15525: rom = 1'b0;
		15526: rom = 1'b0;
		15527: rom = 1'b0;
		15528: rom = 1'b0;
		15529: rom = 1'b0;
		15530: rom = 1'b1;
		15531: rom = 1'b1;
		15532: rom = 1'b1;
		15533: rom = 1'b1;
		15534: rom = 1'b1;
		15535: rom = 1'b1;
		15536: rom = 1'b1;
		15537: rom = 1'b1;
		15538: rom = 1'b1;
		15539: rom = 1'b1;
		15540: rom = 1'b1;
		15541: rom = 1'b1;
		15542: rom = 1'b1;
		15543: rom = 1'b1;
		15544: rom = 1'b1;
		15545: rom = 1'b1;
		15546: rom = 1'b1;
		15547: rom = 1'b1;
		15548: rom = 1'b1;
		15549: rom = 1'b1;
		15550: rom = 1'b1;
		15551: rom = 1'b1;
		15552: rom = 1'b1;
		15553: rom = 1'b1;
		15554: rom = 1'b1;
		15555: rom = 1'b1;
		15556: rom = 1'b1;
		15557: rom = 1'b1;
		15558: rom = 1'b0;
		15559: rom = 1'b0;
		15560: rom = 1'b0;
		15561: rom = 1'b0;
		15562: rom = 1'b0;
		15563: rom = 1'b0;
		15564: rom = 1'b0;
		15565: rom = 1'b0;
		15566: rom = 1'b0;
		15567: rom = 1'b1;
		15568: rom = 1'b1;
		15569: rom = 1'b0;
		15570: rom = 1'b0;
		15571: rom = 1'b0;
		15572: rom = 1'b0;
		15573: rom = 1'b0;
		15574: rom = 1'b0;
		15575: rom = 1'b0;
		15576: rom = 1'b0;
		15577: rom = 1'b0;
		15578: rom = 1'b0;
		15579: rom = 1'b0;
		15580: rom = 1'b0;
		15581: rom = 1'b0;
		15582: rom = 1'b0;
		15583: rom = 1'b0;
		15584: rom = 1'b0;
		15585: rom = 1'b0;
		15586: rom = 1'b0;
		15587: rom = 1'b0;
		15588: rom = 1'b0;
		15589: rom = 1'b0;
		15590: rom = 1'b0;
		15591: rom = 1'b0;
		15592: rom = 1'b0;
		15593: rom = 1'b0;
		15594: rom = 1'b0;
		15595: rom = 1'b0;
		15596: rom = 1'b0;
		15597: rom = 1'b0;
		15598: rom = 1'b0;
		15599: rom = 1'b0;
		15600: rom = 1'b0;
		15601: rom = 1'b0;
		15602: rom = 1'b0;
		15603: rom = 1'b0;
		15604: rom = 1'b0;
		15605: rom = 1'b0;
		15606: rom = 1'b0;
		15607: rom = 1'b0;
		15608: rom = 1'b0;
		15609: rom = 1'b0;
		15610: rom = 1'b0;
		15611: rom = 1'b0;
		15612: rom = 1'b0;
		15613: rom = 1'b0;
		15614: rom = 1'b0;
		15615: rom = 1'b0;
		15616: rom = 1'b0;
		15617: rom = 1'b0;
		15618: rom = 1'b0;
		15619: rom = 1'b0;
		15620: rom = 1'b0;
		15621: rom = 1'b0;
		15622: rom = 1'b0;
		15623: rom = 1'b0;
		15624: rom = 1'b0;
		15625: rom = 1'b0;
		15626: rom = 1'b0;
		15627: rom = 1'b0;
		15628: rom = 1'b0;
		15629: rom = 1'b0;
		15630: rom = 1'b0;
		15631: rom = 1'b0;
		15632: rom = 1'b0;
		15633: rom = 1'b0;
		15634: rom = 1'b0;
		15635: rom = 1'b0;
		15636: rom = 1'b0;
		15637: rom = 1'b0;
		15638: rom = 1'b0;
		15639: rom = 1'b0;
		15640: rom = 1'b0;
		15641: rom = 1'b0;
		15642: rom = 1'b0;
		15643: rom = 1'b0;
		15644: rom = 1'b0;
		15645: rom = 1'b0;
		15646: rom = 1'b0;
		15647: rom = 1'b0;
		15648: rom = 1'b0;
		15649: rom = 1'b0;
		15650: rom = 1'b0;
		15651: rom = 1'b0;
		15652: rom = 1'b0;
		15653: rom = 1'b0;
		15654: rom = 1'b0;
		15655: rom = 1'b0;
		15656: rom = 1'b0;
		15657: rom = 1'b1;
		15658: rom = 1'b1;
		15659: rom = 1'b1;
		15660: rom = 1'b1;
		15661: rom = 1'b1;
		15662: rom = 1'b1;
		15663: rom = 1'b1;
		15664: rom = 1'b1;
		15665: rom = 1'b1;
		15666: rom = 1'b1;
		15667: rom = 1'b1;
		15668: rom = 1'b1;
		15669: rom = 1'b1;
		15670: rom = 1'b1;
		15671: rom = 1'b1;
		15672: rom = 1'b1;
		15673: rom = 1'b1;
		15674: rom = 1'b1;
		15675: rom = 1'b1;
		15676: rom = 1'b1;
		15677: rom = 1'b1;
		15678: rom = 1'b1;
		15679: rom = 1'b1;
		15680: rom = 1'b1;
		15681: rom = 1'b1;
		15682: rom = 1'b1;
		15683: rom = 1'b0;
		15684: rom = 1'b0;
		15685: rom = 1'b0;
		15686: rom = 1'b0;
		15687: rom = 1'b0;
		15688: rom = 1'b0;
		15689: rom = 1'b0;
		15690: rom = 1'b0;
		15691: rom = 1'b0;
		15692: rom = 1'b0;
		15693: rom = 1'b0;
		15694: rom = 1'b0;
		15695: rom = 1'b0;
		15696: rom = 1'b0;
		15697: rom = 1'b0;
		15698: rom = 1'b0;
		15699: rom = 1'b0;
		15700: rom = 1'b0;
		15701: rom = 1'b0;
		15702: rom = 1'b0;
		15703: rom = 1'b0;
		15704: rom = 1'b0;
		15705: rom = 1'b0;
		15706: rom = 1'b0;
		15707: rom = 1'b0;
		15708: rom = 1'b0;
		15709: rom = 1'b0;
		15710: rom = 1'b0;
		15711: rom = 1'b0;
		15712: rom = 1'b0;
		15713: rom = 1'b0;
		15714: rom = 1'b0;
		15715: rom = 1'b0;
		15716: rom = 1'b0;
		15717: rom = 1'b0;
		15718: rom = 1'b0;
		15719: rom = 1'b0;
		15720: rom = 1'b0;
		15721: rom = 1'b0;
		15722: rom = 1'b0;
		15723: rom = 1'b0;
		15724: rom = 1'b0;
		15725: rom = 1'b0;
		15726: rom = 1'b0;
		15727: rom = 1'b0;
		15728: rom = 1'b0;
		15729: rom = 1'b0;
		15730: rom = 1'b0;
		15731: rom = 1'b0;
		15732: rom = 1'b0;
		15733: rom = 1'b0;
		15734: rom = 1'b0;
		15735: rom = 1'b0;
		15736: rom = 1'b0;
		15737: rom = 1'b0;
		15738: rom = 1'b0;
		15739: rom = 1'b0;
		15740: rom = 1'b0;
		15741: rom = 1'b0;
		15742: rom = 1'b0;
		15743: rom = 1'b0;
		15744: rom = 1'b0;
		15745: rom = 1'b0;
		15746: rom = 1'b0;
		15747: rom = 1'b0;
		15748: rom = 1'b0;
		15749: rom = 1'b0;
		15750: rom = 1'b0;
		15751: rom = 1'b0;
		15752: rom = 1'b0;
		15753: rom = 1'b0;
		15754: rom = 1'b0;
		15755: rom = 1'b0;
		15756: rom = 1'b0;
		15757: rom = 1'b0;
		15758: rom = 1'b0;
		15759: rom = 1'b0;
		15760: rom = 1'b0;
		15761: rom = 1'b0;
		15762: rom = 1'b0;
		15763: rom = 1'b0;
		15764: rom = 1'b0;
		15765: rom = 1'b0;
		15766: rom = 1'b0;
		15767: rom = 1'b0;
		15768: rom = 1'b0;
		15769: rom = 1'b0;
		15770: rom = 1'b0;
		15771: rom = 1'b0;
		15772: rom = 1'b0;
		15773: rom = 1'b0;
		15774: rom = 1'b0;
		15775: rom = 1'b0;
		15776: rom = 1'b0;
		15777: rom = 1'b0;
		15778: rom = 1'b0;
		15779: rom = 1'b0;
		15780: rom = 1'b0;
		15781: rom = 1'b0;
		15782: rom = 1'b0;
		15783: rom = 1'b0;
		15784: rom = 1'b1;
		15785: rom = 1'b1;
		15786: rom = 1'b1;
		15787: rom = 1'b1;
		15788: rom = 1'b1;
		15789: rom = 1'b1;
		15790: rom = 1'b1;
		15791: rom = 1'b1;
		15792: rom = 1'b1;
		15793: rom = 1'b1;
		15794: rom = 1'b1;
		15795: rom = 1'b1;
		15796: rom = 1'b1;
		15797: rom = 1'b1;
		15798: rom = 1'b1;
		15799: rom = 1'b1;
		15800: rom = 1'b1;
		15801: rom = 1'b1;
		15802: rom = 1'b1;
		15803: rom = 1'b1;
		15804: rom = 1'b1;
		15805: rom = 1'b1;
		15806: rom = 1'b1;
		15807: rom = 1'b1;
		15808: rom = 1'b0;
		15809: rom = 1'b0;
		15810: rom = 1'b0;
		15811: rom = 1'b0;
		15812: rom = 1'b0;
		15813: rom = 1'b0;
		15814: rom = 1'b0;
		15815: rom = 1'b0;
		15816: rom = 1'b0;
		15817: rom = 1'b0;
		15818: rom = 1'b0;
		15819: rom = 1'b0;
		15820: rom = 1'b0;
		15821: rom = 1'b0;
		15822: rom = 1'b0;
		15823: rom = 1'b0;
		15824: rom = 1'b0;
		15825: rom = 1'b0;
		15826: rom = 1'b0;
		15827: rom = 1'b0;
		15828: rom = 1'b0;
		15829: rom = 1'b0;
		15830: rom = 1'b0;
		15831: rom = 1'b0;
		15832: rom = 1'b0;
		15833: rom = 1'b0;
		15834: rom = 1'b0;
		15835: rom = 1'b0;
		15836: rom = 1'b0;
		15837: rom = 1'b0;
		15838: rom = 1'b0;
		15839: rom = 1'b0;
		15840: rom = 1'b0;
		15841: rom = 1'b0;
		15842: rom = 1'b0;
		15843: rom = 1'b0;
		15844: rom = 1'b0;
		15845: rom = 1'b0;
		15846: rom = 1'b0;
		15847: rom = 1'b0;
		15848: rom = 1'b0;
		15849: rom = 1'b0;
		15850: rom = 1'b0;
		15851: rom = 1'b0;
		15852: rom = 1'b0;
		15853: rom = 1'b0;
		15854: rom = 1'b0;
		15855: rom = 1'b0;
		15856: rom = 1'b0;
		15857: rom = 1'b0;
		15858: rom = 1'b0;
		15859: rom = 1'b0;
		15860: rom = 1'b0;
		15861: rom = 1'b0;
		15862: rom = 1'b0;
		15863: rom = 1'b0;
		15864: rom = 1'b0;
		15865: rom = 1'b0;
		15866: rom = 1'b0;
		15867: rom = 1'b0;
		15868: rom = 1'b0;
		15869: rom = 1'b0;
		15870: rom = 1'b0;
		15871: rom = 1'b0;
		15872: rom = 1'b0;
		15873: rom = 1'b0;
		15874: rom = 1'b0;
		15875: rom = 1'b0;
		15876: rom = 1'b0;
		15877: rom = 1'b0;
		15878: rom = 1'b0;
		15879: rom = 1'b0;
		15880: rom = 1'b0;
		15881: rom = 1'b0;
		15882: rom = 1'b0;
		15883: rom = 1'b0;
		15884: rom = 1'b0;
		15885: rom = 1'b0;
		15886: rom = 1'b0;
		15887: rom = 1'b0;
		15888: rom = 1'b0;
		15889: rom = 1'b0;
		15890: rom = 1'b0;
		15891: rom = 1'b0;
		15892: rom = 1'b0;
		15893: rom = 1'b0;
		15894: rom = 1'b0;
		15895: rom = 1'b0;
		15896: rom = 1'b0;
		15897: rom = 1'b0;
		15898: rom = 1'b0;
		15899: rom = 1'b0;
		15900: rom = 1'b0;
		15901: rom = 1'b0;
		15902: rom = 1'b0;
		15903: rom = 1'b0;
		15904: rom = 1'b0;
		15905: rom = 1'b0;
		15906: rom = 1'b0;
		15907: rom = 1'b0;
		15908: rom = 1'b0;
		15909: rom = 1'b0;
		15910: rom = 1'b0;
		15911: rom = 1'b0;
		15912: rom = 1'b1;
		15913: rom = 1'b1;
		15914: rom = 1'b1;
		15915: rom = 1'b1;
		15916: rom = 1'b1;
		15917: rom = 1'b1;
		15918: rom = 1'b1;
		15919: rom = 1'b1;
		15920: rom = 1'b1;
		15921: rom = 1'b1;
		15922: rom = 1'b1;
		15923: rom = 1'b1;
		15924: rom = 1'b1;
		15925: rom = 1'b1;
		15926: rom = 1'b1;
		15927: rom = 1'b1;
		15928: rom = 1'b1;
		15929: rom = 1'b1;
		15930: rom = 1'b1;
		15931: rom = 1'b0;
		15932: rom = 1'b0;
		15933: rom = 1'b0;
		15934: rom = 1'b0;
		15935: rom = 1'b0;
		15936: rom = 1'b0;
		15937: rom = 1'b0;
		15938: rom = 1'b0;
		15939: rom = 1'b0;
		15940: rom = 1'b0;
		15941: rom = 1'b0;
		15942: rom = 1'b0;
		15943: rom = 1'b0;
		15944: rom = 1'b0;
		15945: rom = 1'b0;
		15946: rom = 1'b0;
		15947: rom = 1'b0;
		15948: rom = 1'b0;
		15949: rom = 1'b0;
		15950: rom = 1'b0;
		15951: rom = 1'b0;
		15952: rom = 1'b0;
		15953: rom = 1'b0;
		15954: rom = 1'b0;
		15955: rom = 1'b0;
		15956: rom = 1'b0;
		15957: rom = 1'b0;
		15958: rom = 1'b0;
		15959: rom = 1'b0;
		15960: rom = 1'b0;
		15961: rom = 1'b0;
		15962: rom = 1'b0;
		15963: rom = 1'b0;
		15964: rom = 1'b0;
		15965: rom = 1'b0;
		15966: rom = 1'b0;
		15967: rom = 1'b0;
		15968: rom = 1'b0;
		15969: rom = 1'b0;
		15970: rom = 1'b0;
		15971: rom = 1'b0;
		15972: rom = 1'b0;
		15973: rom = 1'b0;
		15974: rom = 1'b0;
		15975: rom = 1'b0;
		15976: rom = 1'b0;
		15977: rom = 1'b0;
		15978: rom = 1'b0;
		15979: rom = 1'b0;
		15980: rom = 1'b0;
		15981: rom = 1'b0;
		15982: rom = 1'b0;
		15983: rom = 1'b0;
		15984: rom = 1'b0;
		15985: rom = 1'b0;
		15986: rom = 1'b0;
		15987: rom = 1'b0;
		15988: rom = 1'b0;
		15989: rom = 1'b0;
		15990: rom = 1'b0;
		15991: rom = 1'b0;
		15992: rom = 1'b0;
		15993: rom = 1'b0;
		15994: rom = 1'b0;
		15995: rom = 1'b0;
		15996: rom = 1'b0;
		15997: rom = 1'b0;
		15998: rom = 1'b0;
		15999: rom = 1'b0;
		16000: rom = 1'b0;
		16001: rom = 1'b0;
		16002: rom = 1'b0;
		16003: rom = 1'b0;
		16004: rom = 1'b0;
		16005: rom = 1'b0;
		16006: rom = 1'b0;
		16007: rom = 1'b0;
		16008: rom = 1'b0;
		16009: rom = 1'b0;
		16010: rom = 1'b0;
		16011: rom = 1'b0;
		16012: rom = 1'b0;
		16013: rom = 1'b0;
		16014: rom = 1'b0;
		16015: rom = 1'b0;
		16016: rom = 1'b0;
		16017: rom = 1'b0;
		16018: rom = 1'b0;
		16019: rom = 1'b0;
		16020: rom = 1'b0;
		16021: rom = 1'b0;
		16022: rom = 1'b0;
		16023: rom = 1'b0;
		16024: rom = 1'b0;
		16025: rom = 1'b0;
		16026: rom = 1'b0;
		16027: rom = 1'b0;
		16028: rom = 1'b0;
		16029: rom = 1'b0;
		16030: rom = 1'b0;
		16031: rom = 1'b0;
		16032: rom = 1'b0;
		16033: rom = 1'b0;
		16034: rom = 1'b0;
		16035: rom = 1'b0;
		16036: rom = 1'b0;
		16037: rom = 1'b0;
		16038: rom = 1'b0;
		16039: rom = 1'b0;
		16040: rom = 1'b0;
		16041: rom = 1'b1;
		16042: rom = 1'b1;
		16043: rom = 1'b1;
		16044: rom = 1'b1;
		16045: rom = 1'b1;
		16046: rom = 1'b1;
		16047: rom = 1'b1;
		16048: rom = 1'b0;
		16049: rom = 1'b0;
		16050: rom = 1'b0;
		16051: rom = 1'b0;
		16052: rom = 1'b0;
		16053: rom = 1'b0;
		16054: rom = 1'b0;
		16055: rom = 1'b0;
		16056: rom = 1'b0;
		16057: rom = 1'b0;
		16058: rom = 1'b0;
		16059: rom = 1'b0;
		16060: rom = 1'b0;
		16061: rom = 1'b0;
		16062: rom = 1'b0;
		16063: rom = 1'b0;
		16064: rom = 1'b0;
		16065: rom = 1'b0;
		16066: rom = 1'b0;
		16067: rom = 1'b0;
		16068: rom = 1'b0;
		16069: rom = 1'b0;
		16070: rom = 1'b0;
		16071: rom = 1'b0;
		16072: rom = 1'b0;
		16073: rom = 1'b0;
		16074: rom = 1'b0;
		16075: rom = 1'b0;
		16076: rom = 1'b0;
		16077: rom = 1'b0;
		16078: rom = 1'b0;
		16079: rom = 1'b0;
		16080: rom = 1'b0;
		16081: rom = 1'b0;
		16082: rom = 1'b0;
		16083: rom = 1'b0;
		16084: rom = 1'b0;
		16085: rom = 1'b0;
		16086: rom = 1'b0;
		16087: rom = 1'b0;
		16088: rom = 1'b0;
		16089: rom = 1'b0;
		16090: rom = 1'b0;
		16091: rom = 1'b0;
		16092: rom = 1'b0;
		16093: rom = 1'b0;
		16094: rom = 1'b0;
		16095: rom = 1'b0;
		16096: rom = 1'b0;
		16097: rom = 1'b0;
		16098: rom = 1'b0;
		16099: rom = 1'b0;
		16100: rom = 1'b0;
		16101: rom = 1'b0;
		16102: rom = 1'b0;
		16103: rom = 1'b0;
		16104: rom = 1'b0;
		16105: rom = 1'b0;
		16106: rom = 1'b0;
		16107: rom = 1'b0;
		16108: rom = 1'b0;
		16109: rom = 1'b0;
		16110: rom = 1'b0;
		16111: rom = 1'b0;
		16112: rom = 1'b0;
		16113: rom = 1'b0;
		16114: rom = 1'b0;
		16115: rom = 1'b0;
		16116: rom = 1'b0;
		16117: rom = 1'b0;
		16118: rom = 1'b0;
		16119: rom = 1'b0;
		16120: rom = 1'b0;
		16121: rom = 1'b0;
		16122: rom = 1'b0;
		16123: rom = 1'b0;
		16124: rom = 1'b0;
		16125: rom = 1'b0;
		16126: rom = 1'b0;
		16127: rom = 1'b0;
		16128: rom = 1'b0;
		16129: rom = 1'b0;
		16130: rom = 1'b0;
		16131: rom = 1'b0;
		16132: rom = 1'b0;
		16133: rom = 1'b0;
		16134: rom = 1'b0;
		16135: rom = 1'b0;
		16136: rom = 1'b0;
		16137: rom = 1'b0;
		16138: rom = 1'b0;
		16139: rom = 1'b0;
		16140: rom = 1'b0;
		16141: rom = 1'b0;
		16142: rom = 1'b0;
		16143: rom = 1'b0;
		16144: rom = 1'b0;
		16145: rom = 1'b0;
		16146: rom = 1'b0;
		16147: rom = 1'b0;
		16148: rom = 1'b0;
		16149: rom = 1'b0;
		16150: rom = 1'b0;
		16151: rom = 1'b0;
		16152: rom = 1'b0;
		16153: rom = 1'b0;
		16154: rom = 1'b0;
		16155: rom = 1'b0;
		16156: rom = 1'b0;
		16157: rom = 1'b0;
		16158: rom = 1'b0;
		16159: rom = 1'b0;
		16160: rom = 1'b0;
		16161: rom = 1'b0;
		16162: rom = 1'b0;
		16163: rom = 1'b0;
		16164: rom = 1'b0;
		16165: rom = 1'b0;
		16166: rom = 1'b0;
		16167: rom = 1'b0;
		16168: rom = 1'b0;
		16169: rom = 1'b0;
		16170: rom = 1'b0;
		16171: rom = 1'b0;
		16172: rom = 1'b0;
		16173: rom = 1'b0;
		16174: rom = 1'b0;
		16175: rom = 1'b0;
		16176: rom = 1'b0;
		16177: rom = 1'b0;
		16178: rom = 1'b0;
		16179: rom = 1'b0;
		16180: rom = 1'b0;
		16181: rom = 1'b0;
		16182: rom = 1'b0;
		16183: rom = 1'b0;
		16184: rom = 1'b0;
		16185: rom = 1'b0;
		16186: rom = 1'b0;
		16187: rom = 1'b0;
		16188: rom = 1'b0;
		16189: rom = 1'b0;
		16190: rom = 1'b0;
		16191: rom = 1'b0;
		16192: rom = 1'b0;
		16193: rom = 1'b0;
		16194: rom = 1'b0;
		16195: rom = 1'b0;
		16196: rom = 1'b0;
		16197: rom = 1'b0;
		16198: rom = 1'b0;
		16199: rom = 1'b0;
		16200: rom = 1'b0;
		16201: rom = 1'b0;
		16202: rom = 1'b0;
		16203: rom = 1'b0;
		16204: rom = 1'b0;
		16205: rom = 1'b0;
		16206: rom = 1'b0;
		16207: rom = 1'b0;
		16208: rom = 1'b0;
		16209: rom = 1'b0;
		16210: rom = 1'b0;
		16211: rom = 1'b0;
		16212: rom = 1'b0;
		16213: rom = 1'b0;
		16214: rom = 1'b0;
		16215: rom = 1'b0;
		16216: rom = 1'b0;
		16217: rom = 1'b0;
		16218: rom = 1'b0;
		16219: rom = 1'b0;
		16220: rom = 1'b0;
		16221: rom = 1'b0;
		16222: rom = 1'b0;
		16223: rom = 1'b0;
		16224: rom = 1'b0;
		16225: rom = 1'b0;
		16226: rom = 1'b0;
		16227: rom = 1'b0;
		16228: rom = 1'b0;
		16229: rom = 1'b0;
		16230: rom = 1'b0;
		16231: rom = 1'b0;
		16232: rom = 1'b0;
		16233: rom = 1'b0;
		16234: rom = 1'b0;
		16235: rom = 1'b0;
		16236: rom = 1'b0;
		16237: rom = 1'b0;
		16238: rom = 1'b0;
		16239: rom = 1'b0;
		16240: rom = 1'b0;
		16241: rom = 1'b0;
		16242: rom = 1'b0;
		16243: rom = 1'b0;
		16244: rom = 1'b0;
		16245: rom = 1'b0;
		16246: rom = 1'b0;
		16247: rom = 1'b0;
		16248: rom = 1'b0;
		16249: rom = 1'b0;
		16250: rom = 1'b0;
		16251: rom = 1'b0;
		16252: rom = 1'b0;
		16253: rom = 1'b0;
		16254: rom = 1'b0;
		16255: rom = 1'b0;
		16256: rom = 1'b0;
		16257: rom = 1'b0;
		16258: rom = 1'b0;
		16259: rom = 1'b0;
		16260: rom = 1'b0;
		16261: rom = 1'b0;
		16262: rom = 1'b0;
		16263: rom = 1'b0;
		16264: rom = 1'b0;
		16265: rom = 1'b0;
		16266: rom = 1'b0;
		16267: rom = 1'b0;
		16268: rom = 1'b0;
		16269: rom = 1'b0;
		16270: rom = 1'b0;
		16271: rom = 1'b0;
		16272: rom = 1'b0;
		16273: rom = 1'b0;
		16274: rom = 1'b0;
		16275: rom = 1'b0;
		16276: rom = 1'b0;
		16277: rom = 1'b0;
		16278: rom = 1'b0;
		16279: rom = 1'b0;
		16280: rom = 1'b0;
		16281: rom = 1'b0;
		16282: rom = 1'b0;
		16283: rom = 1'b0;
		16284: rom = 1'b0;
		16285: rom = 1'b0;
		16286: rom = 1'b0;
		16287: rom = 1'b0;
		16288: rom = 1'b0;
		16289: rom = 1'b0;
		16290: rom = 1'b0;
		16291: rom = 1'b0;
		16292: rom = 1'b0;
		16293: rom = 1'b0;
		16294: rom = 1'b0;
		16295: rom = 1'b0;
		16296: rom = 1'b0;
		16297: rom = 1'b0;
		16298: rom = 1'b0;
		16299: rom = 1'b0;
		16300: rom = 1'b0;
		16301: rom = 1'b0;
		16302: rom = 1'b0;
		16303: rom = 1'b0;
		16304: rom = 1'b0;
		16305: rom = 1'b0;
		16306: rom = 1'b0;
		16307: rom = 1'b0;
		16308: rom = 1'b0;
		16309: rom = 1'b0;
		16310: rom = 1'b0;
		16311: rom = 1'b0;
		16312: rom = 1'b0;
		16313: rom = 1'b0;
		16314: rom = 1'b0;
		16315: rom = 1'b0;
		16316: rom = 1'b0;
		16317: rom = 1'b0;
		16318: rom = 1'b0;
		16319: rom = 1'b0;
		16320: rom = 1'b0;
		16321: rom = 1'b0;
		16322: rom = 1'b0;
		16323: rom = 1'b0;
		16324: rom = 1'b0;
		16325: rom = 1'b0;
		16326: rom = 1'b0;
		16327: rom = 1'b0;
		16328: rom = 1'b0;
		16329: rom = 1'b0;
		16330: rom = 1'b0;
		16331: rom = 1'b0;
		16332: rom = 1'b0;
		16333: rom = 1'b0;
		16334: rom = 1'b0;
		16335: rom = 1'b0;
		16336: rom = 1'b0;
		16337: rom = 1'b0;
		16338: rom = 1'b0;
		16339: rom = 1'b0;
		16340: rom = 1'b0;
		16341: rom = 1'b0;
		16342: rom = 1'b0;
		16343: rom = 1'b0;
		16344: rom = 1'b0;
		16345: rom = 1'b0;
		16346: rom = 1'b0;
		16347: rom = 1'b0;
		16348: rom = 1'b0;
		16349: rom = 1'b0;
		16350: rom = 1'b0;
		16351: rom = 1'b0;
		16352: rom = 1'b0;
		16353: rom = 1'b0;
		16354: rom = 1'b0;
		16355: rom = 1'b0;
		16356: rom = 1'b0;
		16357: rom = 1'b0;
		16358: rom = 1'b0;
		16359: rom = 1'b0;
		16360: rom = 1'b0;
		16361: rom = 1'b0;
		16362: rom = 1'b0;
		16363: rom = 1'b0;
		16364: rom = 1'b0;
		16365: rom = 1'b0;
		16366: rom = 1'b0;
		16367: rom = 1'b0;
		16368: rom = 1'b0;
		16369: rom = 1'b0;
		16370: rom = 1'b0;
		16371: rom = 1'b0;
		16372: rom = 1'b0;
		16373: rom = 1'b0;
		16374: rom = 1'b0;
		16375: rom = 1'b0;
		16376: rom = 1'b0;
		16377: rom = 1'b0;
		16378: rom = 1'b0;
		16379: rom = 1'b0;
		16380: rom = 1'b0;
		16381: rom = 1'b0;
		16382: rom = 1'b0;
		16383: rom = 1'b0;
	endcase
end

endmodule
