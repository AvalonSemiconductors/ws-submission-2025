module tholin;
endmodule
