magic
tech gf180mcuD
magscale 1 10
timestamp 1762910469
<< pwell >>
rect -344 -2366 344 2366
<< mvpsubdiff >>
rect -312 2262 312 2334
rect -312 2218 -240 2262
rect -312 -2218 -299 2218
rect -253 -2218 -240 2218
rect 240 2218 312 2262
rect -312 -2262 -240 -2218
rect 240 -2218 253 2218
rect 299 -2218 312 2218
rect 240 -2262 312 -2218
rect -312 -2334 312 -2262
<< mvpsubdiffcont >>
rect -299 -2218 -253 2218
rect 253 -2218 299 2218
<< polysilicon >>
rect -100 2109 100 2122
rect -100 2063 -87 2109
rect 87 2063 100 2109
rect -100 2000 100 2063
rect -100 -2063 100 -2000
rect -100 -2109 -87 -2063
rect 87 -2109 100 -2063
rect -100 -2122 100 -2109
<< polycontact >>
rect -87 2063 87 2109
rect -87 -2109 87 -2063
<< mvnhighres >>
rect -100 -2000 100 2000
<< metal1 >>
rect -299 2275 299 2321
rect -299 2218 -253 2275
rect 253 2218 299 2275
rect -98 2063 -87 2109
rect 87 2063 98 2109
rect -98 -2109 -87 -2063
rect 87 -2109 98 -2063
rect -299 -2275 -253 -2218
rect 253 -2275 299 -2218
rect -299 -2321 299 -2275
<< properties >>
string FIXED_BBOX -276 -2298 276 2298
string gencell ppolyf_u_1k_6p0
string library gf180mcu
string parameters w 1.0 l 20.0 m 1 nx 1 wmin 1.000 lmin 1.000 class resistor rho 1000 val 20.0k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
