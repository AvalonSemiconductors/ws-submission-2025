magic
tech gf180mcuD
timestamp 1638034600
<< fillblock >>
rect 0 0 9000 10566
<< metal4 >>
rect 0 3438 18 3456
rect 0 3456 18 3474
rect 0 3474 18 3492
rect 0 3492 18 3510
rect 0 3510 18 3528
rect 0 3528 18 3546
rect 0 3546 18 3564
rect 0 3564 18 3582
rect 0 3582 18 3600
rect 0 3600 18 3618
rect 0 3618 18 3636
rect 0 3636 18 3654
rect 0 3654 18 3672
rect 0 3672 18 3690
rect 0 3690 18 3708
rect 0 3708 18 3726
rect 0 3726 18 3744
rect 0 3744 18 3762
rect 0 3762 18 3780
rect 0 3780 18 3798
rect 0 3798 18 3816
rect 0 3816 18 3834
rect 18 3222 36 3240
rect 18 3240 36 3258
rect 18 3258 36 3276
rect 18 3276 36 3294
rect 18 3294 36 3312
rect 18 3312 36 3330
rect 18 3330 36 3348
rect 18 3348 36 3366
rect 18 3366 36 3384
rect 18 3384 36 3402
rect 18 3402 36 3420
rect 18 3420 36 3438
rect 18 3438 36 3456
rect 18 3456 36 3474
rect 18 3474 36 3492
rect 18 3492 36 3510
rect 18 3510 36 3528
rect 18 3528 36 3546
rect 18 3546 36 3564
rect 18 3564 36 3582
rect 18 3582 36 3600
rect 18 3600 36 3618
rect 18 3618 36 3636
rect 18 3636 36 3654
rect 18 3654 36 3672
rect 18 3672 36 3690
rect 18 3690 36 3708
rect 18 3708 36 3726
rect 18 3726 36 3744
rect 18 3744 36 3762
rect 18 3762 36 3780
rect 18 3780 36 3798
rect 18 3798 36 3816
rect 18 3816 36 3834
rect 18 3834 36 3852
rect 18 3852 36 3870
rect 18 3870 36 3888
rect 18 3888 36 3906
rect 18 3906 36 3924
rect 18 3924 36 3942
rect 18 3942 36 3960
rect 18 3960 36 3978
rect 18 3978 36 3996
rect 18 3996 36 4014
rect 18 4014 36 4032
rect 18 4032 36 4050
rect 36 3096 54 3114
rect 36 3114 54 3132
rect 36 3132 54 3150
rect 36 3150 54 3168
rect 36 3168 54 3186
rect 36 3186 54 3204
rect 36 3204 54 3222
rect 36 3222 54 3240
rect 36 3240 54 3258
rect 36 3258 54 3276
rect 36 3276 54 3294
rect 36 3294 54 3312
rect 36 3312 54 3330
rect 36 3330 54 3348
rect 36 3348 54 3366
rect 36 3366 54 3384
rect 36 3384 54 3402
rect 36 3402 54 3420
rect 36 3420 54 3438
rect 36 3438 54 3456
rect 36 3456 54 3474
rect 36 3474 54 3492
rect 36 3492 54 3510
rect 36 3510 54 3528
rect 36 3528 54 3546
rect 36 3546 54 3564
rect 36 3564 54 3582
rect 36 3582 54 3600
rect 36 3600 54 3618
rect 36 3618 54 3636
rect 36 3636 54 3654
rect 36 3654 54 3672
rect 36 3672 54 3690
rect 36 3690 54 3708
rect 36 3708 54 3726
rect 36 3726 54 3744
rect 36 3744 54 3762
rect 36 3762 54 3780
rect 36 3780 54 3798
rect 36 3798 54 3816
rect 36 3816 54 3834
rect 36 3834 54 3852
rect 36 3852 54 3870
rect 36 3870 54 3888
rect 36 3888 54 3906
rect 36 3906 54 3924
rect 36 3924 54 3942
rect 36 3942 54 3960
rect 36 3960 54 3978
rect 36 3978 54 3996
rect 36 3996 54 4014
rect 36 4014 54 4032
rect 36 4032 54 4050
rect 36 4050 54 4068
rect 36 4068 54 4086
rect 36 4086 54 4104
rect 36 4104 54 4122
rect 36 4122 54 4140
rect 36 4140 54 4158
rect 36 4158 54 4176
rect 54 2988 72 3006
rect 54 3006 72 3024
rect 54 3024 72 3042
rect 54 3042 72 3060
rect 54 3060 72 3078
rect 54 3078 72 3096
rect 54 3096 72 3114
rect 54 3114 72 3132
rect 54 3132 72 3150
rect 54 3150 72 3168
rect 54 3168 72 3186
rect 54 3186 72 3204
rect 54 3204 72 3222
rect 54 3222 72 3240
rect 54 3240 72 3258
rect 54 3258 72 3276
rect 54 3276 72 3294
rect 54 3294 72 3312
rect 54 3312 72 3330
rect 54 3330 72 3348
rect 54 3348 72 3366
rect 54 3366 72 3384
rect 54 3384 72 3402
rect 54 3402 72 3420
rect 54 3420 72 3438
rect 54 3438 72 3456
rect 54 3456 72 3474
rect 54 3474 72 3492
rect 54 3492 72 3510
rect 54 3510 72 3528
rect 54 3528 72 3546
rect 54 3546 72 3564
rect 54 3564 72 3582
rect 54 3582 72 3600
rect 54 3600 72 3618
rect 54 3618 72 3636
rect 54 3636 72 3654
rect 54 3654 72 3672
rect 54 3672 72 3690
rect 54 3690 72 3708
rect 54 3708 72 3726
rect 54 3726 72 3744
rect 54 3744 72 3762
rect 54 3762 72 3780
rect 54 3780 72 3798
rect 54 3798 72 3816
rect 54 3816 72 3834
rect 54 3834 72 3852
rect 54 3852 72 3870
rect 54 3870 72 3888
rect 54 3888 72 3906
rect 54 3906 72 3924
rect 54 3924 72 3942
rect 54 3942 72 3960
rect 54 3960 72 3978
rect 54 3978 72 3996
rect 54 3996 72 4014
rect 54 4014 72 4032
rect 54 4032 72 4050
rect 54 4050 72 4068
rect 54 4068 72 4086
rect 54 4086 72 4104
rect 54 4104 72 4122
rect 54 4122 72 4140
rect 54 4140 72 4158
rect 54 4158 72 4176
rect 54 4176 72 4194
rect 54 4194 72 4212
rect 54 4212 72 4230
rect 54 4230 72 4248
rect 54 4248 72 4266
rect 54 4266 72 4284
rect 72 2880 90 2898
rect 72 2898 90 2916
rect 72 2916 90 2934
rect 72 2934 90 2952
rect 72 2952 90 2970
rect 72 2970 90 2988
rect 72 2988 90 3006
rect 72 3006 90 3024
rect 72 3024 90 3042
rect 72 3042 90 3060
rect 72 3060 90 3078
rect 72 3078 90 3096
rect 72 3096 90 3114
rect 72 3114 90 3132
rect 72 3132 90 3150
rect 72 3150 90 3168
rect 72 3168 90 3186
rect 72 3186 90 3204
rect 72 3204 90 3222
rect 72 3222 90 3240
rect 72 3240 90 3258
rect 72 3258 90 3276
rect 72 3276 90 3294
rect 72 3294 90 3312
rect 72 3312 90 3330
rect 72 3330 90 3348
rect 72 3348 90 3366
rect 72 3366 90 3384
rect 72 3384 90 3402
rect 72 3402 90 3420
rect 72 3420 90 3438
rect 72 3438 90 3456
rect 72 3456 90 3474
rect 72 3474 90 3492
rect 72 3492 90 3510
rect 72 3510 90 3528
rect 72 3528 90 3546
rect 72 3546 90 3564
rect 72 3564 90 3582
rect 72 3582 90 3600
rect 72 3600 90 3618
rect 72 3618 90 3636
rect 72 3636 90 3654
rect 72 3654 90 3672
rect 72 3672 90 3690
rect 72 3690 90 3708
rect 72 3708 90 3726
rect 72 3726 90 3744
rect 72 3744 90 3762
rect 72 3762 90 3780
rect 72 3780 90 3798
rect 72 3798 90 3816
rect 72 3816 90 3834
rect 72 3834 90 3852
rect 72 3852 90 3870
rect 72 3870 90 3888
rect 72 3888 90 3906
rect 72 3906 90 3924
rect 72 3924 90 3942
rect 72 3942 90 3960
rect 72 3960 90 3978
rect 72 3978 90 3996
rect 72 3996 90 4014
rect 72 4014 90 4032
rect 72 4032 90 4050
rect 72 4050 90 4068
rect 72 4068 90 4086
rect 72 4086 90 4104
rect 72 4104 90 4122
rect 72 4122 90 4140
rect 72 4140 90 4158
rect 72 4158 90 4176
rect 72 4176 90 4194
rect 72 4194 90 4212
rect 72 4212 90 4230
rect 72 4230 90 4248
rect 72 4248 90 4266
rect 72 4266 90 4284
rect 72 4284 90 4302
rect 72 4302 90 4320
rect 72 4320 90 4338
rect 72 4338 90 4356
rect 72 4356 90 4374
rect 90 2808 108 2826
rect 90 2826 108 2844
rect 90 2844 108 2862
rect 90 2862 108 2880
rect 90 2880 108 2898
rect 90 2898 108 2916
rect 90 2916 108 2934
rect 90 2934 108 2952
rect 90 2952 108 2970
rect 90 2970 108 2988
rect 90 2988 108 3006
rect 90 3006 108 3024
rect 90 3024 108 3042
rect 90 3042 108 3060
rect 90 3060 108 3078
rect 90 3078 108 3096
rect 90 3096 108 3114
rect 90 3114 108 3132
rect 90 3132 108 3150
rect 90 3150 108 3168
rect 90 3168 108 3186
rect 90 3186 108 3204
rect 90 3204 108 3222
rect 90 3222 108 3240
rect 90 3240 108 3258
rect 90 3258 108 3276
rect 90 3276 108 3294
rect 90 3294 108 3312
rect 90 3312 108 3330
rect 90 3330 108 3348
rect 90 3348 108 3366
rect 90 3366 108 3384
rect 90 3384 108 3402
rect 90 3402 108 3420
rect 90 3420 108 3438
rect 90 3438 108 3456
rect 90 3456 108 3474
rect 90 3474 108 3492
rect 90 3492 108 3510
rect 90 3510 108 3528
rect 90 3528 108 3546
rect 90 3546 108 3564
rect 90 3564 108 3582
rect 90 3582 108 3600
rect 90 3600 108 3618
rect 90 3618 108 3636
rect 90 3636 108 3654
rect 90 3654 108 3672
rect 90 3672 108 3690
rect 90 3690 108 3708
rect 90 3708 108 3726
rect 90 3726 108 3744
rect 90 3744 108 3762
rect 90 3762 108 3780
rect 90 3780 108 3798
rect 90 3798 108 3816
rect 90 3816 108 3834
rect 90 3834 108 3852
rect 90 3852 108 3870
rect 90 3870 108 3888
rect 90 3888 108 3906
rect 90 3906 108 3924
rect 90 3924 108 3942
rect 90 3942 108 3960
rect 90 3960 108 3978
rect 90 3978 108 3996
rect 90 3996 108 4014
rect 90 4014 108 4032
rect 90 4032 108 4050
rect 90 4050 108 4068
rect 90 4068 108 4086
rect 90 4086 108 4104
rect 90 4104 108 4122
rect 90 4122 108 4140
rect 90 4140 108 4158
rect 90 4158 108 4176
rect 90 4176 108 4194
rect 90 4194 108 4212
rect 90 4212 108 4230
rect 90 4230 108 4248
rect 90 4248 108 4266
rect 90 4266 108 4284
rect 90 4284 108 4302
rect 90 4302 108 4320
rect 90 4320 108 4338
rect 90 4338 108 4356
rect 90 4356 108 4374
rect 90 4374 108 4392
rect 90 4392 108 4410
rect 90 4410 108 4428
rect 90 4428 108 4446
rect 90 4446 108 4464
rect 108 2736 126 2754
rect 108 2754 126 2772
rect 108 2772 126 2790
rect 108 2790 126 2808
rect 108 2808 126 2826
rect 108 2826 126 2844
rect 108 2844 126 2862
rect 108 2862 126 2880
rect 108 2880 126 2898
rect 108 2898 126 2916
rect 108 2916 126 2934
rect 108 2934 126 2952
rect 108 2952 126 2970
rect 108 2970 126 2988
rect 108 2988 126 3006
rect 108 3006 126 3024
rect 108 3024 126 3042
rect 108 3042 126 3060
rect 108 3060 126 3078
rect 108 3078 126 3096
rect 108 3096 126 3114
rect 108 3114 126 3132
rect 108 3132 126 3150
rect 108 3150 126 3168
rect 108 3168 126 3186
rect 108 3186 126 3204
rect 108 3204 126 3222
rect 108 3222 126 3240
rect 108 3240 126 3258
rect 108 3258 126 3276
rect 108 3276 126 3294
rect 108 3294 126 3312
rect 108 3312 126 3330
rect 108 3330 126 3348
rect 108 3348 126 3366
rect 108 3366 126 3384
rect 108 3384 126 3402
rect 108 3402 126 3420
rect 108 3420 126 3438
rect 108 3438 126 3456
rect 108 3456 126 3474
rect 108 3474 126 3492
rect 108 3492 126 3510
rect 108 3510 126 3528
rect 108 3528 126 3546
rect 108 3546 126 3564
rect 108 3564 126 3582
rect 108 3582 126 3600
rect 108 3600 126 3618
rect 108 3618 126 3636
rect 108 3636 126 3654
rect 108 3654 126 3672
rect 108 3672 126 3690
rect 108 3690 126 3708
rect 108 3708 126 3726
rect 108 3726 126 3744
rect 108 3744 126 3762
rect 108 3762 126 3780
rect 108 3780 126 3798
rect 108 3798 126 3816
rect 108 3816 126 3834
rect 108 3834 126 3852
rect 108 3852 126 3870
rect 108 3870 126 3888
rect 108 3888 126 3906
rect 108 3906 126 3924
rect 108 3924 126 3942
rect 108 3942 126 3960
rect 108 3960 126 3978
rect 108 3978 126 3996
rect 108 3996 126 4014
rect 108 4014 126 4032
rect 108 4032 126 4050
rect 108 4050 126 4068
rect 108 4068 126 4086
rect 108 4086 126 4104
rect 108 4104 126 4122
rect 108 4122 126 4140
rect 108 4140 126 4158
rect 108 4158 126 4176
rect 108 4176 126 4194
rect 108 4194 126 4212
rect 108 4212 126 4230
rect 108 4230 126 4248
rect 108 4248 126 4266
rect 108 4266 126 4284
rect 108 4284 126 4302
rect 108 4302 126 4320
rect 108 4320 126 4338
rect 108 4338 126 4356
rect 108 4356 126 4374
rect 108 4374 126 4392
rect 108 4392 126 4410
rect 108 4410 126 4428
rect 108 4428 126 4446
rect 108 4446 126 4464
rect 108 4464 126 4482
rect 108 4482 126 4500
rect 108 4500 126 4518
rect 108 4518 126 4536
rect 126 2664 144 2682
rect 126 2682 144 2700
rect 126 2700 144 2718
rect 126 2718 144 2736
rect 126 2736 144 2754
rect 126 2754 144 2772
rect 126 2772 144 2790
rect 126 2790 144 2808
rect 126 2808 144 2826
rect 126 2826 144 2844
rect 126 2844 144 2862
rect 126 2862 144 2880
rect 126 2880 144 2898
rect 126 2898 144 2916
rect 126 2916 144 2934
rect 126 2934 144 2952
rect 126 2952 144 2970
rect 126 2970 144 2988
rect 126 2988 144 3006
rect 126 3006 144 3024
rect 126 3024 144 3042
rect 126 3042 144 3060
rect 126 3060 144 3078
rect 126 3078 144 3096
rect 126 3096 144 3114
rect 126 3114 144 3132
rect 126 3132 144 3150
rect 126 3150 144 3168
rect 126 3168 144 3186
rect 126 3186 144 3204
rect 126 3204 144 3222
rect 126 3222 144 3240
rect 126 3240 144 3258
rect 126 3258 144 3276
rect 126 3276 144 3294
rect 126 3294 144 3312
rect 126 3312 144 3330
rect 126 3330 144 3348
rect 126 3348 144 3366
rect 126 3366 144 3384
rect 126 3384 144 3402
rect 126 3402 144 3420
rect 126 3420 144 3438
rect 126 3438 144 3456
rect 126 3456 144 3474
rect 126 3474 144 3492
rect 126 3492 144 3510
rect 126 3510 144 3528
rect 126 3528 144 3546
rect 126 3546 144 3564
rect 126 3564 144 3582
rect 126 3582 144 3600
rect 126 3600 144 3618
rect 126 3618 144 3636
rect 126 3636 144 3654
rect 126 3654 144 3672
rect 126 3672 144 3690
rect 126 3690 144 3708
rect 126 3708 144 3726
rect 126 3726 144 3744
rect 126 3744 144 3762
rect 126 3762 144 3780
rect 126 3780 144 3798
rect 126 3798 144 3816
rect 126 3816 144 3834
rect 126 3834 144 3852
rect 126 3852 144 3870
rect 126 3870 144 3888
rect 126 3888 144 3906
rect 126 3906 144 3924
rect 126 3924 144 3942
rect 126 3942 144 3960
rect 126 3960 144 3978
rect 126 3978 144 3996
rect 126 3996 144 4014
rect 126 4014 144 4032
rect 126 4032 144 4050
rect 126 4050 144 4068
rect 126 4068 144 4086
rect 126 4086 144 4104
rect 126 4104 144 4122
rect 126 4122 144 4140
rect 126 4140 144 4158
rect 126 4158 144 4176
rect 126 4176 144 4194
rect 126 4194 144 4212
rect 126 4212 144 4230
rect 126 4230 144 4248
rect 126 4248 144 4266
rect 126 4266 144 4284
rect 126 4284 144 4302
rect 126 4302 144 4320
rect 126 4320 144 4338
rect 126 4338 144 4356
rect 126 4356 144 4374
rect 126 4374 144 4392
rect 126 4392 144 4410
rect 126 4410 144 4428
rect 126 4428 144 4446
rect 126 4446 144 4464
rect 126 4464 144 4482
rect 126 4482 144 4500
rect 126 4500 144 4518
rect 126 4518 144 4536
rect 126 4536 144 4554
rect 126 4554 144 4572
rect 126 4572 144 4590
rect 126 4590 144 4608
rect 144 2610 162 2628
rect 144 2628 162 2646
rect 144 2646 162 2664
rect 144 2664 162 2682
rect 144 2682 162 2700
rect 144 2700 162 2718
rect 144 2718 162 2736
rect 144 2736 162 2754
rect 144 2754 162 2772
rect 144 2772 162 2790
rect 144 2790 162 2808
rect 144 2808 162 2826
rect 144 2826 162 2844
rect 144 2844 162 2862
rect 144 2862 162 2880
rect 144 2880 162 2898
rect 144 2898 162 2916
rect 144 2916 162 2934
rect 144 2934 162 2952
rect 144 2952 162 2970
rect 144 2970 162 2988
rect 144 2988 162 3006
rect 144 3006 162 3024
rect 144 3024 162 3042
rect 144 3042 162 3060
rect 144 3060 162 3078
rect 144 3078 162 3096
rect 144 3096 162 3114
rect 144 3114 162 3132
rect 144 3132 162 3150
rect 144 3150 162 3168
rect 144 3168 162 3186
rect 144 3186 162 3204
rect 144 3204 162 3222
rect 144 3222 162 3240
rect 144 3240 162 3258
rect 144 3258 162 3276
rect 144 3276 162 3294
rect 144 3294 162 3312
rect 144 3312 162 3330
rect 144 3330 162 3348
rect 144 3348 162 3366
rect 144 3366 162 3384
rect 144 3384 162 3402
rect 144 3402 162 3420
rect 144 3420 162 3438
rect 144 3438 162 3456
rect 144 3456 162 3474
rect 144 3474 162 3492
rect 144 3492 162 3510
rect 144 3510 162 3528
rect 144 3528 162 3546
rect 144 3546 162 3564
rect 144 3564 162 3582
rect 144 3582 162 3600
rect 144 3600 162 3618
rect 144 3618 162 3636
rect 144 3636 162 3654
rect 144 3654 162 3672
rect 144 3672 162 3690
rect 144 3690 162 3708
rect 144 3708 162 3726
rect 144 3726 162 3744
rect 144 3744 162 3762
rect 144 3762 162 3780
rect 144 3780 162 3798
rect 144 3798 162 3816
rect 144 3816 162 3834
rect 144 3834 162 3852
rect 144 3852 162 3870
rect 144 3870 162 3888
rect 144 3888 162 3906
rect 144 3906 162 3924
rect 144 3924 162 3942
rect 144 3942 162 3960
rect 144 3960 162 3978
rect 144 3978 162 3996
rect 144 3996 162 4014
rect 144 4014 162 4032
rect 144 4032 162 4050
rect 144 4050 162 4068
rect 144 4068 162 4086
rect 144 4086 162 4104
rect 144 4104 162 4122
rect 144 4122 162 4140
rect 144 4140 162 4158
rect 144 4158 162 4176
rect 144 4176 162 4194
rect 144 4194 162 4212
rect 144 4212 162 4230
rect 144 4230 162 4248
rect 144 4248 162 4266
rect 144 4266 162 4284
rect 144 4284 162 4302
rect 144 4302 162 4320
rect 144 4320 162 4338
rect 144 4338 162 4356
rect 144 4356 162 4374
rect 144 4374 162 4392
rect 144 4392 162 4410
rect 144 4410 162 4428
rect 144 4428 162 4446
rect 144 4446 162 4464
rect 144 4464 162 4482
rect 144 4482 162 4500
rect 144 4500 162 4518
rect 144 4518 162 4536
rect 144 4536 162 4554
rect 144 4554 162 4572
rect 144 4572 162 4590
rect 144 4590 162 4608
rect 144 4608 162 4626
rect 144 4626 162 4644
rect 144 4644 162 4662
rect 162 2538 180 2556
rect 162 2556 180 2574
rect 162 2574 180 2592
rect 162 2592 180 2610
rect 162 2610 180 2628
rect 162 2628 180 2646
rect 162 2646 180 2664
rect 162 2664 180 2682
rect 162 2682 180 2700
rect 162 2700 180 2718
rect 162 2718 180 2736
rect 162 2736 180 2754
rect 162 2754 180 2772
rect 162 2772 180 2790
rect 162 2790 180 2808
rect 162 2808 180 2826
rect 162 2826 180 2844
rect 162 2844 180 2862
rect 162 2862 180 2880
rect 162 2880 180 2898
rect 162 2898 180 2916
rect 162 2916 180 2934
rect 162 2934 180 2952
rect 162 2952 180 2970
rect 162 2970 180 2988
rect 162 2988 180 3006
rect 162 3006 180 3024
rect 162 3024 180 3042
rect 162 3042 180 3060
rect 162 3060 180 3078
rect 162 3078 180 3096
rect 162 3096 180 3114
rect 162 3114 180 3132
rect 162 3132 180 3150
rect 162 3150 180 3168
rect 162 3168 180 3186
rect 162 3186 180 3204
rect 162 3204 180 3222
rect 162 3222 180 3240
rect 162 3240 180 3258
rect 162 3258 180 3276
rect 162 3276 180 3294
rect 162 3294 180 3312
rect 162 3312 180 3330
rect 162 3330 180 3348
rect 162 3348 180 3366
rect 162 3366 180 3384
rect 162 3384 180 3402
rect 162 3402 180 3420
rect 162 3420 180 3438
rect 162 3438 180 3456
rect 162 3456 180 3474
rect 162 3474 180 3492
rect 162 3492 180 3510
rect 162 3510 180 3528
rect 162 3528 180 3546
rect 162 3546 180 3564
rect 162 3564 180 3582
rect 162 3582 180 3600
rect 162 3600 180 3618
rect 162 3618 180 3636
rect 162 3636 180 3654
rect 162 3654 180 3672
rect 162 3672 180 3690
rect 162 3690 180 3708
rect 162 3708 180 3726
rect 162 3726 180 3744
rect 162 3744 180 3762
rect 162 3762 180 3780
rect 162 3780 180 3798
rect 162 3798 180 3816
rect 162 3816 180 3834
rect 162 3834 180 3852
rect 162 3852 180 3870
rect 162 3870 180 3888
rect 162 3888 180 3906
rect 162 3906 180 3924
rect 162 3924 180 3942
rect 162 3942 180 3960
rect 162 3960 180 3978
rect 162 3978 180 3996
rect 162 3996 180 4014
rect 162 4014 180 4032
rect 162 4032 180 4050
rect 162 4050 180 4068
rect 162 4068 180 4086
rect 162 4086 180 4104
rect 162 4104 180 4122
rect 162 4122 180 4140
rect 162 4140 180 4158
rect 162 4158 180 4176
rect 162 4176 180 4194
rect 162 4194 180 4212
rect 162 4212 180 4230
rect 162 4230 180 4248
rect 162 4248 180 4266
rect 162 4266 180 4284
rect 162 4284 180 4302
rect 162 4302 180 4320
rect 162 4320 180 4338
rect 162 4338 180 4356
rect 162 4356 180 4374
rect 162 4374 180 4392
rect 162 4392 180 4410
rect 162 4410 180 4428
rect 162 4428 180 4446
rect 162 4446 180 4464
rect 162 4464 180 4482
rect 162 4482 180 4500
rect 162 4500 180 4518
rect 162 4518 180 4536
rect 162 4536 180 4554
rect 162 4554 180 4572
rect 162 4572 180 4590
rect 162 4590 180 4608
rect 162 4608 180 4626
rect 162 4626 180 4644
rect 162 4644 180 4662
rect 162 4662 180 4680
rect 162 4680 180 4698
rect 162 4698 180 4716
rect 162 4716 180 4734
rect 180 2484 198 2502
rect 180 2502 198 2520
rect 180 2520 198 2538
rect 180 2538 198 2556
rect 180 2556 198 2574
rect 180 2574 198 2592
rect 180 2592 198 2610
rect 180 2610 198 2628
rect 180 2628 198 2646
rect 180 2646 198 2664
rect 180 2664 198 2682
rect 180 2682 198 2700
rect 180 2700 198 2718
rect 180 2718 198 2736
rect 180 2736 198 2754
rect 180 2754 198 2772
rect 180 2772 198 2790
rect 180 2790 198 2808
rect 180 2808 198 2826
rect 180 2826 198 2844
rect 180 2844 198 2862
rect 180 2862 198 2880
rect 180 2880 198 2898
rect 180 2898 198 2916
rect 180 2916 198 2934
rect 180 2934 198 2952
rect 180 2952 198 2970
rect 180 2970 198 2988
rect 180 2988 198 3006
rect 180 3006 198 3024
rect 180 3024 198 3042
rect 180 3042 198 3060
rect 180 3060 198 3078
rect 180 3078 198 3096
rect 180 3096 198 3114
rect 180 3114 198 3132
rect 180 3132 198 3150
rect 180 3150 198 3168
rect 180 3168 198 3186
rect 180 3186 198 3204
rect 180 3204 198 3222
rect 180 3222 198 3240
rect 180 3240 198 3258
rect 180 3258 198 3276
rect 180 3276 198 3294
rect 180 3294 198 3312
rect 180 3312 198 3330
rect 180 3330 198 3348
rect 180 3348 198 3366
rect 180 3366 198 3384
rect 180 3384 198 3402
rect 180 3402 198 3420
rect 180 3420 198 3438
rect 180 3438 198 3456
rect 180 3456 198 3474
rect 180 3474 198 3492
rect 180 3492 198 3510
rect 180 3510 198 3528
rect 180 3528 198 3546
rect 180 3546 198 3564
rect 180 3564 198 3582
rect 180 3582 198 3600
rect 180 3600 198 3618
rect 180 3618 198 3636
rect 180 3636 198 3654
rect 180 3654 198 3672
rect 180 3672 198 3690
rect 180 3690 198 3708
rect 180 3708 198 3726
rect 180 3726 198 3744
rect 180 3744 198 3762
rect 180 3762 198 3780
rect 180 3780 198 3798
rect 180 3798 198 3816
rect 180 3816 198 3834
rect 180 3834 198 3852
rect 180 3852 198 3870
rect 180 3870 198 3888
rect 180 3888 198 3906
rect 180 3906 198 3924
rect 180 3924 198 3942
rect 180 3942 198 3960
rect 180 3960 198 3978
rect 180 3978 198 3996
rect 180 3996 198 4014
rect 180 4014 198 4032
rect 180 4032 198 4050
rect 180 4050 198 4068
rect 180 4068 198 4086
rect 180 4086 198 4104
rect 180 4104 198 4122
rect 180 4122 198 4140
rect 180 4140 198 4158
rect 180 4158 198 4176
rect 180 4176 198 4194
rect 180 4194 198 4212
rect 180 4212 198 4230
rect 180 4230 198 4248
rect 180 4248 198 4266
rect 180 4266 198 4284
rect 180 4284 198 4302
rect 180 4302 198 4320
rect 180 4320 198 4338
rect 180 4338 198 4356
rect 180 4356 198 4374
rect 180 4374 198 4392
rect 180 4392 198 4410
rect 180 4410 198 4428
rect 180 4428 198 4446
rect 180 4446 198 4464
rect 180 4464 198 4482
rect 180 4482 198 4500
rect 180 4500 198 4518
rect 180 4518 198 4536
rect 180 4536 198 4554
rect 180 4554 198 4572
rect 180 4572 198 4590
rect 180 4590 198 4608
rect 180 4608 198 4626
rect 180 4626 198 4644
rect 180 4644 198 4662
rect 180 4662 198 4680
rect 180 4680 198 4698
rect 180 4698 198 4716
rect 180 4716 198 4734
rect 180 4734 198 4752
rect 180 4752 198 4770
rect 180 4770 198 4788
rect 198 2430 216 2448
rect 198 2448 216 2466
rect 198 2466 216 2484
rect 198 2484 216 2502
rect 198 2502 216 2520
rect 198 2520 216 2538
rect 198 2538 216 2556
rect 198 2556 216 2574
rect 198 2574 216 2592
rect 198 2592 216 2610
rect 198 2610 216 2628
rect 198 2628 216 2646
rect 198 2646 216 2664
rect 198 2664 216 2682
rect 198 2682 216 2700
rect 198 2700 216 2718
rect 198 2718 216 2736
rect 198 2736 216 2754
rect 198 2754 216 2772
rect 198 2772 216 2790
rect 198 2790 216 2808
rect 198 2808 216 2826
rect 198 2826 216 2844
rect 198 2844 216 2862
rect 198 2862 216 2880
rect 198 2880 216 2898
rect 198 2898 216 2916
rect 198 2916 216 2934
rect 198 2934 216 2952
rect 198 2952 216 2970
rect 198 2970 216 2988
rect 198 2988 216 3006
rect 198 3006 216 3024
rect 198 3024 216 3042
rect 198 3042 216 3060
rect 198 3060 216 3078
rect 198 3078 216 3096
rect 198 3096 216 3114
rect 198 3114 216 3132
rect 198 3132 216 3150
rect 198 3150 216 3168
rect 198 3168 216 3186
rect 198 3186 216 3204
rect 198 3204 216 3222
rect 198 3222 216 3240
rect 198 3240 216 3258
rect 198 3258 216 3276
rect 198 3276 216 3294
rect 198 3294 216 3312
rect 198 3312 216 3330
rect 198 3330 216 3348
rect 198 3348 216 3366
rect 198 3366 216 3384
rect 198 3384 216 3402
rect 198 3402 216 3420
rect 198 3420 216 3438
rect 198 3438 216 3456
rect 198 3456 216 3474
rect 198 3474 216 3492
rect 198 3492 216 3510
rect 198 3510 216 3528
rect 198 3528 216 3546
rect 198 3546 216 3564
rect 198 3564 216 3582
rect 198 3582 216 3600
rect 198 3600 216 3618
rect 198 3618 216 3636
rect 198 3636 216 3654
rect 198 3654 216 3672
rect 198 3672 216 3690
rect 198 3690 216 3708
rect 198 3708 216 3726
rect 198 3726 216 3744
rect 198 3744 216 3762
rect 198 3762 216 3780
rect 198 3780 216 3798
rect 198 3798 216 3816
rect 198 3816 216 3834
rect 198 3834 216 3852
rect 198 3852 216 3870
rect 198 3870 216 3888
rect 198 3888 216 3906
rect 198 3906 216 3924
rect 198 3924 216 3942
rect 198 3942 216 3960
rect 198 3960 216 3978
rect 198 3978 216 3996
rect 198 3996 216 4014
rect 198 4014 216 4032
rect 198 4032 216 4050
rect 198 4050 216 4068
rect 198 4068 216 4086
rect 198 4086 216 4104
rect 198 4104 216 4122
rect 198 4122 216 4140
rect 198 4140 216 4158
rect 198 4158 216 4176
rect 198 4176 216 4194
rect 198 4194 216 4212
rect 198 4212 216 4230
rect 198 4230 216 4248
rect 198 4248 216 4266
rect 198 4266 216 4284
rect 198 4284 216 4302
rect 198 4302 216 4320
rect 198 4320 216 4338
rect 198 4338 216 4356
rect 198 4356 216 4374
rect 198 4374 216 4392
rect 198 4392 216 4410
rect 198 4410 216 4428
rect 198 4428 216 4446
rect 198 4446 216 4464
rect 198 4464 216 4482
rect 198 4482 216 4500
rect 198 4500 216 4518
rect 198 4518 216 4536
rect 198 4536 216 4554
rect 198 4554 216 4572
rect 198 4572 216 4590
rect 198 4590 216 4608
rect 198 4608 216 4626
rect 198 4626 216 4644
rect 198 4644 216 4662
rect 198 4662 216 4680
rect 198 4680 216 4698
rect 198 4698 216 4716
rect 198 4716 216 4734
rect 198 4734 216 4752
rect 198 4752 216 4770
rect 198 4770 216 4788
rect 198 4788 216 4806
rect 198 4806 216 4824
rect 198 4824 216 4842
rect 216 2394 234 2412
rect 216 2412 234 2430
rect 216 2430 234 2448
rect 216 2448 234 2466
rect 216 2466 234 2484
rect 216 2484 234 2502
rect 216 2502 234 2520
rect 216 2520 234 2538
rect 216 2538 234 2556
rect 216 2556 234 2574
rect 216 2574 234 2592
rect 216 2592 234 2610
rect 216 2610 234 2628
rect 216 2628 234 2646
rect 216 2646 234 2664
rect 216 2664 234 2682
rect 216 2682 234 2700
rect 216 2700 234 2718
rect 216 2718 234 2736
rect 216 2736 234 2754
rect 216 2754 234 2772
rect 216 2772 234 2790
rect 216 2790 234 2808
rect 216 2808 234 2826
rect 216 2826 234 2844
rect 216 2844 234 2862
rect 216 2862 234 2880
rect 216 2880 234 2898
rect 216 2898 234 2916
rect 216 2916 234 2934
rect 216 2934 234 2952
rect 216 2952 234 2970
rect 216 2970 234 2988
rect 216 2988 234 3006
rect 216 3006 234 3024
rect 216 3024 234 3042
rect 216 3042 234 3060
rect 216 3060 234 3078
rect 216 3078 234 3096
rect 216 3096 234 3114
rect 216 3114 234 3132
rect 216 3132 234 3150
rect 216 3150 234 3168
rect 216 3168 234 3186
rect 216 3186 234 3204
rect 216 3204 234 3222
rect 216 3222 234 3240
rect 216 3240 234 3258
rect 216 3258 234 3276
rect 216 3276 234 3294
rect 216 3294 234 3312
rect 216 3312 234 3330
rect 216 3330 234 3348
rect 216 3348 234 3366
rect 216 3366 234 3384
rect 216 3384 234 3402
rect 216 3402 234 3420
rect 216 3420 234 3438
rect 216 3438 234 3456
rect 216 3456 234 3474
rect 216 3474 234 3492
rect 216 3492 234 3510
rect 216 3510 234 3528
rect 216 3528 234 3546
rect 216 3546 234 3564
rect 216 3564 234 3582
rect 216 3582 234 3600
rect 216 3600 234 3618
rect 216 3618 234 3636
rect 216 3636 234 3654
rect 216 3654 234 3672
rect 216 3672 234 3690
rect 216 3690 234 3708
rect 216 3708 234 3726
rect 216 3726 234 3744
rect 216 3744 234 3762
rect 216 3762 234 3780
rect 216 3780 234 3798
rect 216 3798 234 3816
rect 216 3816 234 3834
rect 216 3834 234 3852
rect 216 3852 234 3870
rect 216 3870 234 3888
rect 216 3888 234 3906
rect 216 3906 234 3924
rect 216 3924 234 3942
rect 216 3942 234 3960
rect 216 3960 234 3978
rect 216 3978 234 3996
rect 216 3996 234 4014
rect 216 4014 234 4032
rect 216 4032 234 4050
rect 216 4050 234 4068
rect 216 4068 234 4086
rect 216 4086 234 4104
rect 216 4104 234 4122
rect 216 4122 234 4140
rect 216 4140 234 4158
rect 216 4158 234 4176
rect 216 4176 234 4194
rect 216 4194 234 4212
rect 216 4212 234 4230
rect 216 4230 234 4248
rect 216 4248 234 4266
rect 216 4266 234 4284
rect 216 4284 234 4302
rect 216 4302 234 4320
rect 216 4320 234 4338
rect 216 4338 234 4356
rect 216 4356 234 4374
rect 216 4374 234 4392
rect 216 4392 234 4410
rect 216 4410 234 4428
rect 216 4428 234 4446
rect 216 4446 234 4464
rect 216 4464 234 4482
rect 216 4482 234 4500
rect 216 4500 234 4518
rect 216 4518 234 4536
rect 216 4536 234 4554
rect 216 4554 234 4572
rect 216 4572 234 4590
rect 216 4590 234 4608
rect 216 4608 234 4626
rect 216 4626 234 4644
rect 216 4644 234 4662
rect 216 4662 234 4680
rect 216 4680 234 4698
rect 216 4698 234 4716
rect 216 4716 234 4734
rect 216 4734 234 4752
rect 216 4752 234 4770
rect 216 4770 234 4788
rect 216 4788 234 4806
rect 216 4806 234 4824
rect 216 4824 234 4842
rect 216 4842 234 4860
rect 216 4860 234 4878
rect 234 2340 252 2358
rect 234 2358 252 2376
rect 234 2376 252 2394
rect 234 2394 252 2412
rect 234 2412 252 2430
rect 234 2430 252 2448
rect 234 2448 252 2466
rect 234 2466 252 2484
rect 234 2484 252 2502
rect 234 2502 252 2520
rect 234 2520 252 2538
rect 234 2538 252 2556
rect 234 2556 252 2574
rect 234 2574 252 2592
rect 234 2592 252 2610
rect 234 2610 252 2628
rect 234 2628 252 2646
rect 234 2646 252 2664
rect 234 2664 252 2682
rect 234 2682 252 2700
rect 234 2700 252 2718
rect 234 2718 252 2736
rect 234 2736 252 2754
rect 234 2754 252 2772
rect 234 2772 252 2790
rect 234 2790 252 2808
rect 234 2808 252 2826
rect 234 2826 252 2844
rect 234 2844 252 2862
rect 234 2862 252 2880
rect 234 2880 252 2898
rect 234 2898 252 2916
rect 234 2916 252 2934
rect 234 2934 252 2952
rect 234 2952 252 2970
rect 234 2970 252 2988
rect 234 2988 252 3006
rect 234 3006 252 3024
rect 234 3024 252 3042
rect 234 3042 252 3060
rect 234 3060 252 3078
rect 234 3078 252 3096
rect 234 3096 252 3114
rect 234 3114 252 3132
rect 234 3132 252 3150
rect 234 3150 252 3168
rect 234 3168 252 3186
rect 234 3186 252 3204
rect 234 3204 252 3222
rect 234 3222 252 3240
rect 234 3240 252 3258
rect 234 3258 252 3276
rect 234 3276 252 3294
rect 234 3294 252 3312
rect 234 3312 252 3330
rect 234 3330 252 3348
rect 234 3348 252 3366
rect 234 3366 252 3384
rect 234 3384 252 3402
rect 234 3402 252 3420
rect 234 3420 252 3438
rect 234 3438 252 3456
rect 234 3456 252 3474
rect 234 3474 252 3492
rect 234 3492 252 3510
rect 234 3510 252 3528
rect 234 3528 252 3546
rect 234 3546 252 3564
rect 234 3564 252 3582
rect 234 3582 252 3600
rect 234 3600 252 3618
rect 234 3618 252 3636
rect 234 3636 252 3654
rect 234 3654 252 3672
rect 234 3672 252 3690
rect 234 3690 252 3708
rect 234 3708 252 3726
rect 234 3726 252 3744
rect 234 3744 252 3762
rect 234 3762 252 3780
rect 234 3780 252 3798
rect 234 3798 252 3816
rect 234 3816 252 3834
rect 234 3834 252 3852
rect 234 3852 252 3870
rect 234 3870 252 3888
rect 234 3888 252 3906
rect 234 3906 252 3924
rect 234 3924 252 3942
rect 234 3942 252 3960
rect 234 3960 252 3978
rect 234 3978 252 3996
rect 234 3996 252 4014
rect 234 4014 252 4032
rect 234 4032 252 4050
rect 234 4050 252 4068
rect 234 4068 252 4086
rect 234 4086 252 4104
rect 234 4104 252 4122
rect 234 4122 252 4140
rect 234 4140 252 4158
rect 234 4158 252 4176
rect 234 4176 252 4194
rect 234 4194 252 4212
rect 234 4212 252 4230
rect 234 4230 252 4248
rect 234 4248 252 4266
rect 234 4266 252 4284
rect 234 4284 252 4302
rect 234 4302 252 4320
rect 234 4320 252 4338
rect 234 4338 252 4356
rect 234 4356 252 4374
rect 234 4374 252 4392
rect 234 4392 252 4410
rect 234 4410 252 4428
rect 234 4428 252 4446
rect 234 4446 252 4464
rect 234 4464 252 4482
rect 234 4482 252 4500
rect 234 4500 252 4518
rect 234 4518 252 4536
rect 234 4536 252 4554
rect 234 4554 252 4572
rect 234 4572 252 4590
rect 234 4590 252 4608
rect 234 4608 252 4626
rect 234 4626 252 4644
rect 234 4644 252 4662
rect 234 4662 252 4680
rect 234 4680 252 4698
rect 234 4698 252 4716
rect 234 4716 252 4734
rect 234 4734 252 4752
rect 234 4752 252 4770
rect 234 4770 252 4788
rect 234 4788 252 4806
rect 234 4806 252 4824
rect 234 4824 252 4842
rect 234 4842 252 4860
rect 234 4860 252 4878
rect 234 4878 252 4896
rect 234 4896 252 4914
rect 234 4914 252 4932
rect 252 2286 270 2304
rect 252 2304 270 2322
rect 252 2322 270 2340
rect 252 2340 270 2358
rect 252 2358 270 2376
rect 252 2376 270 2394
rect 252 2394 270 2412
rect 252 2412 270 2430
rect 252 2430 270 2448
rect 252 2448 270 2466
rect 252 2466 270 2484
rect 252 2484 270 2502
rect 252 2502 270 2520
rect 252 2520 270 2538
rect 252 2538 270 2556
rect 252 2556 270 2574
rect 252 2574 270 2592
rect 252 2592 270 2610
rect 252 2610 270 2628
rect 252 2628 270 2646
rect 252 2646 270 2664
rect 252 2664 270 2682
rect 252 2682 270 2700
rect 252 2700 270 2718
rect 252 2718 270 2736
rect 252 2736 270 2754
rect 252 2754 270 2772
rect 252 2772 270 2790
rect 252 2790 270 2808
rect 252 2808 270 2826
rect 252 2826 270 2844
rect 252 2844 270 2862
rect 252 2862 270 2880
rect 252 2880 270 2898
rect 252 2898 270 2916
rect 252 2916 270 2934
rect 252 2934 270 2952
rect 252 2952 270 2970
rect 252 2970 270 2988
rect 252 2988 270 3006
rect 252 3006 270 3024
rect 252 3024 270 3042
rect 252 3042 270 3060
rect 252 3060 270 3078
rect 252 3078 270 3096
rect 252 3096 270 3114
rect 252 3114 270 3132
rect 252 3132 270 3150
rect 252 3150 270 3168
rect 252 3168 270 3186
rect 252 3186 270 3204
rect 252 3204 270 3222
rect 252 3222 270 3240
rect 252 3240 270 3258
rect 252 3258 270 3276
rect 252 3276 270 3294
rect 252 3294 270 3312
rect 252 3312 270 3330
rect 252 3330 270 3348
rect 252 3348 270 3366
rect 252 3366 270 3384
rect 252 3384 270 3402
rect 252 3402 270 3420
rect 252 3420 270 3438
rect 252 3438 270 3456
rect 252 3456 270 3474
rect 252 3474 270 3492
rect 252 3492 270 3510
rect 252 3510 270 3528
rect 252 3528 270 3546
rect 252 3546 270 3564
rect 252 3564 270 3582
rect 252 3582 270 3600
rect 252 3600 270 3618
rect 252 3618 270 3636
rect 252 3636 270 3654
rect 252 3654 270 3672
rect 252 3672 270 3690
rect 252 3690 270 3708
rect 252 3708 270 3726
rect 252 3726 270 3744
rect 252 3744 270 3762
rect 252 3762 270 3780
rect 252 3780 270 3798
rect 252 3798 270 3816
rect 252 3816 270 3834
rect 252 3834 270 3852
rect 252 3852 270 3870
rect 252 3870 270 3888
rect 252 3888 270 3906
rect 252 3906 270 3924
rect 252 3924 270 3942
rect 252 3942 270 3960
rect 252 3960 270 3978
rect 252 3978 270 3996
rect 252 3996 270 4014
rect 252 4014 270 4032
rect 252 4032 270 4050
rect 252 4050 270 4068
rect 252 4068 270 4086
rect 252 4086 270 4104
rect 252 4104 270 4122
rect 252 4122 270 4140
rect 252 4140 270 4158
rect 252 4158 270 4176
rect 252 4176 270 4194
rect 252 4194 270 4212
rect 252 4212 270 4230
rect 252 4230 270 4248
rect 252 4248 270 4266
rect 252 4266 270 4284
rect 252 4284 270 4302
rect 252 4302 270 4320
rect 252 4320 270 4338
rect 252 4338 270 4356
rect 252 4356 270 4374
rect 252 4374 270 4392
rect 252 4392 270 4410
rect 252 4410 270 4428
rect 252 4428 270 4446
rect 252 4446 270 4464
rect 252 4464 270 4482
rect 252 4482 270 4500
rect 252 4500 270 4518
rect 252 4518 270 4536
rect 252 4536 270 4554
rect 252 4554 270 4572
rect 252 4572 270 4590
rect 252 4590 270 4608
rect 252 4608 270 4626
rect 252 4626 270 4644
rect 252 4644 270 4662
rect 252 4662 270 4680
rect 252 4680 270 4698
rect 252 4698 270 4716
rect 252 4716 270 4734
rect 252 4734 270 4752
rect 252 4752 270 4770
rect 252 4770 270 4788
rect 252 4788 270 4806
rect 252 4806 270 4824
rect 252 4824 270 4842
rect 252 4842 270 4860
rect 252 4860 270 4878
rect 252 4878 270 4896
rect 252 4896 270 4914
rect 252 4914 270 4932
rect 252 4932 270 4950
rect 252 4950 270 4968
rect 252 4968 270 4986
rect 270 2250 288 2268
rect 270 2268 288 2286
rect 270 2286 288 2304
rect 270 2304 288 2322
rect 270 2322 288 2340
rect 270 2340 288 2358
rect 270 2358 288 2376
rect 270 2376 288 2394
rect 270 2394 288 2412
rect 270 2412 288 2430
rect 270 2430 288 2448
rect 270 2448 288 2466
rect 270 2466 288 2484
rect 270 2484 288 2502
rect 270 2502 288 2520
rect 270 2520 288 2538
rect 270 2538 288 2556
rect 270 2556 288 2574
rect 270 2574 288 2592
rect 270 2592 288 2610
rect 270 2610 288 2628
rect 270 2628 288 2646
rect 270 2646 288 2664
rect 270 2664 288 2682
rect 270 2682 288 2700
rect 270 2700 288 2718
rect 270 2718 288 2736
rect 270 2736 288 2754
rect 270 2754 288 2772
rect 270 2772 288 2790
rect 270 2790 288 2808
rect 270 2808 288 2826
rect 270 2826 288 2844
rect 270 2844 288 2862
rect 270 2862 288 2880
rect 270 2880 288 2898
rect 270 2898 288 2916
rect 270 2916 288 2934
rect 270 2934 288 2952
rect 270 2952 288 2970
rect 270 2970 288 2988
rect 270 2988 288 3006
rect 270 3006 288 3024
rect 270 3024 288 3042
rect 270 3042 288 3060
rect 270 3060 288 3078
rect 270 3078 288 3096
rect 270 3096 288 3114
rect 270 3114 288 3132
rect 270 3132 288 3150
rect 270 3150 288 3168
rect 270 3168 288 3186
rect 270 3186 288 3204
rect 270 3204 288 3222
rect 270 3222 288 3240
rect 270 3240 288 3258
rect 270 3258 288 3276
rect 270 3276 288 3294
rect 270 3294 288 3312
rect 270 3312 288 3330
rect 270 3330 288 3348
rect 270 3348 288 3366
rect 270 3366 288 3384
rect 270 3384 288 3402
rect 270 3402 288 3420
rect 270 3420 288 3438
rect 270 3438 288 3456
rect 270 3456 288 3474
rect 270 3474 288 3492
rect 270 3492 288 3510
rect 270 3510 288 3528
rect 270 3528 288 3546
rect 270 3546 288 3564
rect 270 3564 288 3582
rect 270 3582 288 3600
rect 270 3600 288 3618
rect 270 3618 288 3636
rect 270 3636 288 3654
rect 270 3654 288 3672
rect 270 3672 288 3690
rect 270 3690 288 3708
rect 270 3708 288 3726
rect 270 3726 288 3744
rect 270 3744 288 3762
rect 270 3762 288 3780
rect 270 3780 288 3798
rect 270 3798 288 3816
rect 270 3816 288 3834
rect 270 3834 288 3852
rect 270 3852 288 3870
rect 270 3870 288 3888
rect 270 3888 288 3906
rect 270 3906 288 3924
rect 270 3924 288 3942
rect 270 3942 288 3960
rect 270 3960 288 3978
rect 270 3978 288 3996
rect 270 3996 288 4014
rect 270 4014 288 4032
rect 270 4032 288 4050
rect 270 4050 288 4068
rect 270 4068 288 4086
rect 270 4086 288 4104
rect 270 4104 288 4122
rect 270 4122 288 4140
rect 270 4140 288 4158
rect 270 4158 288 4176
rect 270 4176 288 4194
rect 270 4194 288 4212
rect 270 4212 288 4230
rect 270 4230 288 4248
rect 270 4248 288 4266
rect 270 4266 288 4284
rect 270 4284 288 4302
rect 270 4302 288 4320
rect 270 4320 288 4338
rect 270 4338 288 4356
rect 270 4356 288 4374
rect 270 4374 288 4392
rect 270 4392 288 4410
rect 270 4410 288 4428
rect 270 4428 288 4446
rect 270 4446 288 4464
rect 270 4464 288 4482
rect 270 4482 288 4500
rect 270 4500 288 4518
rect 270 4518 288 4536
rect 270 4536 288 4554
rect 270 4554 288 4572
rect 270 4572 288 4590
rect 270 4590 288 4608
rect 270 4608 288 4626
rect 270 4626 288 4644
rect 270 4644 288 4662
rect 270 4662 288 4680
rect 270 4680 288 4698
rect 270 4698 288 4716
rect 270 4716 288 4734
rect 270 4734 288 4752
rect 270 4752 288 4770
rect 270 4770 288 4788
rect 270 4788 288 4806
rect 270 4806 288 4824
rect 270 4824 288 4842
rect 270 4842 288 4860
rect 270 4860 288 4878
rect 270 4878 288 4896
rect 270 4896 288 4914
rect 270 4914 288 4932
rect 270 4932 288 4950
rect 270 4950 288 4968
rect 270 4968 288 4986
rect 270 4986 288 5004
rect 270 5004 288 5022
rect 288 2196 306 2214
rect 288 2214 306 2232
rect 288 2232 306 2250
rect 288 2250 306 2268
rect 288 2268 306 2286
rect 288 2286 306 2304
rect 288 2304 306 2322
rect 288 2322 306 2340
rect 288 2340 306 2358
rect 288 2358 306 2376
rect 288 2376 306 2394
rect 288 2394 306 2412
rect 288 2412 306 2430
rect 288 2430 306 2448
rect 288 2448 306 2466
rect 288 2466 306 2484
rect 288 2484 306 2502
rect 288 2502 306 2520
rect 288 2520 306 2538
rect 288 2538 306 2556
rect 288 2556 306 2574
rect 288 2574 306 2592
rect 288 2592 306 2610
rect 288 2610 306 2628
rect 288 2628 306 2646
rect 288 2646 306 2664
rect 288 2664 306 2682
rect 288 2682 306 2700
rect 288 2700 306 2718
rect 288 2718 306 2736
rect 288 2736 306 2754
rect 288 2754 306 2772
rect 288 2772 306 2790
rect 288 2790 306 2808
rect 288 2808 306 2826
rect 288 2826 306 2844
rect 288 2844 306 2862
rect 288 2862 306 2880
rect 288 2880 306 2898
rect 288 2898 306 2916
rect 288 2916 306 2934
rect 288 2934 306 2952
rect 288 2952 306 2970
rect 288 2970 306 2988
rect 288 2988 306 3006
rect 288 3006 306 3024
rect 288 3024 306 3042
rect 288 3042 306 3060
rect 288 3060 306 3078
rect 288 3078 306 3096
rect 288 3096 306 3114
rect 288 3114 306 3132
rect 288 3132 306 3150
rect 288 3150 306 3168
rect 288 3168 306 3186
rect 288 3186 306 3204
rect 288 3204 306 3222
rect 288 3222 306 3240
rect 288 3240 306 3258
rect 288 3258 306 3276
rect 288 3276 306 3294
rect 288 3294 306 3312
rect 288 3312 306 3330
rect 288 3330 306 3348
rect 288 3348 306 3366
rect 288 3366 306 3384
rect 288 3384 306 3402
rect 288 3402 306 3420
rect 288 3420 306 3438
rect 288 3438 306 3456
rect 288 3456 306 3474
rect 288 3474 306 3492
rect 288 3492 306 3510
rect 288 3510 306 3528
rect 288 3528 306 3546
rect 288 3546 306 3564
rect 288 3564 306 3582
rect 288 3582 306 3600
rect 288 3600 306 3618
rect 288 3618 306 3636
rect 288 3636 306 3654
rect 288 3654 306 3672
rect 288 3672 306 3690
rect 288 3690 306 3708
rect 288 3708 306 3726
rect 288 3726 306 3744
rect 288 3744 306 3762
rect 288 3762 306 3780
rect 288 3780 306 3798
rect 288 3798 306 3816
rect 288 3816 306 3834
rect 288 3834 306 3852
rect 288 3852 306 3870
rect 288 3870 306 3888
rect 288 3888 306 3906
rect 288 3906 306 3924
rect 288 3924 306 3942
rect 288 3942 306 3960
rect 288 3960 306 3978
rect 288 3978 306 3996
rect 288 3996 306 4014
rect 288 4014 306 4032
rect 288 4032 306 4050
rect 288 4050 306 4068
rect 288 4068 306 4086
rect 288 4086 306 4104
rect 288 4104 306 4122
rect 288 4122 306 4140
rect 288 4140 306 4158
rect 288 4158 306 4176
rect 288 4176 306 4194
rect 288 4194 306 4212
rect 288 4212 306 4230
rect 288 4230 306 4248
rect 288 4248 306 4266
rect 288 4266 306 4284
rect 288 4284 306 4302
rect 288 4302 306 4320
rect 288 4320 306 4338
rect 288 4338 306 4356
rect 288 4356 306 4374
rect 288 4374 306 4392
rect 288 4392 306 4410
rect 288 4410 306 4428
rect 288 4428 306 4446
rect 288 4446 306 4464
rect 288 4464 306 4482
rect 288 4482 306 4500
rect 288 4500 306 4518
rect 288 4518 306 4536
rect 288 4536 306 4554
rect 288 4554 306 4572
rect 288 4572 306 4590
rect 288 4590 306 4608
rect 288 4608 306 4626
rect 288 4626 306 4644
rect 288 4644 306 4662
rect 288 4662 306 4680
rect 288 4680 306 4698
rect 288 4698 306 4716
rect 288 4716 306 4734
rect 288 4734 306 4752
rect 288 4752 306 4770
rect 288 4770 306 4788
rect 288 4788 306 4806
rect 288 4806 306 4824
rect 288 4824 306 4842
rect 288 4842 306 4860
rect 288 4860 306 4878
rect 288 4878 306 4896
rect 288 4896 306 4914
rect 288 4914 306 4932
rect 288 4932 306 4950
rect 288 4950 306 4968
rect 288 4968 306 4986
rect 288 4986 306 5004
rect 288 5004 306 5022
rect 288 5022 306 5040
rect 288 5040 306 5058
rect 306 2160 324 2178
rect 306 2178 324 2196
rect 306 2196 324 2214
rect 306 2214 324 2232
rect 306 2232 324 2250
rect 306 2250 324 2268
rect 306 2268 324 2286
rect 306 2286 324 2304
rect 306 2304 324 2322
rect 306 2322 324 2340
rect 306 2340 324 2358
rect 306 2358 324 2376
rect 306 2376 324 2394
rect 306 2394 324 2412
rect 306 2412 324 2430
rect 306 2430 324 2448
rect 306 2448 324 2466
rect 306 2466 324 2484
rect 306 2484 324 2502
rect 306 2502 324 2520
rect 306 2520 324 2538
rect 306 2538 324 2556
rect 306 2556 324 2574
rect 306 2574 324 2592
rect 306 2592 324 2610
rect 306 2610 324 2628
rect 306 2628 324 2646
rect 306 2646 324 2664
rect 306 2664 324 2682
rect 306 2682 324 2700
rect 306 2700 324 2718
rect 306 2718 324 2736
rect 306 2736 324 2754
rect 306 2754 324 2772
rect 306 2772 324 2790
rect 306 2790 324 2808
rect 306 2808 324 2826
rect 306 2826 324 2844
rect 306 2844 324 2862
rect 306 2862 324 2880
rect 306 2880 324 2898
rect 306 2898 324 2916
rect 306 2916 324 2934
rect 306 2934 324 2952
rect 306 2952 324 2970
rect 306 2970 324 2988
rect 306 2988 324 3006
rect 306 3006 324 3024
rect 306 3024 324 3042
rect 306 3042 324 3060
rect 306 3060 324 3078
rect 306 3078 324 3096
rect 306 3096 324 3114
rect 306 3114 324 3132
rect 306 3132 324 3150
rect 306 3150 324 3168
rect 306 3168 324 3186
rect 306 3186 324 3204
rect 306 3204 324 3222
rect 306 3222 324 3240
rect 306 3240 324 3258
rect 306 3258 324 3276
rect 306 3276 324 3294
rect 306 3294 324 3312
rect 306 3312 324 3330
rect 306 3330 324 3348
rect 306 3348 324 3366
rect 306 3366 324 3384
rect 306 3384 324 3402
rect 306 3402 324 3420
rect 306 3420 324 3438
rect 306 3438 324 3456
rect 306 3456 324 3474
rect 306 3474 324 3492
rect 306 3492 324 3510
rect 306 3510 324 3528
rect 306 3528 324 3546
rect 306 3546 324 3564
rect 306 3564 324 3582
rect 306 3582 324 3600
rect 306 3600 324 3618
rect 306 3618 324 3636
rect 306 3636 324 3654
rect 306 3654 324 3672
rect 306 3672 324 3690
rect 306 3690 324 3708
rect 306 3708 324 3726
rect 306 3726 324 3744
rect 306 3744 324 3762
rect 306 3762 324 3780
rect 306 3780 324 3798
rect 306 3798 324 3816
rect 306 3816 324 3834
rect 306 3834 324 3852
rect 306 3852 324 3870
rect 306 3870 324 3888
rect 306 3888 324 3906
rect 306 3906 324 3924
rect 306 3924 324 3942
rect 306 3942 324 3960
rect 306 3960 324 3978
rect 306 3978 324 3996
rect 306 3996 324 4014
rect 306 4014 324 4032
rect 306 4032 324 4050
rect 306 4050 324 4068
rect 306 4068 324 4086
rect 306 4086 324 4104
rect 306 4104 324 4122
rect 306 4122 324 4140
rect 306 4140 324 4158
rect 306 4158 324 4176
rect 306 4176 324 4194
rect 306 4194 324 4212
rect 306 4212 324 4230
rect 306 4230 324 4248
rect 306 4248 324 4266
rect 306 4266 324 4284
rect 306 4284 324 4302
rect 306 4302 324 4320
rect 306 4320 324 4338
rect 306 4338 324 4356
rect 306 4356 324 4374
rect 306 4374 324 4392
rect 306 4392 324 4410
rect 306 4410 324 4428
rect 306 4428 324 4446
rect 306 4446 324 4464
rect 306 4464 324 4482
rect 306 4482 324 4500
rect 306 4500 324 4518
rect 306 4518 324 4536
rect 306 4536 324 4554
rect 306 4554 324 4572
rect 306 4572 324 4590
rect 306 4590 324 4608
rect 306 4608 324 4626
rect 306 4626 324 4644
rect 306 4644 324 4662
rect 306 4662 324 4680
rect 306 4680 324 4698
rect 306 4698 324 4716
rect 306 4716 324 4734
rect 306 4734 324 4752
rect 306 4752 324 4770
rect 306 4770 324 4788
rect 306 4788 324 4806
rect 306 4806 324 4824
rect 306 4824 324 4842
rect 306 4842 324 4860
rect 306 4860 324 4878
rect 306 4878 324 4896
rect 306 4896 324 4914
rect 306 4914 324 4932
rect 306 4932 324 4950
rect 306 4950 324 4968
rect 306 4968 324 4986
rect 306 4986 324 5004
rect 306 5004 324 5022
rect 306 5022 324 5040
rect 306 5040 324 5058
rect 306 5058 324 5076
rect 306 5076 324 5094
rect 306 5094 324 5112
rect 324 2124 342 2142
rect 324 2142 342 2160
rect 324 2160 342 2178
rect 324 2178 342 2196
rect 324 2196 342 2214
rect 324 2214 342 2232
rect 324 2232 342 2250
rect 324 2250 342 2268
rect 324 2268 342 2286
rect 324 2286 342 2304
rect 324 2304 342 2322
rect 324 2322 342 2340
rect 324 2340 342 2358
rect 324 2358 342 2376
rect 324 2376 342 2394
rect 324 2394 342 2412
rect 324 2412 342 2430
rect 324 2430 342 2448
rect 324 2448 342 2466
rect 324 2466 342 2484
rect 324 2484 342 2502
rect 324 2502 342 2520
rect 324 2520 342 2538
rect 324 2538 342 2556
rect 324 2556 342 2574
rect 324 2574 342 2592
rect 324 2592 342 2610
rect 324 2610 342 2628
rect 324 2628 342 2646
rect 324 2646 342 2664
rect 324 2664 342 2682
rect 324 2682 342 2700
rect 324 2700 342 2718
rect 324 2718 342 2736
rect 324 2736 342 2754
rect 324 2754 342 2772
rect 324 2772 342 2790
rect 324 2790 342 2808
rect 324 2808 342 2826
rect 324 2826 342 2844
rect 324 2844 342 2862
rect 324 2862 342 2880
rect 324 2880 342 2898
rect 324 2898 342 2916
rect 324 2916 342 2934
rect 324 2934 342 2952
rect 324 2952 342 2970
rect 324 2970 342 2988
rect 324 2988 342 3006
rect 324 3006 342 3024
rect 324 3024 342 3042
rect 324 3042 342 3060
rect 324 3060 342 3078
rect 324 3078 342 3096
rect 324 3096 342 3114
rect 324 3114 342 3132
rect 324 3132 342 3150
rect 324 3150 342 3168
rect 324 3168 342 3186
rect 324 3186 342 3204
rect 324 3204 342 3222
rect 324 3222 342 3240
rect 324 3240 342 3258
rect 324 3258 342 3276
rect 324 3276 342 3294
rect 324 3294 342 3312
rect 324 3312 342 3330
rect 324 3330 342 3348
rect 324 3348 342 3366
rect 324 3366 342 3384
rect 324 3384 342 3402
rect 324 3402 342 3420
rect 324 3420 342 3438
rect 324 3438 342 3456
rect 324 3456 342 3474
rect 324 3474 342 3492
rect 324 3492 342 3510
rect 324 3510 342 3528
rect 324 3528 342 3546
rect 324 3546 342 3564
rect 324 3564 342 3582
rect 324 3582 342 3600
rect 324 3600 342 3618
rect 324 3618 342 3636
rect 324 3636 342 3654
rect 324 3654 342 3672
rect 324 3672 342 3690
rect 324 3690 342 3708
rect 324 3708 342 3726
rect 324 3726 342 3744
rect 324 3744 342 3762
rect 324 3762 342 3780
rect 324 3780 342 3798
rect 324 3798 342 3816
rect 324 3816 342 3834
rect 324 3834 342 3852
rect 324 3852 342 3870
rect 324 3870 342 3888
rect 324 3888 342 3906
rect 324 3906 342 3924
rect 324 3924 342 3942
rect 324 3942 342 3960
rect 324 3960 342 3978
rect 324 3978 342 3996
rect 324 3996 342 4014
rect 324 4014 342 4032
rect 324 4032 342 4050
rect 324 4050 342 4068
rect 324 4068 342 4086
rect 324 4086 342 4104
rect 324 4104 342 4122
rect 324 4122 342 4140
rect 324 4140 342 4158
rect 324 4158 342 4176
rect 324 4176 342 4194
rect 324 4194 342 4212
rect 324 4212 342 4230
rect 324 4230 342 4248
rect 324 4248 342 4266
rect 324 4266 342 4284
rect 324 4284 342 4302
rect 324 4302 342 4320
rect 324 4320 342 4338
rect 324 4338 342 4356
rect 324 4356 342 4374
rect 324 4374 342 4392
rect 324 4392 342 4410
rect 324 4410 342 4428
rect 324 4428 342 4446
rect 324 4446 342 4464
rect 324 4464 342 4482
rect 324 4482 342 4500
rect 324 4500 342 4518
rect 324 4518 342 4536
rect 324 4536 342 4554
rect 324 4554 342 4572
rect 324 4572 342 4590
rect 324 4590 342 4608
rect 324 4608 342 4626
rect 324 4626 342 4644
rect 324 4644 342 4662
rect 324 4662 342 4680
rect 324 4680 342 4698
rect 324 4698 342 4716
rect 324 4716 342 4734
rect 324 4734 342 4752
rect 324 4752 342 4770
rect 324 4770 342 4788
rect 324 4788 342 4806
rect 324 4806 342 4824
rect 324 4824 342 4842
rect 324 4842 342 4860
rect 324 4860 342 4878
rect 324 4878 342 4896
rect 324 4896 342 4914
rect 324 4914 342 4932
rect 324 4932 342 4950
rect 324 4950 342 4968
rect 324 4968 342 4986
rect 324 4986 342 5004
rect 324 5004 342 5022
rect 324 5022 342 5040
rect 324 5040 342 5058
rect 324 5058 342 5076
rect 324 5076 342 5094
rect 324 5094 342 5112
rect 324 5112 342 5130
rect 324 5130 342 5148
rect 342 2088 360 2106
rect 342 2106 360 2124
rect 342 2124 360 2142
rect 342 2142 360 2160
rect 342 2160 360 2178
rect 342 2178 360 2196
rect 342 2196 360 2214
rect 342 2214 360 2232
rect 342 2232 360 2250
rect 342 2250 360 2268
rect 342 2268 360 2286
rect 342 2286 360 2304
rect 342 2304 360 2322
rect 342 2322 360 2340
rect 342 2340 360 2358
rect 342 2358 360 2376
rect 342 2376 360 2394
rect 342 2394 360 2412
rect 342 2412 360 2430
rect 342 2430 360 2448
rect 342 2448 360 2466
rect 342 2466 360 2484
rect 342 2484 360 2502
rect 342 2502 360 2520
rect 342 2520 360 2538
rect 342 2538 360 2556
rect 342 2556 360 2574
rect 342 2574 360 2592
rect 342 2592 360 2610
rect 342 2610 360 2628
rect 342 2628 360 2646
rect 342 2646 360 2664
rect 342 2664 360 2682
rect 342 2682 360 2700
rect 342 2700 360 2718
rect 342 2718 360 2736
rect 342 2736 360 2754
rect 342 2754 360 2772
rect 342 2772 360 2790
rect 342 2790 360 2808
rect 342 2808 360 2826
rect 342 2826 360 2844
rect 342 2844 360 2862
rect 342 2862 360 2880
rect 342 2880 360 2898
rect 342 2898 360 2916
rect 342 2916 360 2934
rect 342 2934 360 2952
rect 342 2952 360 2970
rect 342 2970 360 2988
rect 342 2988 360 3006
rect 342 3006 360 3024
rect 342 3024 360 3042
rect 342 3042 360 3060
rect 342 3060 360 3078
rect 342 3078 360 3096
rect 342 3096 360 3114
rect 342 3114 360 3132
rect 342 3132 360 3150
rect 342 3150 360 3168
rect 342 3168 360 3186
rect 342 3186 360 3204
rect 342 3204 360 3222
rect 342 3222 360 3240
rect 342 3240 360 3258
rect 342 3258 360 3276
rect 342 3276 360 3294
rect 342 3294 360 3312
rect 342 3312 360 3330
rect 342 3330 360 3348
rect 342 3348 360 3366
rect 342 3366 360 3384
rect 342 3384 360 3402
rect 342 3402 360 3420
rect 342 3420 360 3438
rect 342 3438 360 3456
rect 342 3456 360 3474
rect 342 3474 360 3492
rect 342 3492 360 3510
rect 342 3510 360 3528
rect 342 3528 360 3546
rect 342 3546 360 3564
rect 342 3564 360 3582
rect 342 3582 360 3600
rect 342 3600 360 3618
rect 342 3618 360 3636
rect 342 3636 360 3654
rect 342 3654 360 3672
rect 342 3672 360 3690
rect 342 3690 360 3708
rect 342 3708 360 3726
rect 342 3726 360 3744
rect 342 3744 360 3762
rect 342 3762 360 3780
rect 342 3780 360 3798
rect 342 3798 360 3816
rect 342 3816 360 3834
rect 342 3834 360 3852
rect 342 3852 360 3870
rect 342 3870 360 3888
rect 342 3888 360 3906
rect 342 3906 360 3924
rect 342 3924 360 3942
rect 342 3942 360 3960
rect 342 3960 360 3978
rect 342 3978 360 3996
rect 342 3996 360 4014
rect 342 4014 360 4032
rect 342 4032 360 4050
rect 342 4050 360 4068
rect 342 4068 360 4086
rect 342 4086 360 4104
rect 342 4104 360 4122
rect 342 4122 360 4140
rect 342 4140 360 4158
rect 342 4158 360 4176
rect 342 4176 360 4194
rect 342 4194 360 4212
rect 342 4212 360 4230
rect 342 4230 360 4248
rect 342 4248 360 4266
rect 342 4266 360 4284
rect 342 4284 360 4302
rect 342 4302 360 4320
rect 342 4320 360 4338
rect 342 4338 360 4356
rect 342 4356 360 4374
rect 342 4374 360 4392
rect 342 4392 360 4410
rect 342 4410 360 4428
rect 342 4428 360 4446
rect 342 4446 360 4464
rect 342 4464 360 4482
rect 342 4482 360 4500
rect 342 4500 360 4518
rect 342 4518 360 4536
rect 342 4536 360 4554
rect 342 4554 360 4572
rect 342 4572 360 4590
rect 342 4590 360 4608
rect 342 4608 360 4626
rect 342 4626 360 4644
rect 342 4644 360 4662
rect 342 4662 360 4680
rect 342 4680 360 4698
rect 342 4698 360 4716
rect 342 4716 360 4734
rect 342 4734 360 4752
rect 342 4752 360 4770
rect 342 4770 360 4788
rect 342 4788 360 4806
rect 342 4806 360 4824
rect 342 4824 360 4842
rect 342 4842 360 4860
rect 342 4860 360 4878
rect 342 4878 360 4896
rect 342 4896 360 4914
rect 342 4914 360 4932
rect 342 4932 360 4950
rect 342 4950 360 4968
rect 342 4968 360 4986
rect 342 4986 360 5004
rect 342 5004 360 5022
rect 342 5022 360 5040
rect 342 5040 360 5058
rect 342 5058 360 5076
rect 342 5076 360 5094
rect 342 5094 360 5112
rect 342 5112 360 5130
rect 342 5130 360 5148
rect 342 5148 360 5166
rect 342 5166 360 5184
rect 360 2052 378 2070
rect 360 2070 378 2088
rect 360 2088 378 2106
rect 360 2106 378 2124
rect 360 2124 378 2142
rect 360 2142 378 2160
rect 360 2160 378 2178
rect 360 2178 378 2196
rect 360 2196 378 2214
rect 360 2214 378 2232
rect 360 2232 378 2250
rect 360 2250 378 2268
rect 360 2268 378 2286
rect 360 2286 378 2304
rect 360 2304 378 2322
rect 360 2322 378 2340
rect 360 2340 378 2358
rect 360 2358 378 2376
rect 360 2376 378 2394
rect 360 2394 378 2412
rect 360 2412 378 2430
rect 360 2430 378 2448
rect 360 2448 378 2466
rect 360 2466 378 2484
rect 360 2484 378 2502
rect 360 2502 378 2520
rect 360 2520 378 2538
rect 360 2538 378 2556
rect 360 2556 378 2574
rect 360 2574 378 2592
rect 360 2592 378 2610
rect 360 2610 378 2628
rect 360 2628 378 2646
rect 360 2646 378 2664
rect 360 2664 378 2682
rect 360 2682 378 2700
rect 360 2700 378 2718
rect 360 2718 378 2736
rect 360 2736 378 2754
rect 360 2754 378 2772
rect 360 2772 378 2790
rect 360 2790 378 2808
rect 360 2808 378 2826
rect 360 2826 378 2844
rect 360 2844 378 2862
rect 360 2862 378 2880
rect 360 2880 378 2898
rect 360 2898 378 2916
rect 360 2916 378 2934
rect 360 2934 378 2952
rect 360 2952 378 2970
rect 360 2970 378 2988
rect 360 2988 378 3006
rect 360 3006 378 3024
rect 360 3024 378 3042
rect 360 3042 378 3060
rect 360 3060 378 3078
rect 360 3078 378 3096
rect 360 3096 378 3114
rect 360 3114 378 3132
rect 360 3132 378 3150
rect 360 3150 378 3168
rect 360 3168 378 3186
rect 360 3186 378 3204
rect 360 3204 378 3222
rect 360 3222 378 3240
rect 360 3240 378 3258
rect 360 3258 378 3276
rect 360 3276 378 3294
rect 360 3294 378 3312
rect 360 3312 378 3330
rect 360 3330 378 3348
rect 360 3348 378 3366
rect 360 3366 378 3384
rect 360 3384 378 3402
rect 360 3402 378 3420
rect 360 3420 378 3438
rect 360 3438 378 3456
rect 360 3456 378 3474
rect 360 3474 378 3492
rect 360 3492 378 3510
rect 360 3510 378 3528
rect 360 3528 378 3546
rect 360 3546 378 3564
rect 360 3564 378 3582
rect 360 3582 378 3600
rect 360 3600 378 3618
rect 360 3618 378 3636
rect 360 3636 378 3654
rect 360 3654 378 3672
rect 360 3672 378 3690
rect 360 3690 378 3708
rect 360 3708 378 3726
rect 360 3726 378 3744
rect 360 3744 378 3762
rect 360 3762 378 3780
rect 360 3780 378 3798
rect 360 3798 378 3816
rect 360 3816 378 3834
rect 360 3834 378 3852
rect 360 3852 378 3870
rect 360 3870 378 3888
rect 360 3888 378 3906
rect 360 3906 378 3924
rect 360 3924 378 3942
rect 360 3942 378 3960
rect 360 3960 378 3978
rect 360 3978 378 3996
rect 360 3996 378 4014
rect 360 4014 378 4032
rect 360 4032 378 4050
rect 360 4050 378 4068
rect 360 4068 378 4086
rect 360 4086 378 4104
rect 360 4104 378 4122
rect 360 4122 378 4140
rect 360 4140 378 4158
rect 360 4158 378 4176
rect 360 4176 378 4194
rect 360 4194 378 4212
rect 360 4212 378 4230
rect 360 4230 378 4248
rect 360 4248 378 4266
rect 360 4266 378 4284
rect 360 4284 378 4302
rect 360 4302 378 4320
rect 360 4320 378 4338
rect 360 4338 378 4356
rect 360 4356 378 4374
rect 360 4374 378 4392
rect 360 4392 378 4410
rect 360 4410 378 4428
rect 360 4428 378 4446
rect 360 4446 378 4464
rect 360 4464 378 4482
rect 360 4482 378 4500
rect 360 4500 378 4518
rect 360 4518 378 4536
rect 360 4536 378 4554
rect 360 4554 378 4572
rect 360 4572 378 4590
rect 360 4590 378 4608
rect 360 4608 378 4626
rect 360 4626 378 4644
rect 360 4644 378 4662
rect 360 4662 378 4680
rect 360 4680 378 4698
rect 360 4698 378 4716
rect 360 4716 378 4734
rect 360 4734 378 4752
rect 360 4752 378 4770
rect 360 4770 378 4788
rect 360 4788 378 4806
rect 360 4806 378 4824
rect 360 4824 378 4842
rect 360 4842 378 4860
rect 360 4860 378 4878
rect 360 4878 378 4896
rect 360 4896 378 4914
rect 360 4914 378 4932
rect 360 4932 378 4950
rect 360 4950 378 4968
rect 360 4968 378 4986
rect 360 4986 378 5004
rect 360 5004 378 5022
rect 360 5022 378 5040
rect 360 5040 378 5058
rect 360 5058 378 5076
rect 360 5076 378 5094
rect 360 5094 378 5112
rect 360 5112 378 5130
rect 360 5130 378 5148
rect 360 5148 378 5166
rect 360 5166 378 5184
rect 360 5184 378 5202
rect 360 5202 378 5220
rect 378 2016 396 2034
rect 378 2034 396 2052
rect 378 2052 396 2070
rect 378 2070 396 2088
rect 378 2088 396 2106
rect 378 2106 396 2124
rect 378 2124 396 2142
rect 378 2142 396 2160
rect 378 2160 396 2178
rect 378 2178 396 2196
rect 378 2196 396 2214
rect 378 2214 396 2232
rect 378 2232 396 2250
rect 378 2250 396 2268
rect 378 2268 396 2286
rect 378 2286 396 2304
rect 378 2304 396 2322
rect 378 2322 396 2340
rect 378 2340 396 2358
rect 378 2358 396 2376
rect 378 2376 396 2394
rect 378 2394 396 2412
rect 378 2412 396 2430
rect 378 2430 396 2448
rect 378 2448 396 2466
rect 378 2466 396 2484
rect 378 2484 396 2502
rect 378 2502 396 2520
rect 378 2520 396 2538
rect 378 2538 396 2556
rect 378 2556 396 2574
rect 378 2574 396 2592
rect 378 2592 396 2610
rect 378 2610 396 2628
rect 378 2628 396 2646
rect 378 2646 396 2664
rect 378 2664 396 2682
rect 378 2682 396 2700
rect 378 2700 396 2718
rect 378 2718 396 2736
rect 378 2736 396 2754
rect 378 2754 396 2772
rect 378 2772 396 2790
rect 378 2790 396 2808
rect 378 2808 396 2826
rect 378 2826 396 2844
rect 378 2844 396 2862
rect 378 2862 396 2880
rect 378 2880 396 2898
rect 378 2898 396 2916
rect 378 2916 396 2934
rect 378 2934 396 2952
rect 378 2952 396 2970
rect 378 2970 396 2988
rect 378 2988 396 3006
rect 378 3006 396 3024
rect 378 3024 396 3042
rect 378 3042 396 3060
rect 378 3060 396 3078
rect 378 3078 396 3096
rect 378 3096 396 3114
rect 378 3114 396 3132
rect 378 3132 396 3150
rect 378 3150 396 3168
rect 378 3168 396 3186
rect 378 3186 396 3204
rect 378 3204 396 3222
rect 378 3222 396 3240
rect 378 3240 396 3258
rect 378 3258 396 3276
rect 378 3276 396 3294
rect 378 3294 396 3312
rect 378 3312 396 3330
rect 378 3330 396 3348
rect 378 3348 396 3366
rect 378 3366 396 3384
rect 378 3384 396 3402
rect 378 3402 396 3420
rect 378 3420 396 3438
rect 378 3438 396 3456
rect 378 3456 396 3474
rect 378 3474 396 3492
rect 378 3492 396 3510
rect 378 3510 396 3528
rect 378 3528 396 3546
rect 378 3546 396 3564
rect 378 3564 396 3582
rect 378 3582 396 3600
rect 378 3600 396 3618
rect 378 3618 396 3636
rect 378 3636 396 3654
rect 378 3654 396 3672
rect 378 3672 396 3690
rect 378 3690 396 3708
rect 378 3708 396 3726
rect 378 3726 396 3744
rect 378 3744 396 3762
rect 378 3762 396 3780
rect 378 3780 396 3798
rect 378 3798 396 3816
rect 378 3816 396 3834
rect 378 3834 396 3852
rect 378 3852 396 3870
rect 378 3870 396 3888
rect 378 3888 396 3906
rect 378 3906 396 3924
rect 378 3924 396 3942
rect 378 3942 396 3960
rect 378 3960 396 3978
rect 378 3978 396 3996
rect 378 3996 396 4014
rect 378 4014 396 4032
rect 378 4032 396 4050
rect 378 4050 396 4068
rect 378 4068 396 4086
rect 378 4086 396 4104
rect 378 4104 396 4122
rect 378 4122 396 4140
rect 378 4140 396 4158
rect 378 4158 396 4176
rect 378 4176 396 4194
rect 378 4194 396 4212
rect 378 4212 396 4230
rect 378 4230 396 4248
rect 378 4248 396 4266
rect 378 4266 396 4284
rect 378 4284 396 4302
rect 378 4302 396 4320
rect 378 4320 396 4338
rect 378 4338 396 4356
rect 378 4356 396 4374
rect 378 4374 396 4392
rect 378 4392 396 4410
rect 378 4410 396 4428
rect 378 4428 396 4446
rect 378 4446 396 4464
rect 378 4464 396 4482
rect 378 4482 396 4500
rect 378 4500 396 4518
rect 378 4518 396 4536
rect 378 4536 396 4554
rect 378 4554 396 4572
rect 378 4572 396 4590
rect 378 4590 396 4608
rect 378 4608 396 4626
rect 378 4626 396 4644
rect 378 4644 396 4662
rect 378 4662 396 4680
rect 378 4680 396 4698
rect 378 4698 396 4716
rect 378 4716 396 4734
rect 378 4734 396 4752
rect 378 4752 396 4770
rect 378 4770 396 4788
rect 378 4788 396 4806
rect 378 4806 396 4824
rect 378 4824 396 4842
rect 378 4842 396 4860
rect 378 4860 396 4878
rect 378 4878 396 4896
rect 378 4896 396 4914
rect 378 4914 396 4932
rect 378 4932 396 4950
rect 378 4950 396 4968
rect 378 4968 396 4986
rect 378 4986 396 5004
rect 378 5004 396 5022
rect 378 5022 396 5040
rect 378 5040 396 5058
rect 378 5058 396 5076
rect 378 5076 396 5094
rect 378 5094 396 5112
rect 378 5112 396 5130
rect 378 5130 396 5148
rect 378 5148 396 5166
rect 378 5166 396 5184
rect 378 5184 396 5202
rect 378 5202 396 5220
rect 378 5220 396 5238
rect 378 5238 396 5256
rect 396 1980 414 1998
rect 396 1998 414 2016
rect 396 2016 414 2034
rect 396 2034 414 2052
rect 396 2052 414 2070
rect 396 2070 414 2088
rect 396 2088 414 2106
rect 396 2106 414 2124
rect 396 2124 414 2142
rect 396 2142 414 2160
rect 396 2160 414 2178
rect 396 2178 414 2196
rect 396 2196 414 2214
rect 396 2214 414 2232
rect 396 2232 414 2250
rect 396 2250 414 2268
rect 396 2268 414 2286
rect 396 2286 414 2304
rect 396 2304 414 2322
rect 396 2322 414 2340
rect 396 2340 414 2358
rect 396 2358 414 2376
rect 396 2376 414 2394
rect 396 2394 414 2412
rect 396 2412 414 2430
rect 396 2430 414 2448
rect 396 2448 414 2466
rect 396 2466 414 2484
rect 396 2484 414 2502
rect 396 2502 414 2520
rect 396 2520 414 2538
rect 396 2538 414 2556
rect 396 2556 414 2574
rect 396 2574 414 2592
rect 396 2592 414 2610
rect 396 2610 414 2628
rect 396 2628 414 2646
rect 396 2646 414 2664
rect 396 2664 414 2682
rect 396 2682 414 2700
rect 396 2700 414 2718
rect 396 2718 414 2736
rect 396 2736 414 2754
rect 396 2754 414 2772
rect 396 2772 414 2790
rect 396 2790 414 2808
rect 396 2808 414 2826
rect 396 2826 414 2844
rect 396 2844 414 2862
rect 396 2862 414 2880
rect 396 2880 414 2898
rect 396 2898 414 2916
rect 396 2916 414 2934
rect 396 2934 414 2952
rect 396 2952 414 2970
rect 396 2970 414 2988
rect 396 2988 414 3006
rect 396 3006 414 3024
rect 396 3024 414 3042
rect 396 3042 414 3060
rect 396 3060 414 3078
rect 396 3078 414 3096
rect 396 3096 414 3114
rect 396 3114 414 3132
rect 396 3132 414 3150
rect 396 3150 414 3168
rect 396 3168 414 3186
rect 396 3186 414 3204
rect 396 3204 414 3222
rect 396 3222 414 3240
rect 396 3240 414 3258
rect 396 3258 414 3276
rect 396 3276 414 3294
rect 396 3294 414 3312
rect 396 3312 414 3330
rect 396 3330 414 3348
rect 396 3348 414 3366
rect 396 3366 414 3384
rect 396 3384 414 3402
rect 396 3402 414 3420
rect 396 3420 414 3438
rect 396 3438 414 3456
rect 396 3456 414 3474
rect 396 3474 414 3492
rect 396 3492 414 3510
rect 396 3510 414 3528
rect 396 3528 414 3546
rect 396 3546 414 3564
rect 396 3564 414 3582
rect 396 3582 414 3600
rect 396 3600 414 3618
rect 396 3618 414 3636
rect 396 3636 414 3654
rect 396 3654 414 3672
rect 396 3672 414 3690
rect 396 3690 414 3708
rect 396 3708 414 3726
rect 396 3726 414 3744
rect 396 3744 414 3762
rect 396 3762 414 3780
rect 396 3780 414 3798
rect 396 3798 414 3816
rect 396 3816 414 3834
rect 396 3834 414 3852
rect 396 3852 414 3870
rect 396 3870 414 3888
rect 396 3888 414 3906
rect 396 3906 414 3924
rect 396 3924 414 3942
rect 396 3942 414 3960
rect 396 3960 414 3978
rect 396 3978 414 3996
rect 396 3996 414 4014
rect 396 4014 414 4032
rect 396 4032 414 4050
rect 396 4050 414 4068
rect 396 4068 414 4086
rect 396 4086 414 4104
rect 396 4104 414 4122
rect 396 4122 414 4140
rect 396 4140 414 4158
rect 396 4158 414 4176
rect 396 4176 414 4194
rect 396 4194 414 4212
rect 396 4212 414 4230
rect 396 4230 414 4248
rect 396 4248 414 4266
rect 396 4266 414 4284
rect 396 4284 414 4302
rect 396 4302 414 4320
rect 396 4320 414 4338
rect 396 4338 414 4356
rect 396 4356 414 4374
rect 396 4374 414 4392
rect 396 4392 414 4410
rect 396 4410 414 4428
rect 396 4428 414 4446
rect 396 4446 414 4464
rect 396 4464 414 4482
rect 396 4482 414 4500
rect 396 4500 414 4518
rect 396 4518 414 4536
rect 396 4536 414 4554
rect 396 4554 414 4572
rect 396 4572 414 4590
rect 396 4590 414 4608
rect 396 4608 414 4626
rect 396 4626 414 4644
rect 396 4644 414 4662
rect 396 4662 414 4680
rect 396 4680 414 4698
rect 396 4698 414 4716
rect 396 4716 414 4734
rect 396 4734 414 4752
rect 396 4752 414 4770
rect 396 4770 414 4788
rect 396 4788 414 4806
rect 396 4806 414 4824
rect 396 4824 414 4842
rect 396 4842 414 4860
rect 396 4860 414 4878
rect 396 4878 414 4896
rect 396 4896 414 4914
rect 396 4914 414 4932
rect 396 4932 414 4950
rect 396 4950 414 4968
rect 396 4968 414 4986
rect 396 4986 414 5004
rect 396 5004 414 5022
rect 396 5022 414 5040
rect 396 5040 414 5058
rect 396 5058 414 5076
rect 396 5076 414 5094
rect 396 5094 414 5112
rect 396 5112 414 5130
rect 396 5130 414 5148
rect 396 5148 414 5166
rect 396 5166 414 5184
rect 396 5184 414 5202
rect 396 5202 414 5220
rect 396 5220 414 5238
rect 396 5238 414 5256
rect 396 5256 414 5274
rect 396 5274 414 5292
rect 414 1944 432 1962
rect 414 1962 432 1980
rect 414 1980 432 1998
rect 414 1998 432 2016
rect 414 2016 432 2034
rect 414 2034 432 2052
rect 414 2052 432 2070
rect 414 2070 432 2088
rect 414 2088 432 2106
rect 414 2106 432 2124
rect 414 2124 432 2142
rect 414 2142 432 2160
rect 414 2160 432 2178
rect 414 2178 432 2196
rect 414 2196 432 2214
rect 414 2214 432 2232
rect 414 2232 432 2250
rect 414 2250 432 2268
rect 414 2268 432 2286
rect 414 2286 432 2304
rect 414 2304 432 2322
rect 414 2322 432 2340
rect 414 2340 432 2358
rect 414 2358 432 2376
rect 414 2376 432 2394
rect 414 2394 432 2412
rect 414 2412 432 2430
rect 414 2430 432 2448
rect 414 2448 432 2466
rect 414 2466 432 2484
rect 414 2484 432 2502
rect 414 2502 432 2520
rect 414 2520 432 2538
rect 414 2538 432 2556
rect 414 2556 432 2574
rect 414 2574 432 2592
rect 414 2592 432 2610
rect 414 2610 432 2628
rect 414 2628 432 2646
rect 414 2646 432 2664
rect 414 2664 432 2682
rect 414 2682 432 2700
rect 414 2700 432 2718
rect 414 2718 432 2736
rect 414 2736 432 2754
rect 414 2754 432 2772
rect 414 2772 432 2790
rect 414 2790 432 2808
rect 414 2808 432 2826
rect 414 2826 432 2844
rect 414 2844 432 2862
rect 414 2862 432 2880
rect 414 2880 432 2898
rect 414 2898 432 2916
rect 414 2916 432 2934
rect 414 2934 432 2952
rect 414 2952 432 2970
rect 414 2970 432 2988
rect 414 2988 432 3006
rect 414 3006 432 3024
rect 414 3024 432 3042
rect 414 3042 432 3060
rect 414 3060 432 3078
rect 414 3078 432 3096
rect 414 3096 432 3114
rect 414 3114 432 3132
rect 414 3132 432 3150
rect 414 3150 432 3168
rect 414 3168 432 3186
rect 414 3186 432 3204
rect 414 3204 432 3222
rect 414 3222 432 3240
rect 414 3240 432 3258
rect 414 3258 432 3276
rect 414 3276 432 3294
rect 414 3294 432 3312
rect 414 3312 432 3330
rect 414 3330 432 3348
rect 414 3348 432 3366
rect 414 3366 432 3384
rect 414 3384 432 3402
rect 414 3402 432 3420
rect 414 3420 432 3438
rect 414 3438 432 3456
rect 414 3456 432 3474
rect 414 3474 432 3492
rect 414 3492 432 3510
rect 414 3510 432 3528
rect 414 3528 432 3546
rect 414 3546 432 3564
rect 414 3564 432 3582
rect 414 3582 432 3600
rect 414 3600 432 3618
rect 414 3618 432 3636
rect 414 3636 432 3654
rect 414 3654 432 3672
rect 414 3672 432 3690
rect 414 3690 432 3708
rect 414 3708 432 3726
rect 414 3726 432 3744
rect 414 3744 432 3762
rect 414 3762 432 3780
rect 414 3780 432 3798
rect 414 3798 432 3816
rect 414 3816 432 3834
rect 414 3834 432 3852
rect 414 3852 432 3870
rect 414 3870 432 3888
rect 414 3888 432 3906
rect 414 3906 432 3924
rect 414 3924 432 3942
rect 414 3942 432 3960
rect 414 3960 432 3978
rect 414 3978 432 3996
rect 414 3996 432 4014
rect 414 4014 432 4032
rect 414 4032 432 4050
rect 414 4050 432 4068
rect 414 4068 432 4086
rect 414 4086 432 4104
rect 414 4104 432 4122
rect 414 4122 432 4140
rect 414 4140 432 4158
rect 414 4158 432 4176
rect 414 4176 432 4194
rect 414 4194 432 4212
rect 414 4212 432 4230
rect 414 4230 432 4248
rect 414 4248 432 4266
rect 414 4266 432 4284
rect 414 4284 432 4302
rect 414 4302 432 4320
rect 414 4320 432 4338
rect 414 4338 432 4356
rect 414 4356 432 4374
rect 414 4374 432 4392
rect 414 4392 432 4410
rect 414 4410 432 4428
rect 414 4428 432 4446
rect 414 4446 432 4464
rect 414 4464 432 4482
rect 414 4482 432 4500
rect 414 4500 432 4518
rect 414 4518 432 4536
rect 414 4536 432 4554
rect 414 4554 432 4572
rect 414 4572 432 4590
rect 414 4590 432 4608
rect 414 4608 432 4626
rect 414 4626 432 4644
rect 414 4644 432 4662
rect 414 4662 432 4680
rect 414 4680 432 4698
rect 414 4698 432 4716
rect 414 4716 432 4734
rect 414 4734 432 4752
rect 414 4752 432 4770
rect 414 4770 432 4788
rect 414 4788 432 4806
rect 414 4806 432 4824
rect 414 4824 432 4842
rect 414 4842 432 4860
rect 414 4860 432 4878
rect 414 4878 432 4896
rect 414 4896 432 4914
rect 414 4914 432 4932
rect 414 4932 432 4950
rect 414 4950 432 4968
rect 414 4968 432 4986
rect 414 4986 432 5004
rect 414 5004 432 5022
rect 414 5022 432 5040
rect 414 5040 432 5058
rect 414 5058 432 5076
rect 414 5076 432 5094
rect 414 5094 432 5112
rect 414 5112 432 5130
rect 414 5130 432 5148
rect 414 5148 432 5166
rect 414 5166 432 5184
rect 414 5184 432 5202
rect 414 5202 432 5220
rect 414 5220 432 5238
rect 414 5238 432 5256
rect 414 5256 432 5274
rect 414 5274 432 5292
rect 414 5292 432 5310
rect 414 5310 432 5328
rect 432 1908 450 1926
rect 432 1926 450 1944
rect 432 1944 450 1962
rect 432 1962 450 1980
rect 432 1980 450 1998
rect 432 1998 450 2016
rect 432 2016 450 2034
rect 432 2034 450 2052
rect 432 2052 450 2070
rect 432 2070 450 2088
rect 432 2088 450 2106
rect 432 2106 450 2124
rect 432 2124 450 2142
rect 432 2142 450 2160
rect 432 2160 450 2178
rect 432 2178 450 2196
rect 432 2196 450 2214
rect 432 2214 450 2232
rect 432 2232 450 2250
rect 432 2250 450 2268
rect 432 2268 450 2286
rect 432 2286 450 2304
rect 432 2304 450 2322
rect 432 2322 450 2340
rect 432 2340 450 2358
rect 432 2358 450 2376
rect 432 2376 450 2394
rect 432 2394 450 2412
rect 432 2412 450 2430
rect 432 2430 450 2448
rect 432 2448 450 2466
rect 432 2466 450 2484
rect 432 2484 450 2502
rect 432 2502 450 2520
rect 432 2520 450 2538
rect 432 2538 450 2556
rect 432 2556 450 2574
rect 432 2574 450 2592
rect 432 2592 450 2610
rect 432 2610 450 2628
rect 432 2628 450 2646
rect 432 2646 450 2664
rect 432 2664 450 2682
rect 432 2682 450 2700
rect 432 2700 450 2718
rect 432 2718 450 2736
rect 432 2736 450 2754
rect 432 2754 450 2772
rect 432 2772 450 2790
rect 432 2790 450 2808
rect 432 2808 450 2826
rect 432 2826 450 2844
rect 432 2844 450 2862
rect 432 2862 450 2880
rect 432 2880 450 2898
rect 432 2898 450 2916
rect 432 2916 450 2934
rect 432 2934 450 2952
rect 432 2952 450 2970
rect 432 2970 450 2988
rect 432 2988 450 3006
rect 432 3006 450 3024
rect 432 3024 450 3042
rect 432 3042 450 3060
rect 432 3060 450 3078
rect 432 3078 450 3096
rect 432 3096 450 3114
rect 432 3114 450 3132
rect 432 3132 450 3150
rect 432 3150 450 3168
rect 432 3168 450 3186
rect 432 3186 450 3204
rect 432 3204 450 3222
rect 432 3222 450 3240
rect 432 3240 450 3258
rect 432 3258 450 3276
rect 432 3276 450 3294
rect 432 3294 450 3312
rect 432 3312 450 3330
rect 432 3330 450 3348
rect 432 3348 450 3366
rect 432 3366 450 3384
rect 432 3384 450 3402
rect 432 3402 450 3420
rect 432 3420 450 3438
rect 432 3438 450 3456
rect 432 3456 450 3474
rect 432 3474 450 3492
rect 432 3492 450 3510
rect 432 3510 450 3528
rect 432 3528 450 3546
rect 432 3546 450 3564
rect 432 3564 450 3582
rect 432 3582 450 3600
rect 432 3600 450 3618
rect 432 3618 450 3636
rect 432 3636 450 3654
rect 432 3654 450 3672
rect 432 3672 450 3690
rect 432 3690 450 3708
rect 432 3708 450 3726
rect 432 3726 450 3744
rect 432 3744 450 3762
rect 432 3762 450 3780
rect 432 3780 450 3798
rect 432 3798 450 3816
rect 432 3816 450 3834
rect 432 3834 450 3852
rect 432 3852 450 3870
rect 432 3870 450 3888
rect 432 3888 450 3906
rect 432 3906 450 3924
rect 432 3924 450 3942
rect 432 3942 450 3960
rect 432 3960 450 3978
rect 432 3978 450 3996
rect 432 3996 450 4014
rect 432 4014 450 4032
rect 432 4032 450 4050
rect 432 4050 450 4068
rect 432 4068 450 4086
rect 432 4086 450 4104
rect 432 4104 450 4122
rect 432 4122 450 4140
rect 432 4140 450 4158
rect 432 4158 450 4176
rect 432 4176 450 4194
rect 432 4194 450 4212
rect 432 4212 450 4230
rect 432 4230 450 4248
rect 432 4248 450 4266
rect 432 4266 450 4284
rect 432 4284 450 4302
rect 432 4302 450 4320
rect 432 4320 450 4338
rect 432 4338 450 4356
rect 432 4356 450 4374
rect 432 4374 450 4392
rect 432 4392 450 4410
rect 432 4410 450 4428
rect 432 4428 450 4446
rect 432 4446 450 4464
rect 432 4464 450 4482
rect 432 4482 450 4500
rect 432 4500 450 4518
rect 432 4518 450 4536
rect 432 4536 450 4554
rect 432 4554 450 4572
rect 432 4572 450 4590
rect 432 4590 450 4608
rect 432 4608 450 4626
rect 432 4626 450 4644
rect 432 4644 450 4662
rect 432 4662 450 4680
rect 432 4680 450 4698
rect 432 4698 450 4716
rect 432 4716 450 4734
rect 432 4734 450 4752
rect 432 4752 450 4770
rect 432 4770 450 4788
rect 432 4788 450 4806
rect 432 4806 450 4824
rect 432 4824 450 4842
rect 432 4842 450 4860
rect 432 4860 450 4878
rect 432 4878 450 4896
rect 432 4896 450 4914
rect 432 4914 450 4932
rect 432 4932 450 4950
rect 432 4950 450 4968
rect 432 4968 450 4986
rect 432 4986 450 5004
rect 432 5004 450 5022
rect 432 5022 450 5040
rect 432 5040 450 5058
rect 432 5058 450 5076
rect 432 5076 450 5094
rect 432 5094 450 5112
rect 432 5112 450 5130
rect 432 5130 450 5148
rect 432 5148 450 5166
rect 432 5166 450 5184
rect 432 5184 450 5202
rect 432 5202 450 5220
rect 432 5220 450 5238
rect 432 5238 450 5256
rect 432 5256 450 5274
rect 432 5274 450 5292
rect 432 5292 450 5310
rect 432 5310 450 5328
rect 432 5328 450 5346
rect 432 5346 450 5364
rect 450 1872 468 1890
rect 450 1890 468 1908
rect 450 1908 468 1926
rect 450 1926 468 1944
rect 450 1944 468 1962
rect 450 1962 468 1980
rect 450 1980 468 1998
rect 450 1998 468 2016
rect 450 2016 468 2034
rect 450 2034 468 2052
rect 450 2052 468 2070
rect 450 2070 468 2088
rect 450 2088 468 2106
rect 450 2106 468 2124
rect 450 2124 468 2142
rect 450 2142 468 2160
rect 450 2160 468 2178
rect 450 2178 468 2196
rect 450 2196 468 2214
rect 450 2214 468 2232
rect 450 2232 468 2250
rect 450 2250 468 2268
rect 450 2268 468 2286
rect 450 2286 468 2304
rect 450 2304 468 2322
rect 450 2322 468 2340
rect 450 2340 468 2358
rect 450 2358 468 2376
rect 450 2376 468 2394
rect 450 2394 468 2412
rect 450 2412 468 2430
rect 450 2430 468 2448
rect 450 2448 468 2466
rect 450 2466 468 2484
rect 450 2484 468 2502
rect 450 2502 468 2520
rect 450 2520 468 2538
rect 450 2538 468 2556
rect 450 2556 468 2574
rect 450 2574 468 2592
rect 450 2592 468 2610
rect 450 2610 468 2628
rect 450 2628 468 2646
rect 450 2646 468 2664
rect 450 2664 468 2682
rect 450 2682 468 2700
rect 450 2700 468 2718
rect 450 2718 468 2736
rect 450 2736 468 2754
rect 450 2754 468 2772
rect 450 2772 468 2790
rect 450 2790 468 2808
rect 450 2808 468 2826
rect 450 2826 468 2844
rect 450 2844 468 2862
rect 450 2862 468 2880
rect 450 2880 468 2898
rect 450 2898 468 2916
rect 450 2916 468 2934
rect 450 2934 468 2952
rect 450 2952 468 2970
rect 450 2970 468 2988
rect 450 2988 468 3006
rect 450 3006 468 3024
rect 450 3024 468 3042
rect 450 3042 468 3060
rect 450 3060 468 3078
rect 450 3078 468 3096
rect 450 3096 468 3114
rect 450 3114 468 3132
rect 450 3132 468 3150
rect 450 3150 468 3168
rect 450 3168 468 3186
rect 450 3186 468 3204
rect 450 3204 468 3222
rect 450 3222 468 3240
rect 450 3240 468 3258
rect 450 3258 468 3276
rect 450 3276 468 3294
rect 450 3294 468 3312
rect 450 3312 468 3330
rect 450 3330 468 3348
rect 450 3348 468 3366
rect 450 3366 468 3384
rect 450 3384 468 3402
rect 450 3402 468 3420
rect 450 3420 468 3438
rect 450 3438 468 3456
rect 450 3456 468 3474
rect 450 3474 468 3492
rect 450 3492 468 3510
rect 450 3510 468 3528
rect 450 3528 468 3546
rect 450 3546 468 3564
rect 450 3564 468 3582
rect 450 3582 468 3600
rect 450 3600 468 3618
rect 450 3618 468 3636
rect 450 3636 468 3654
rect 450 3654 468 3672
rect 450 3672 468 3690
rect 450 3690 468 3708
rect 450 3708 468 3726
rect 450 3726 468 3744
rect 450 3744 468 3762
rect 450 3762 468 3780
rect 450 3780 468 3798
rect 450 3798 468 3816
rect 450 3816 468 3834
rect 450 3834 468 3852
rect 450 3852 468 3870
rect 450 3870 468 3888
rect 450 3888 468 3906
rect 450 3906 468 3924
rect 450 3924 468 3942
rect 450 3942 468 3960
rect 450 3960 468 3978
rect 450 3978 468 3996
rect 450 3996 468 4014
rect 450 4014 468 4032
rect 450 4032 468 4050
rect 450 4050 468 4068
rect 450 4068 468 4086
rect 450 4086 468 4104
rect 450 4104 468 4122
rect 450 4122 468 4140
rect 450 4140 468 4158
rect 450 4158 468 4176
rect 450 4176 468 4194
rect 450 4194 468 4212
rect 450 4212 468 4230
rect 450 4230 468 4248
rect 450 4248 468 4266
rect 450 4266 468 4284
rect 450 4284 468 4302
rect 450 4302 468 4320
rect 450 4320 468 4338
rect 450 4338 468 4356
rect 450 4356 468 4374
rect 450 4374 468 4392
rect 450 4392 468 4410
rect 450 4410 468 4428
rect 450 4428 468 4446
rect 450 4446 468 4464
rect 450 4464 468 4482
rect 450 4482 468 4500
rect 450 4500 468 4518
rect 450 4518 468 4536
rect 450 4536 468 4554
rect 450 4554 468 4572
rect 450 4572 468 4590
rect 450 4590 468 4608
rect 450 4608 468 4626
rect 450 4626 468 4644
rect 450 4644 468 4662
rect 450 4662 468 4680
rect 450 4680 468 4698
rect 450 4698 468 4716
rect 450 4716 468 4734
rect 450 4734 468 4752
rect 450 4752 468 4770
rect 450 4770 468 4788
rect 450 4788 468 4806
rect 450 4806 468 4824
rect 450 4824 468 4842
rect 450 4842 468 4860
rect 450 4860 468 4878
rect 450 4878 468 4896
rect 450 4896 468 4914
rect 450 4914 468 4932
rect 450 4932 468 4950
rect 450 4950 468 4968
rect 450 4968 468 4986
rect 450 4986 468 5004
rect 450 5004 468 5022
rect 450 5022 468 5040
rect 450 5040 468 5058
rect 450 5058 468 5076
rect 450 5076 468 5094
rect 450 5094 468 5112
rect 450 5112 468 5130
rect 450 5130 468 5148
rect 450 5148 468 5166
rect 450 5166 468 5184
rect 450 5184 468 5202
rect 450 5202 468 5220
rect 450 5220 468 5238
rect 450 5238 468 5256
rect 450 5256 468 5274
rect 450 5274 468 5292
rect 450 5292 468 5310
rect 450 5310 468 5328
rect 450 5328 468 5346
rect 450 5346 468 5364
rect 450 5364 468 5382
rect 450 5382 468 5400
rect 468 1836 486 1854
rect 468 1854 486 1872
rect 468 1872 486 1890
rect 468 1890 486 1908
rect 468 1908 486 1926
rect 468 1926 486 1944
rect 468 1944 486 1962
rect 468 1962 486 1980
rect 468 1980 486 1998
rect 468 1998 486 2016
rect 468 2016 486 2034
rect 468 2034 486 2052
rect 468 2052 486 2070
rect 468 2070 486 2088
rect 468 2088 486 2106
rect 468 2106 486 2124
rect 468 2124 486 2142
rect 468 2142 486 2160
rect 468 2160 486 2178
rect 468 2178 486 2196
rect 468 2196 486 2214
rect 468 2214 486 2232
rect 468 2232 486 2250
rect 468 2250 486 2268
rect 468 2268 486 2286
rect 468 2286 486 2304
rect 468 2304 486 2322
rect 468 2322 486 2340
rect 468 2340 486 2358
rect 468 2358 486 2376
rect 468 2376 486 2394
rect 468 2394 486 2412
rect 468 2412 486 2430
rect 468 2430 486 2448
rect 468 2448 486 2466
rect 468 2466 486 2484
rect 468 2484 486 2502
rect 468 2502 486 2520
rect 468 2520 486 2538
rect 468 2538 486 2556
rect 468 2556 486 2574
rect 468 2574 486 2592
rect 468 2592 486 2610
rect 468 2610 486 2628
rect 468 2628 486 2646
rect 468 2646 486 2664
rect 468 2664 486 2682
rect 468 2682 486 2700
rect 468 2700 486 2718
rect 468 2718 486 2736
rect 468 2736 486 2754
rect 468 2754 486 2772
rect 468 2772 486 2790
rect 468 2790 486 2808
rect 468 2808 486 2826
rect 468 2826 486 2844
rect 468 2844 486 2862
rect 468 2862 486 2880
rect 468 2880 486 2898
rect 468 2898 486 2916
rect 468 2916 486 2934
rect 468 2934 486 2952
rect 468 2952 486 2970
rect 468 2970 486 2988
rect 468 2988 486 3006
rect 468 3006 486 3024
rect 468 3024 486 3042
rect 468 3042 486 3060
rect 468 3060 486 3078
rect 468 3078 486 3096
rect 468 3096 486 3114
rect 468 3114 486 3132
rect 468 3132 486 3150
rect 468 3150 486 3168
rect 468 3168 486 3186
rect 468 3186 486 3204
rect 468 3204 486 3222
rect 468 3222 486 3240
rect 468 3240 486 3258
rect 468 3258 486 3276
rect 468 3276 486 3294
rect 468 3294 486 3312
rect 468 3312 486 3330
rect 468 3330 486 3348
rect 468 3348 486 3366
rect 468 3366 486 3384
rect 468 3384 486 3402
rect 468 3402 486 3420
rect 468 3420 486 3438
rect 468 3438 486 3456
rect 468 3456 486 3474
rect 468 3474 486 3492
rect 468 3492 486 3510
rect 468 3510 486 3528
rect 468 3528 486 3546
rect 468 3546 486 3564
rect 468 3564 486 3582
rect 468 3582 486 3600
rect 468 3600 486 3618
rect 468 3618 486 3636
rect 468 3636 486 3654
rect 468 3654 486 3672
rect 468 3672 486 3690
rect 468 3690 486 3708
rect 468 3708 486 3726
rect 468 3726 486 3744
rect 468 3744 486 3762
rect 468 3762 486 3780
rect 468 3780 486 3798
rect 468 3798 486 3816
rect 468 3816 486 3834
rect 468 3834 486 3852
rect 468 3852 486 3870
rect 468 3870 486 3888
rect 468 3888 486 3906
rect 468 3906 486 3924
rect 468 3924 486 3942
rect 468 3942 486 3960
rect 468 3960 486 3978
rect 468 3978 486 3996
rect 468 3996 486 4014
rect 468 4014 486 4032
rect 468 4032 486 4050
rect 468 4050 486 4068
rect 468 4068 486 4086
rect 468 4086 486 4104
rect 468 4104 486 4122
rect 468 4122 486 4140
rect 468 4140 486 4158
rect 468 4158 486 4176
rect 468 4176 486 4194
rect 468 4194 486 4212
rect 468 4212 486 4230
rect 468 4230 486 4248
rect 468 4248 486 4266
rect 468 4266 486 4284
rect 468 4284 486 4302
rect 468 4302 486 4320
rect 468 4320 486 4338
rect 468 4338 486 4356
rect 468 4356 486 4374
rect 468 4374 486 4392
rect 468 4392 486 4410
rect 468 4410 486 4428
rect 468 4428 486 4446
rect 468 4446 486 4464
rect 468 4464 486 4482
rect 468 4482 486 4500
rect 468 4500 486 4518
rect 468 4518 486 4536
rect 468 4536 486 4554
rect 468 4554 486 4572
rect 468 4572 486 4590
rect 468 4590 486 4608
rect 468 4608 486 4626
rect 468 4626 486 4644
rect 468 4644 486 4662
rect 468 4662 486 4680
rect 468 4680 486 4698
rect 468 4698 486 4716
rect 468 4716 486 4734
rect 468 4734 486 4752
rect 468 4752 486 4770
rect 468 4770 486 4788
rect 468 4788 486 4806
rect 468 4806 486 4824
rect 468 4824 486 4842
rect 468 4842 486 4860
rect 468 4860 486 4878
rect 468 4878 486 4896
rect 468 4896 486 4914
rect 468 4914 486 4932
rect 468 4932 486 4950
rect 468 4950 486 4968
rect 468 4968 486 4986
rect 468 4986 486 5004
rect 468 5004 486 5022
rect 468 5022 486 5040
rect 468 5040 486 5058
rect 468 5058 486 5076
rect 468 5076 486 5094
rect 468 5094 486 5112
rect 468 5112 486 5130
rect 468 5130 486 5148
rect 468 5148 486 5166
rect 468 5166 486 5184
rect 468 5184 486 5202
rect 468 5202 486 5220
rect 468 5220 486 5238
rect 468 5238 486 5256
rect 468 5256 486 5274
rect 468 5274 486 5292
rect 468 5292 486 5310
rect 468 5310 486 5328
rect 468 5328 486 5346
rect 468 5346 486 5364
rect 468 5364 486 5382
rect 468 5382 486 5400
rect 468 5400 486 5418
rect 468 5418 486 5436
rect 486 1818 504 1836
rect 486 1836 504 1854
rect 486 1854 504 1872
rect 486 1872 504 1890
rect 486 1890 504 1908
rect 486 1908 504 1926
rect 486 1926 504 1944
rect 486 1944 504 1962
rect 486 1962 504 1980
rect 486 1980 504 1998
rect 486 1998 504 2016
rect 486 2016 504 2034
rect 486 2034 504 2052
rect 486 2052 504 2070
rect 486 2070 504 2088
rect 486 2088 504 2106
rect 486 2106 504 2124
rect 486 2124 504 2142
rect 486 2142 504 2160
rect 486 2160 504 2178
rect 486 2178 504 2196
rect 486 2196 504 2214
rect 486 2214 504 2232
rect 486 2232 504 2250
rect 486 2250 504 2268
rect 486 2268 504 2286
rect 486 2286 504 2304
rect 486 2304 504 2322
rect 486 2322 504 2340
rect 486 2340 504 2358
rect 486 2358 504 2376
rect 486 2376 504 2394
rect 486 2394 504 2412
rect 486 2412 504 2430
rect 486 2430 504 2448
rect 486 2448 504 2466
rect 486 2466 504 2484
rect 486 2484 504 2502
rect 486 2502 504 2520
rect 486 2520 504 2538
rect 486 2538 504 2556
rect 486 2556 504 2574
rect 486 2574 504 2592
rect 486 2592 504 2610
rect 486 2610 504 2628
rect 486 2628 504 2646
rect 486 2646 504 2664
rect 486 2664 504 2682
rect 486 2682 504 2700
rect 486 2700 504 2718
rect 486 2718 504 2736
rect 486 2736 504 2754
rect 486 2754 504 2772
rect 486 2772 504 2790
rect 486 2790 504 2808
rect 486 2808 504 2826
rect 486 2826 504 2844
rect 486 2844 504 2862
rect 486 2862 504 2880
rect 486 2880 504 2898
rect 486 2898 504 2916
rect 486 2916 504 2934
rect 486 2934 504 2952
rect 486 2952 504 2970
rect 486 2970 504 2988
rect 486 2988 504 3006
rect 486 3006 504 3024
rect 486 3024 504 3042
rect 486 3042 504 3060
rect 486 3060 504 3078
rect 486 3078 504 3096
rect 486 3096 504 3114
rect 486 3114 504 3132
rect 486 3132 504 3150
rect 486 3150 504 3168
rect 486 3168 504 3186
rect 486 3186 504 3204
rect 486 3204 504 3222
rect 486 3222 504 3240
rect 486 3240 504 3258
rect 486 3258 504 3276
rect 486 3276 504 3294
rect 486 3294 504 3312
rect 486 3312 504 3330
rect 486 3330 504 3348
rect 486 3348 504 3366
rect 486 3366 504 3384
rect 486 3384 504 3402
rect 486 3402 504 3420
rect 486 3420 504 3438
rect 486 3438 504 3456
rect 486 3456 504 3474
rect 486 3474 504 3492
rect 486 3492 504 3510
rect 486 3510 504 3528
rect 486 3528 504 3546
rect 486 3546 504 3564
rect 486 3564 504 3582
rect 486 3582 504 3600
rect 486 3600 504 3618
rect 486 3618 504 3636
rect 486 3636 504 3654
rect 486 3654 504 3672
rect 486 3672 504 3690
rect 486 3690 504 3708
rect 486 3708 504 3726
rect 486 3726 504 3744
rect 486 3744 504 3762
rect 486 3762 504 3780
rect 486 3780 504 3798
rect 486 3798 504 3816
rect 486 3816 504 3834
rect 486 3834 504 3852
rect 486 3852 504 3870
rect 486 3870 504 3888
rect 486 3888 504 3906
rect 486 3906 504 3924
rect 486 3924 504 3942
rect 486 3942 504 3960
rect 486 3960 504 3978
rect 486 3978 504 3996
rect 486 3996 504 4014
rect 486 4014 504 4032
rect 486 4032 504 4050
rect 486 4050 504 4068
rect 486 4068 504 4086
rect 486 4086 504 4104
rect 486 4104 504 4122
rect 486 4122 504 4140
rect 486 4140 504 4158
rect 486 4158 504 4176
rect 486 4176 504 4194
rect 486 4194 504 4212
rect 486 4212 504 4230
rect 486 4230 504 4248
rect 486 4248 504 4266
rect 486 4266 504 4284
rect 486 4284 504 4302
rect 486 4302 504 4320
rect 486 4320 504 4338
rect 486 4338 504 4356
rect 486 4356 504 4374
rect 486 4374 504 4392
rect 486 4392 504 4410
rect 486 4410 504 4428
rect 486 4428 504 4446
rect 486 4446 504 4464
rect 486 4464 504 4482
rect 486 4482 504 4500
rect 486 4500 504 4518
rect 486 4518 504 4536
rect 486 4536 504 4554
rect 486 4554 504 4572
rect 486 4572 504 4590
rect 486 4590 504 4608
rect 486 4608 504 4626
rect 486 4626 504 4644
rect 486 4644 504 4662
rect 486 4662 504 4680
rect 486 4680 504 4698
rect 486 4698 504 4716
rect 486 4716 504 4734
rect 486 4734 504 4752
rect 486 4752 504 4770
rect 486 4770 504 4788
rect 486 4788 504 4806
rect 486 4806 504 4824
rect 486 4824 504 4842
rect 486 4842 504 4860
rect 486 4860 504 4878
rect 486 4878 504 4896
rect 486 4896 504 4914
rect 486 4914 504 4932
rect 486 4932 504 4950
rect 486 4950 504 4968
rect 486 4968 504 4986
rect 486 4986 504 5004
rect 486 5004 504 5022
rect 486 5022 504 5040
rect 486 5040 504 5058
rect 486 5058 504 5076
rect 486 5076 504 5094
rect 486 5094 504 5112
rect 486 5112 504 5130
rect 486 5130 504 5148
rect 486 5148 504 5166
rect 486 5166 504 5184
rect 486 5184 504 5202
rect 486 5202 504 5220
rect 486 5220 504 5238
rect 486 5238 504 5256
rect 486 5256 504 5274
rect 486 5274 504 5292
rect 486 5292 504 5310
rect 486 5310 504 5328
rect 486 5328 504 5346
rect 486 5346 504 5364
rect 486 5364 504 5382
rect 486 5382 504 5400
rect 486 5400 504 5418
rect 486 5418 504 5436
rect 486 5436 504 5454
rect 504 1782 522 1800
rect 504 1800 522 1818
rect 504 1818 522 1836
rect 504 1836 522 1854
rect 504 1854 522 1872
rect 504 1872 522 1890
rect 504 1890 522 1908
rect 504 1908 522 1926
rect 504 1926 522 1944
rect 504 1944 522 1962
rect 504 1962 522 1980
rect 504 1980 522 1998
rect 504 1998 522 2016
rect 504 2016 522 2034
rect 504 2034 522 2052
rect 504 2052 522 2070
rect 504 2070 522 2088
rect 504 2088 522 2106
rect 504 2106 522 2124
rect 504 2124 522 2142
rect 504 2142 522 2160
rect 504 2160 522 2178
rect 504 2178 522 2196
rect 504 2196 522 2214
rect 504 2214 522 2232
rect 504 2232 522 2250
rect 504 2250 522 2268
rect 504 2268 522 2286
rect 504 2286 522 2304
rect 504 2304 522 2322
rect 504 2322 522 2340
rect 504 2340 522 2358
rect 504 2358 522 2376
rect 504 2376 522 2394
rect 504 2394 522 2412
rect 504 2412 522 2430
rect 504 2430 522 2448
rect 504 2448 522 2466
rect 504 2466 522 2484
rect 504 2484 522 2502
rect 504 2502 522 2520
rect 504 2520 522 2538
rect 504 2538 522 2556
rect 504 2556 522 2574
rect 504 2574 522 2592
rect 504 2592 522 2610
rect 504 2610 522 2628
rect 504 2628 522 2646
rect 504 2646 522 2664
rect 504 2664 522 2682
rect 504 2682 522 2700
rect 504 2700 522 2718
rect 504 2718 522 2736
rect 504 2736 522 2754
rect 504 2754 522 2772
rect 504 2772 522 2790
rect 504 2790 522 2808
rect 504 2808 522 2826
rect 504 2826 522 2844
rect 504 2844 522 2862
rect 504 2862 522 2880
rect 504 2880 522 2898
rect 504 2898 522 2916
rect 504 2916 522 2934
rect 504 2934 522 2952
rect 504 2952 522 2970
rect 504 2970 522 2988
rect 504 2988 522 3006
rect 504 3006 522 3024
rect 504 3024 522 3042
rect 504 3042 522 3060
rect 504 3060 522 3078
rect 504 3078 522 3096
rect 504 3096 522 3114
rect 504 3114 522 3132
rect 504 3132 522 3150
rect 504 3150 522 3168
rect 504 3168 522 3186
rect 504 3186 522 3204
rect 504 3204 522 3222
rect 504 3222 522 3240
rect 504 3240 522 3258
rect 504 3258 522 3276
rect 504 3276 522 3294
rect 504 3294 522 3312
rect 504 3312 522 3330
rect 504 3330 522 3348
rect 504 3348 522 3366
rect 504 3366 522 3384
rect 504 3384 522 3402
rect 504 3402 522 3420
rect 504 3420 522 3438
rect 504 3438 522 3456
rect 504 3456 522 3474
rect 504 3474 522 3492
rect 504 3492 522 3510
rect 504 3510 522 3528
rect 504 3528 522 3546
rect 504 3546 522 3564
rect 504 3564 522 3582
rect 504 3582 522 3600
rect 504 3600 522 3618
rect 504 3618 522 3636
rect 504 3636 522 3654
rect 504 3654 522 3672
rect 504 3672 522 3690
rect 504 3690 522 3708
rect 504 3708 522 3726
rect 504 3726 522 3744
rect 504 3744 522 3762
rect 504 3762 522 3780
rect 504 3780 522 3798
rect 504 3798 522 3816
rect 504 3816 522 3834
rect 504 3834 522 3852
rect 504 3852 522 3870
rect 504 3870 522 3888
rect 504 3888 522 3906
rect 504 3906 522 3924
rect 504 3924 522 3942
rect 504 3942 522 3960
rect 504 3960 522 3978
rect 504 3978 522 3996
rect 504 3996 522 4014
rect 504 4014 522 4032
rect 504 4032 522 4050
rect 504 4050 522 4068
rect 504 4068 522 4086
rect 504 4086 522 4104
rect 504 4104 522 4122
rect 504 4122 522 4140
rect 504 4140 522 4158
rect 504 4158 522 4176
rect 504 4176 522 4194
rect 504 4194 522 4212
rect 504 4212 522 4230
rect 504 4230 522 4248
rect 504 4248 522 4266
rect 504 4266 522 4284
rect 504 4284 522 4302
rect 504 4302 522 4320
rect 504 4320 522 4338
rect 504 4338 522 4356
rect 504 4356 522 4374
rect 504 4374 522 4392
rect 504 4392 522 4410
rect 504 4410 522 4428
rect 504 4428 522 4446
rect 504 4446 522 4464
rect 504 4464 522 4482
rect 504 4482 522 4500
rect 504 4500 522 4518
rect 504 4518 522 4536
rect 504 4536 522 4554
rect 504 4554 522 4572
rect 504 4572 522 4590
rect 504 4590 522 4608
rect 504 4608 522 4626
rect 504 4626 522 4644
rect 504 4644 522 4662
rect 504 4662 522 4680
rect 504 4680 522 4698
rect 504 4698 522 4716
rect 504 4716 522 4734
rect 504 4734 522 4752
rect 504 4752 522 4770
rect 504 4770 522 4788
rect 504 4788 522 4806
rect 504 4806 522 4824
rect 504 4824 522 4842
rect 504 4842 522 4860
rect 504 4860 522 4878
rect 504 4878 522 4896
rect 504 4896 522 4914
rect 504 4914 522 4932
rect 504 4932 522 4950
rect 504 4950 522 4968
rect 504 4968 522 4986
rect 504 4986 522 5004
rect 504 5004 522 5022
rect 504 5022 522 5040
rect 504 5040 522 5058
rect 504 5058 522 5076
rect 504 5076 522 5094
rect 504 5094 522 5112
rect 504 5112 522 5130
rect 504 5130 522 5148
rect 504 5148 522 5166
rect 504 5166 522 5184
rect 504 5184 522 5202
rect 504 5202 522 5220
rect 504 5220 522 5238
rect 504 5238 522 5256
rect 504 5256 522 5274
rect 504 5274 522 5292
rect 504 5292 522 5310
rect 504 5310 522 5328
rect 504 5328 522 5346
rect 504 5346 522 5364
rect 504 5364 522 5382
rect 504 5382 522 5400
rect 504 5400 522 5418
rect 504 5418 522 5436
rect 504 5436 522 5454
rect 504 5454 522 5472
rect 504 5472 522 5490
rect 522 1746 540 1764
rect 522 1764 540 1782
rect 522 1782 540 1800
rect 522 1800 540 1818
rect 522 1818 540 1836
rect 522 1836 540 1854
rect 522 1854 540 1872
rect 522 1872 540 1890
rect 522 1890 540 1908
rect 522 1908 540 1926
rect 522 1926 540 1944
rect 522 1944 540 1962
rect 522 1962 540 1980
rect 522 1980 540 1998
rect 522 1998 540 2016
rect 522 2016 540 2034
rect 522 2034 540 2052
rect 522 2052 540 2070
rect 522 2070 540 2088
rect 522 2088 540 2106
rect 522 2106 540 2124
rect 522 2124 540 2142
rect 522 2142 540 2160
rect 522 2160 540 2178
rect 522 2178 540 2196
rect 522 2196 540 2214
rect 522 2214 540 2232
rect 522 2232 540 2250
rect 522 2250 540 2268
rect 522 2268 540 2286
rect 522 2286 540 2304
rect 522 2304 540 2322
rect 522 2322 540 2340
rect 522 2340 540 2358
rect 522 2358 540 2376
rect 522 2376 540 2394
rect 522 2394 540 2412
rect 522 2412 540 2430
rect 522 2430 540 2448
rect 522 2448 540 2466
rect 522 2466 540 2484
rect 522 2484 540 2502
rect 522 2502 540 2520
rect 522 2520 540 2538
rect 522 2538 540 2556
rect 522 2556 540 2574
rect 522 2574 540 2592
rect 522 2592 540 2610
rect 522 2610 540 2628
rect 522 2628 540 2646
rect 522 2646 540 2664
rect 522 2664 540 2682
rect 522 2682 540 2700
rect 522 2700 540 2718
rect 522 2718 540 2736
rect 522 2736 540 2754
rect 522 2754 540 2772
rect 522 2772 540 2790
rect 522 2790 540 2808
rect 522 2808 540 2826
rect 522 2826 540 2844
rect 522 2844 540 2862
rect 522 2862 540 2880
rect 522 2880 540 2898
rect 522 2898 540 2916
rect 522 2916 540 2934
rect 522 2934 540 2952
rect 522 2952 540 2970
rect 522 2970 540 2988
rect 522 2988 540 3006
rect 522 3006 540 3024
rect 522 3024 540 3042
rect 522 3042 540 3060
rect 522 3060 540 3078
rect 522 3078 540 3096
rect 522 3096 540 3114
rect 522 3114 540 3132
rect 522 3132 540 3150
rect 522 3150 540 3168
rect 522 3168 540 3186
rect 522 3186 540 3204
rect 522 3204 540 3222
rect 522 3222 540 3240
rect 522 3240 540 3258
rect 522 3258 540 3276
rect 522 3276 540 3294
rect 522 3294 540 3312
rect 522 3312 540 3330
rect 522 3330 540 3348
rect 522 3348 540 3366
rect 522 3366 540 3384
rect 522 3384 540 3402
rect 522 3402 540 3420
rect 522 3420 540 3438
rect 522 3438 540 3456
rect 522 3456 540 3474
rect 522 3474 540 3492
rect 522 3492 540 3510
rect 522 3510 540 3528
rect 522 3528 540 3546
rect 522 3546 540 3564
rect 522 3564 540 3582
rect 522 3582 540 3600
rect 522 3600 540 3618
rect 522 3618 540 3636
rect 522 3636 540 3654
rect 522 3654 540 3672
rect 522 3672 540 3690
rect 522 3690 540 3708
rect 522 3708 540 3726
rect 522 3726 540 3744
rect 522 3744 540 3762
rect 522 3762 540 3780
rect 522 3780 540 3798
rect 522 3798 540 3816
rect 522 3816 540 3834
rect 522 3834 540 3852
rect 522 3852 540 3870
rect 522 3870 540 3888
rect 522 3888 540 3906
rect 522 3906 540 3924
rect 522 3924 540 3942
rect 522 3942 540 3960
rect 522 3960 540 3978
rect 522 3978 540 3996
rect 522 3996 540 4014
rect 522 4014 540 4032
rect 522 4032 540 4050
rect 522 4050 540 4068
rect 522 4068 540 4086
rect 522 4086 540 4104
rect 522 4104 540 4122
rect 522 4122 540 4140
rect 522 4140 540 4158
rect 522 4158 540 4176
rect 522 4176 540 4194
rect 522 4194 540 4212
rect 522 4212 540 4230
rect 522 4230 540 4248
rect 522 4248 540 4266
rect 522 4266 540 4284
rect 522 4284 540 4302
rect 522 4302 540 4320
rect 522 4320 540 4338
rect 522 4338 540 4356
rect 522 4356 540 4374
rect 522 4374 540 4392
rect 522 4392 540 4410
rect 522 4410 540 4428
rect 522 4428 540 4446
rect 522 4446 540 4464
rect 522 4464 540 4482
rect 522 4482 540 4500
rect 522 4500 540 4518
rect 522 4518 540 4536
rect 522 4536 540 4554
rect 522 4554 540 4572
rect 522 4572 540 4590
rect 522 4590 540 4608
rect 522 4608 540 4626
rect 522 4626 540 4644
rect 522 4644 540 4662
rect 522 4662 540 4680
rect 522 4680 540 4698
rect 522 4698 540 4716
rect 522 4716 540 4734
rect 522 4734 540 4752
rect 522 4752 540 4770
rect 522 4770 540 4788
rect 522 4788 540 4806
rect 522 4806 540 4824
rect 522 4824 540 4842
rect 522 4842 540 4860
rect 522 4860 540 4878
rect 522 4878 540 4896
rect 522 4896 540 4914
rect 522 4914 540 4932
rect 522 4932 540 4950
rect 522 4950 540 4968
rect 522 4968 540 4986
rect 522 4986 540 5004
rect 522 5004 540 5022
rect 522 5022 540 5040
rect 522 5040 540 5058
rect 522 5058 540 5076
rect 522 5076 540 5094
rect 522 5094 540 5112
rect 522 5112 540 5130
rect 522 5130 540 5148
rect 522 5148 540 5166
rect 522 5166 540 5184
rect 522 5184 540 5202
rect 522 5202 540 5220
rect 522 5220 540 5238
rect 522 5238 540 5256
rect 522 5256 540 5274
rect 522 5274 540 5292
rect 522 5292 540 5310
rect 522 5310 540 5328
rect 522 5328 540 5346
rect 522 5346 540 5364
rect 522 5364 540 5382
rect 522 5382 540 5400
rect 522 5400 540 5418
rect 522 5418 540 5436
rect 522 5436 540 5454
rect 522 5454 540 5472
rect 522 5472 540 5490
rect 522 5490 540 5508
rect 522 5508 540 5526
rect 540 1728 558 1746
rect 540 1746 558 1764
rect 540 1764 558 1782
rect 540 1782 558 1800
rect 540 1800 558 1818
rect 540 1818 558 1836
rect 540 1836 558 1854
rect 540 1854 558 1872
rect 540 1872 558 1890
rect 540 1890 558 1908
rect 540 1908 558 1926
rect 540 1926 558 1944
rect 540 1944 558 1962
rect 540 1962 558 1980
rect 540 1980 558 1998
rect 540 1998 558 2016
rect 540 2016 558 2034
rect 540 2034 558 2052
rect 540 2052 558 2070
rect 540 2070 558 2088
rect 540 2088 558 2106
rect 540 2106 558 2124
rect 540 2124 558 2142
rect 540 2142 558 2160
rect 540 2160 558 2178
rect 540 2178 558 2196
rect 540 2196 558 2214
rect 540 2214 558 2232
rect 540 2232 558 2250
rect 540 2250 558 2268
rect 540 2268 558 2286
rect 540 2286 558 2304
rect 540 2304 558 2322
rect 540 2322 558 2340
rect 540 2340 558 2358
rect 540 2358 558 2376
rect 540 2376 558 2394
rect 540 2394 558 2412
rect 540 2412 558 2430
rect 540 2430 558 2448
rect 540 2448 558 2466
rect 540 2466 558 2484
rect 540 2484 558 2502
rect 540 2502 558 2520
rect 540 2520 558 2538
rect 540 2538 558 2556
rect 540 2556 558 2574
rect 540 2574 558 2592
rect 540 2592 558 2610
rect 540 2610 558 2628
rect 540 2628 558 2646
rect 540 2646 558 2664
rect 540 2664 558 2682
rect 540 2682 558 2700
rect 540 2700 558 2718
rect 540 2718 558 2736
rect 540 2736 558 2754
rect 540 2754 558 2772
rect 540 2772 558 2790
rect 540 2790 558 2808
rect 540 2808 558 2826
rect 540 2826 558 2844
rect 540 2844 558 2862
rect 540 2862 558 2880
rect 540 2880 558 2898
rect 540 2898 558 2916
rect 540 2916 558 2934
rect 540 2934 558 2952
rect 540 2952 558 2970
rect 540 2970 558 2988
rect 540 2988 558 3006
rect 540 3006 558 3024
rect 540 3024 558 3042
rect 540 3042 558 3060
rect 540 3060 558 3078
rect 540 3078 558 3096
rect 540 3096 558 3114
rect 540 3114 558 3132
rect 540 3132 558 3150
rect 540 3150 558 3168
rect 540 3168 558 3186
rect 540 3186 558 3204
rect 540 3204 558 3222
rect 540 3222 558 3240
rect 540 3240 558 3258
rect 540 3258 558 3276
rect 540 3276 558 3294
rect 540 3294 558 3312
rect 540 3312 558 3330
rect 540 3330 558 3348
rect 540 3348 558 3366
rect 540 3366 558 3384
rect 540 3384 558 3402
rect 540 3402 558 3420
rect 540 3420 558 3438
rect 540 3438 558 3456
rect 540 3456 558 3474
rect 540 3474 558 3492
rect 540 3492 558 3510
rect 540 3510 558 3528
rect 540 3528 558 3546
rect 540 3546 558 3564
rect 540 3564 558 3582
rect 540 3582 558 3600
rect 540 3600 558 3618
rect 540 3618 558 3636
rect 540 3636 558 3654
rect 540 3654 558 3672
rect 540 3672 558 3690
rect 540 3690 558 3708
rect 540 3708 558 3726
rect 540 3726 558 3744
rect 540 3744 558 3762
rect 540 3762 558 3780
rect 540 3780 558 3798
rect 540 3798 558 3816
rect 540 3816 558 3834
rect 540 3834 558 3852
rect 540 3852 558 3870
rect 540 3870 558 3888
rect 540 3888 558 3906
rect 540 3906 558 3924
rect 540 3924 558 3942
rect 540 3942 558 3960
rect 540 3960 558 3978
rect 540 3978 558 3996
rect 540 3996 558 4014
rect 540 4014 558 4032
rect 540 4032 558 4050
rect 540 4050 558 4068
rect 540 4068 558 4086
rect 540 4086 558 4104
rect 540 4104 558 4122
rect 540 4122 558 4140
rect 540 4140 558 4158
rect 540 4158 558 4176
rect 540 4176 558 4194
rect 540 4194 558 4212
rect 540 4212 558 4230
rect 540 4230 558 4248
rect 540 4248 558 4266
rect 540 4266 558 4284
rect 540 4284 558 4302
rect 540 4302 558 4320
rect 540 4320 558 4338
rect 540 4338 558 4356
rect 540 4356 558 4374
rect 540 4374 558 4392
rect 540 4392 558 4410
rect 540 4410 558 4428
rect 540 4428 558 4446
rect 540 4446 558 4464
rect 540 4464 558 4482
rect 540 4482 558 4500
rect 540 4500 558 4518
rect 540 4518 558 4536
rect 540 4536 558 4554
rect 540 4554 558 4572
rect 540 4572 558 4590
rect 540 4590 558 4608
rect 540 4608 558 4626
rect 540 4626 558 4644
rect 540 4644 558 4662
rect 540 4662 558 4680
rect 540 4680 558 4698
rect 540 4698 558 4716
rect 540 4716 558 4734
rect 540 4734 558 4752
rect 540 4752 558 4770
rect 540 4770 558 4788
rect 540 4788 558 4806
rect 540 4806 558 4824
rect 540 4824 558 4842
rect 540 4842 558 4860
rect 540 4860 558 4878
rect 540 4878 558 4896
rect 540 4896 558 4914
rect 540 4914 558 4932
rect 540 4932 558 4950
rect 540 4950 558 4968
rect 540 4968 558 4986
rect 540 4986 558 5004
rect 540 5004 558 5022
rect 540 5022 558 5040
rect 540 5040 558 5058
rect 540 5058 558 5076
rect 540 5076 558 5094
rect 540 5094 558 5112
rect 540 5112 558 5130
rect 540 5130 558 5148
rect 540 5148 558 5166
rect 540 5166 558 5184
rect 540 5184 558 5202
rect 540 5202 558 5220
rect 540 5220 558 5238
rect 540 5238 558 5256
rect 540 5256 558 5274
rect 540 5274 558 5292
rect 540 5292 558 5310
rect 540 5310 558 5328
rect 540 5328 558 5346
rect 540 5346 558 5364
rect 540 5364 558 5382
rect 540 5382 558 5400
rect 540 5400 558 5418
rect 540 5418 558 5436
rect 540 5436 558 5454
rect 540 5454 558 5472
rect 540 5472 558 5490
rect 540 5490 558 5508
rect 540 5508 558 5526
rect 540 5526 558 5544
rect 558 1692 576 1710
rect 558 1710 576 1728
rect 558 1728 576 1746
rect 558 1746 576 1764
rect 558 1764 576 1782
rect 558 1782 576 1800
rect 558 1800 576 1818
rect 558 1818 576 1836
rect 558 1836 576 1854
rect 558 1854 576 1872
rect 558 1872 576 1890
rect 558 1890 576 1908
rect 558 1908 576 1926
rect 558 1926 576 1944
rect 558 1944 576 1962
rect 558 1962 576 1980
rect 558 1980 576 1998
rect 558 1998 576 2016
rect 558 2016 576 2034
rect 558 2034 576 2052
rect 558 2052 576 2070
rect 558 2070 576 2088
rect 558 2088 576 2106
rect 558 2106 576 2124
rect 558 2124 576 2142
rect 558 2142 576 2160
rect 558 2160 576 2178
rect 558 2178 576 2196
rect 558 2196 576 2214
rect 558 2214 576 2232
rect 558 2232 576 2250
rect 558 2250 576 2268
rect 558 2268 576 2286
rect 558 2286 576 2304
rect 558 2304 576 2322
rect 558 2322 576 2340
rect 558 2340 576 2358
rect 558 2358 576 2376
rect 558 2376 576 2394
rect 558 2394 576 2412
rect 558 2412 576 2430
rect 558 2430 576 2448
rect 558 2448 576 2466
rect 558 2466 576 2484
rect 558 2484 576 2502
rect 558 2502 576 2520
rect 558 2520 576 2538
rect 558 2538 576 2556
rect 558 2556 576 2574
rect 558 2574 576 2592
rect 558 2592 576 2610
rect 558 2610 576 2628
rect 558 2628 576 2646
rect 558 2646 576 2664
rect 558 2664 576 2682
rect 558 2682 576 2700
rect 558 2700 576 2718
rect 558 2718 576 2736
rect 558 2736 576 2754
rect 558 2754 576 2772
rect 558 2772 576 2790
rect 558 2790 576 2808
rect 558 2808 576 2826
rect 558 2826 576 2844
rect 558 2844 576 2862
rect 558 2862 576 2880
rect 558 2880 576 2898
rect 558 2898 576 2916
rect 558 2916 576 2934
rect 558 2934 576 2952
rect 558 2952 576 2970
rect 558 2970 576 2988
rect 558 2988 576 3006
rect 558 3006 576 3024
rect 558 3024 576 3042
rect 558 3042 576 3060
rect 558 3060 576 3078
rect 558 3078 576 3096
rect 558 3096 576 3114
rect 558 3114 576 3132
rect 558 3132 576 3150
rect 558 3150 576 3168
rect 558 3168 576 3186
rect 558 3186 576 3204
rect 558 3204 576 3222
rect 558 3222 576 3240
rect 558 3240 576 3258
rect 558 3258 576 3276
rect 558 3276 576 3294
rect 558 3294 576 3312
rect 558 3312 576 3330
rect 558 3330 576 3348
rect 558 3348 576 3366
rect 558 3366 576 3384
rect 558 3384 576 3402
rect 558 3402 576 3420
rect 558 3420 576 3438
rect 558 3438 576 3456
rect 558 3456 576 3474
rect 558 3474 576 3492
rect 558 3492 576 3510
rect 558 3510 576 3528
rect 558 3528 576 3546
rect 558 3546 576 3564
rect 558 3564 576 3582
rect 558 3582 576 3600
rect 558 3600 576 3618
rect 558 3618 576 3636
rect 558 3636 576 3654
rect 558 3654 576 3672
rect 558 3672 576 3690
rect 558 3690 576 3708
rect 558 3708 576 3726
rect 558 3726 576 3744
rect 558 3744 576 3762
rect 558 3762 576 3780
rect 558 3780 576 3798
rect 558 3798 576 3816
rect 558 3816 576 3834
rect 558 3834 576 3852
rect 558 3852 576 3870
rect 558 3870 576 3888
rect 558 3888 576 3906
rect 558 3906 576 3924
rect 558 3924 576 3942
rect 558 3942 576 3960
rect 558 3960 576 3978
rect 558 3978 576 3996
rect 558 3996 576 4014
rect 558 4014 576 4032
rect 558 4032 576 4050
rect 558 4050 576 4068
rect 558 4068 576 4086
rect 558 4086 576 4104
rect 558 4104 576 4122
rect 558 4122 576 4140
rect 558 4140 576 4158
rect 558 4158 576 4176
rect 558 4176 576 4194
rect 558 4194 576 4212
rect 558 4212 576 4230
rect 558 4230 576 4248
rect 558 4248 576 4266
rect 558 4266 576 4284
rect 558 4284 576 4302
rect 558 4302 576 4320
rect 558 4320 576 4338
rect 558 4338 576 4356
rect 558 4356 576 4374
rect 558 4374 576 4392
rect 558 4392 576 4410
rect 558 4410 576 4428
rect 558 4428 576 4446
rect 558 4446 576 4464
rect 558 4464 576 4482
rect 558 4482 576 4500
rect 558 4500 576 4518
rect 558 4518 576 4536
rect 558 4536 576 4554
rect 558 4554 576 4572
rect 558 4572 576 4590
rect 558 4590 576 4608
rect 558 4608 576 4626
rect 558 4626 576 4644
rect 558 4644 576 4662
rect 558 4662 576 4680
rect 558 4680 576 4698
rect 558 4698 576 4716
rect 558 4716 576 4734
rect 558 4734 576 4752
rect 558 4752 576 4770
rect 558 4770 576 4788
rect 558 4788 576 4806
rect 558 4806 576 4824
rect 558 4824 576 4842
rect 558 4842 576 4860
rect 558 4860 576 4878
rect 558 4878 576 4896
rect 558 4896 576 4914
rect 558 4914 576 4932
rect 558 4932 576 4950
rect 558 4950 576 4968
rect 558 4968 576 4986
rect 558 4986 576 5004
rect 558 5004 576 5022
rect 558 5022 576 5040
rect 558 5040 576 5058
rect 558 5058 576 5076
rect 558 5076 576 5094
rect 558 5094 576 5112
rect 558 5112 576 5130
rect 558 5130 576 5148
rect 558 5148 576 5166
rect 558 5166 576 5184
rect 558 5184 576 5202
rect 558 5202 576 5220
rect 558 5220 576 5238
rect 558 5238 576 5256
rect 558 5256 576 5274
rect 558 5274 576 5292
rect 558 5292 576 5310
rect 558 5310 576 5328
rect 558 5328 576 5346
rect 558 5346 576 5364
rect 558 5364 576 5382
rect 558 5382 576 5400
rect 558 5400 576 5418
rect 558 5418 576 5436
rect 558 5436 576 5454
rect 558 5454 576 5472
rect 558 5472 576 5490
rect 558 5490 576 5508
rect 558 5508 576 5526
rect 558 5526 576 5544
rect 558 5544 576 5562
rect 558 5562 576 5580
rect 576 1656 594 1674
rect 576 1674 594 1692
rect 576 1692 594 1710
rect 576 1710 594 1728
rect 576 1728 594 1746
rect 576 1746 594 1764
rect 576 1764 594 1782
rect 576 1782 594 1800
rect 576 1800 594 1818
rect 576 1818 594 1836
rect 576 1836 594 1854
rect 576 1854 594 1872
rect 576 1872 594 1890
rect 576 1890 594 1908
rect 576 1908 594 1926
rect 576 1926 594 1944
rect 576 1944 594 1962
rect 576 1962 594 1980
rect 576 1980 594 1998
rect 576 1998 594 2016
rect 576 2016 594 2034
rect 576 2034 594 2052
rect 576 2052 594 2070
rect 576 2070 594 2088
rect 576 2088 594 2106
rect 576 2106 594 2124
rect 576 2124 594 2142
rect 576 2142 594 2160
rect 576 2160 594 2178
rect 576 2178 594 2196
rect 576 2196 594 2214
rect 576 2214 594 2232
rect 576 2232 594 2250
rect 576 2250 594 2268
rect 576 2268 594 2286
rect 576 2286 594 2304
rect 576 2304 594 2322
rect 576 2322 594 2340
rect 576 2340 594 2358
rect 576 2358 594 2376
rect 576 2376 594 2394
rect 576 2394 594 2412
rect 576 2412 594 2430
rect 576 2430 594 2448
rect 576 2448 594 2466
rect 576 2466 594 2484
rect 576 2484 594 2502
rect 576 2502 594 2520
rect 576 2520 594 2538
rect 576 2538 594 2556
rect 576 2556 594 2574
rect 576 2574 594 2592
rect 576 2592 594 2610
rect 576 2610 594 2628
rect 576 2628 594 2646
rect 576 2646 594 2664
rect 576 2664 594 2682
rect 576 2682 594 2700
rect 576 2700 594 2718
rect 576 2718 594 2736
rect 576 2736 594 2754
rect 576 2754 594 2772
rect 576 2772 594 2790
rect 576 2790 594 2808
rect 576 2808 594 2826
rect 576 2826 594 2844
rect 576 2844 594 2862
rect 576 2862 594 2880
rect 576 2880 594 2898
rect 576 2898 594 2916
rect 576 2916 594 2934
rect 576 2934 594 2952
rect 576 2952 594 2970
rect 576 2970 594 2988
rect 576 2988 594 3006
rect 576 3006 594 3024
rect 576 3024 594 3042
rect 576 3042 594 3060
rect 576 3060 594 3078
rect 576 3078 594 3096
rect 576 3096 594 3114
rect 576 3114 594 3132
rect 576 3132 594 3150
rect 576 3150 594 3168
rect 576 3168 594 3186
rect 576 3186 594 3204
rect 576 3204 594 3222
rect 576 3222 594 3240
rect 576 3240 594 3258
rect 576 3258 594 3276
rect 576 3276 594 3294
rect 576 3294 594 3312
rect 576 3312 594 3330
rect 576 3330 594 3348
rect 576 3348 594 3366
rect 576 3366 594 3384
rect 576 3384 594 3402
rect 576 3402 594 3420
rect 576 3420 594 3438
rect 576 3438 594 3456
rect 576 3456 594 3474
rect 576 3474 594 3492
rect 576 3492 594 3510
rect 576 3510 594 3528
rect 576 3528 594 3546
rect 576 3546 594 3564
rect 576 3564 594 3582
rect 576 3582 594 3600
rect 576 3600 594 3618
rect 576 3618 594 3636
rect 576 3636 594 3654
rect 576 3654 594 3672
rect 576 3672 594 3690
rect 576 3690 594 3708
rect 576 3708 594 3726
rect 576 3726 594 3744
rect 576 3744 594 3762
rect 576 3762 594 3780
rect 576 3780 594 3798
rect 576 3798 594 3816
rect 576 3816 594 3834
rect 576 3834 594 3852
rect 576 3852 594 3870
rect 576 3870 594 3888
rect 576 3888 594 3906
rect 576 3906 594 3924
rect 576 3924 594 3942
rect 576 3942 594 3960
rect 576 3960 594 3978
rect 576 3978 594 3996
rect 576 3996 594 4014
rect 576 4014 594 4032
rect 576 4032 594 4050
rect 576 4050 594 4068
rect 576 4068 594 4086
rect 576 4086 594 4104
rect 576 4104 594 4122
rect 576 4122 594 4140
rect 576 4140 594 4158
rect 576 4158 594 4176
rect 576 4176 594 4194
rect 576 4194 594 4212
rect 576 4212 594 4230
rect 576 4230 594 4248
rect 576 4248 594 4266
rect 576 4266 594 4284
rect 576 4284 594 4302
rect 576 4302 594 4320
rect 576 4320 594 4338
rect 576 4338 594 4356
rect 576 4356 594 4374
rect 576 4374 594 4392
rect 576 4392 594 4410
rect 576 4410 594 4428
rect 576 4428 594 4446
rect 576 4446 594 4464
rect 576 4464 594 4482
rect 576 4482 594 4500
rect 576 4500 594 4518
rect 576 4518 594 4536
rect 576 4536 594 4554
rect 576 4554 594 4572
rect 576 4572 594 4590
rect 576 4590 594 4608
rect 576 4608 594 4626
rect 576 4626 594 4644
rect 576 4644 594 4662
rect 576 4662 594 4680
rect 576 4680 594 4698
rect 576 4698 594 4716
rect 576 4716 594 4734
rect 576 4734 594 4752
rect 576 4752 594 4770
rect 576 4770 594 4788
rect 576 4788 594 4806
rect 576 4806 594 4824
rect 576 4824 594 4842
rect 576 4842 594 4860
rect 576 4860 594 4878
rect 576 4878 594 4896
rect 576 4896 594 4914
rect 576 4914 594 4932
rect 576 4932 594 4950
rect 576 4950 594 4968
rect 576 4968 594 4986
rect 576 4986 594 5004
rect 576 5004 594 5022
rect 576 5022 594 5040
rect 576 5040 594 5058
rect 576 5058 594 5076
rect 576 5076 594 5094
rect 576 5094 594 5112
rect 576 5112 594 5130
rect 576 5130 594 5148
rect 576 5148 594 5166
rect 576 5166 594 5184
rect 576 5184 594 5202
rect 576 5202 594 5220
rect 576 5220 594 5238
rect 576 5238 594 5256
rect 576 5256 594 5274
rect 576 5274 594 5292
rect 576 5292 594 5310
rect 576 5310 594 5328
rect 576 5328 594 5346
rect 576 5346 594 5364
rect 576 5364 594 5382
rect 576 5382 594 5400
rect 576 5400 594 5418
rect 576 5418 594 5436
rect 576 5436 594 5454
rect 576 5454 594 5472
rect 576 5472 594 5490
rect 576 5490 594 5508
rect 576 5508 594 5526
rect 576 5526 594 5544
rect 576 5544 594 5562
rect 576 5562 594 5580
rect 576 5580 594 5598
rect 594 1638 612 1656
rect 594 1656 612 1674
rect 594 1674 612 1692
rect 594 1692 612 1710
rect 594 1710 612 1728
rect 594 1728 612 1746
rect 594 1746 612 1764
rect 594 1764 612 1782
rect 594 1782 612 1800
rect 594 1800 612 1818
rect 594 1818 612 1836
rect 594 1836 612 1854
rect 594 1854 612 1872
rect 594 1872 612 1890
rect 594 1890 612 1908
rect 594 1908 612 1926
rect 594 1926 612 1944
rect 594 1944 612 1962
rect 594 1962 612 1980
rect 594 1980 612 1998
rect 594 1998 612 2016
rect 594 2016 612 2034
rect 594 2034 612 2052
rect 594 2052 612 2070
rect 594 2070 612 2088
rect 594 2088 612 2106
rect 594 2106 612 2124
rect 594 2124 612 2142
rect 594 2142 612 2160
rect 594 2160 612 2178
rect 594 2178 612 2196
rect 594 2196 612 2214
rect 594 2214 612 2232
rect 594 2232 612 2250
rect 594 2250 612 2268
rect 594 2268 612 2286
rect 594 2286 612 2304
rect 594 2304 612 2322
rect 594 2322 612 2340
rect 594 2340 612 2358
rect 594 2358 612 2376
rect 594 2376 612 2394
rect 594 2394 612 2412
rect 594 2412 612 2430
rect 594 2430 612 2448
rect 594 2448 612 2466
rect 594 2466 612 2484
rect 594 2484 612 2502
rect 594 2502 612 2520
rect 594 2520 612 2538
rect 594 2538 612 2556
rect 594 2556 612 2574
rect 594 2574 612 2592
rect 594 2592 612 2610
rect 594 2610 612 2628
rect 594 2628 612 2646
rect 594 2646 612 2664
rect 594 2664 612 2682
rect 594 2682 612 2700
rect 594 2700 612 2718
rect 594 2718 612 2736
rect 594 2736 612 2754
rect 594 2754 612 2772
rect 594 2772 612 2790
rect 594 2790 612 2808
rect 594 2808 612 2826
rect 594 2826 612 2844
rect 594 2844 612 2862
rect 594 2862 612 2880
rect 594 2880 612 2898
rect 594 2898 612 2916
rect 594 2916 612 2934
rect 594 2934 612 2952
rect 594 2952 612 2970
rect 594 2970 612 2988
rect 594 2988 612 3006
rect 594 3006 612 3024
rect 594 3024 612 3042
rect 594 3042 612 3060
rect 594 3060 612 3078
rect 594 3078 612 3096
rect 594 3096 612 3114
rect 594 3114 612 3132
rect 594 3132 612 3150
rect 594 3150 612 3168
rect 594 3168 612 3186
rect 594 3186 612 3204
rect 594 3204 612 3222
rect 594 3222 612 3240
rect 594 3240 612 3258
rect 594 3258 612 3276
rect 594 3276 612 3294
rect 594 3294 612 3312
rect 594 3312 612 3330
rect 594 3330 612 3348
rect 594 3348 612 3366
rect 594 3366 612 3384
rect 594 3384 612 3402
rect 594 3402 612 3420
rect 594 3420 612 3438
rect 594 3438 612 3456
rect 594 3456 612 3474
rect 594 3474 612 3492
rect 594 3492 612 3510
rect 594 3510 612 3528
rect 594 3528 612 3546
rect 594 3546 612 3564
rect 594 3564 612 3582
rect 594 3582 612 3600
rect 594 3600 612 3618
rect 594 3618 612 3636
rect 594 3636 612 3654
rect 594 3654 612 3672
rect 594 3672 612 3690
rect 594 3690 612 3708
rect 594 3708 612 3726
rect 594 3726 612 3744
rect 594 3744 612 3762
rect 594 3762 612 3780
rect 594 3780 612 3798
rect 594 3798 612 3816
rect 594 3816 612 3834
rect 594 3834 612 3852
rect 594 3852 612 3870
rect 594 3870 612 3888
rect 594 3888 612 3906
rect 594 3906 612 3924
rect 594 3924 612 3942
rect 594 3942 612 3960
rect 594 3960 612 3978
rect 594 3978 612 3996
rect 594 3996 612 4014
rect 594 4014 612 4032
rect 594 4032 612 4050
rect 594 4050 612 4068
rect 594 4068 612 4086
rect 594 4086 612 4104
rect 594 4104 612 4122
rect 594 4122 612 4140
rect 594 4140 612 4158
rect 594 4158 612 4176
rect 594 4176 612 4194
rect 594 4194 612 4212
rect 594 4212 612 4230
rect 594 4230 612 4248
rect 594 4248 612 4266
rect 594 4266 612 4284
rect 594 4284 612 4302
rect 594 4302 612 4320
rect 594 4320 612 4338
rect 594 4338 612 4356
rect 594 4356 612 4374
rect 594 4374 612 4392
rect 594 4392 612 4410
rect 594 4410 612 4428
rect 594 4428 612 4446
rect 594 4446 612 4464
rect 594 4464 612 4482
rect 594 4482 612 4500
rect 594 4500 612 4518
rect 594 4518 612 4536
rect 594 4536 612 4554
rect 594 4554 612 4572
rect 594 4572 612 4590
rect 594 4590 612 4608
rect 594 4608 612 4626
rect 594 4626 612 4644
rect 594 4644 612 4662
rect 594 4662 612 4680
rect 594 4680 612 4698
rect 594 4698 612 4716
rect 594 4716 612 4734
rect 594 4734 612 4752
rect 594 4752 612 4770
rect 594 4770 612 4788
rect 594 4788 612 4806
rect 594 4806 612 4824
rect 594 4824 612 4842
rect 594 4842 612 4860
rect 594 4860 612 4878
rect 594 4878 612 4896
rect 594 4896 612 4914
rect 594 4914 612 4932
rect 594 4932 612 4950
rect 594 4950 612 4968
rect 594 4968 612 4986
rect 594 4986 612 5004
rect 594 5004 612 5022
rect 594 5022 612 5040
rect 594 5040 612 5058
rect 594 5058 612 5076
rect 594 5076 612 5094
rect 594 5094 612 5112
rect 594 5112 612 5130
rect 594 5130 612 5148
rect 594 5148 612 5166
rect 594 5166 612 5184
rect 594 5184 612 5202
rect 594 5202 612 5220
rect 594 5220 612 5238
rect 594 5238 612 5256
rect 594 5256 612 5274
rect 594 5274 612 5292
rect 594 5292 612 5310
rect 594 5310 612 5328
rect 594 5328 612 5346
rect 594 5346 612 5364
rect 594 5364 612 5382
rect 594 5382 612 5400
rect 594 5400 612 5418
rect 594 5418 612 5436
rect 594 5436 612 5454
rect 594 5454 612 5472
rect 594 5472 612 5490
rect 594 5490 612 5508
rect 594 5508 612 5526
rect 594 5526 612 5544
rect 594 5544 612 5562
rect 594 5562 612 5580
rect 594 5580 612 5598
rect 594 5598 612 5616
rect 594 5616 612 5634
rect 612 1602 630 1620
rect 612 1620 630 1638
rect 612 1638 630 1656
rect 612 1656 630 1674
rect 612 1674 630 1692
rect 612 1692 630 1710
rect 612 1710 630 1728
rect 612 1728 630 1746
rect 612 1746 630 1764
rect 612 1764 630 1782
rect 612 1782 630 1800
rect 612 1800 630 1818
rect 612 1818 630 1836
rect 612 1836 630 1854
rect 612 1854 630 1872
rect 612 1872 630 1890
rect 612 1890 630 1908
rect 612 1908 630 1926
rect 612 1926 630 1944
rect 612 1944 630 1962
rect 612 1962 630 1980
rect 612 1980 630 1998
rect 612 1998 630 2016
rect 612 2016 630 2034
rect 612 2034 630 2052
rect 612 2052 630 2070
rect 612 2070 630 2088
rect 612 2088 630 2106
rect 612 2106 630 2124
rect 612 2124 630 2142
rect 612 2142 630 2160
rect 612 2160 630 2178
rect 612 2178 630 2196
rect 612 2196 630 2214
rect 612 2214 630 2232
rect 612 2232 630 2250
rect 612 2250 630 2268
rect 612 2268 630 2286
rect 612 2286 630 2304
rect 612 2304 630 2322
rect 612 2322 630 2340
rect 612 2340 630 2358
rect 612 2358 630 2376
rect 612 2376 630 2394
rect 612 2394 630 2412
rect 612 2412 630 2430
rect 612 2430 630 2448
rect 612 2448 630 2466
rect 612 2466 630 2484
rect 612 2484 630 2502
rect 612 2502 630 2520
rect 612 2520 630 2538
rect 612 2538 630 2556
rect 612 2556 630 2574
rect 612 2574 630 2592
rect 612 2592 630 2610
rect 612 2610 630 2628
rect 612 2628 630 2646
rect 612 2646 630 2664
rect 612 2664 630 2682
rect 612 2682 630 2700
rect 612 2700 630 2718
rect 612 2718 630 2736
rect 612 2736 630 2754
rect 612 2754 630 2772
rect 612 2772 630 2790
rect 612 2790 630 2808
rect 612 2808 630 2826
rect 612 2826 630 2844
rect 612 2844 630 2862
rect 612 2862 630 2880
rect 612 2880 630 2898
rect 612 2898 630 2916
rect 612 2916 630 2934
rect 612 2934 630 2952
rect 612 2952 630 2970
rect 612 2970 630 2988
rect 612 2988 630 3006
rect 612 3006 630 3024
rect 612 3024 630 3042
rect 612 3042 630 3060
rect 612 3060 630 3078
rect 612 3078 630 3096
rect 612 3096 630 3114
rect 612 3114 630 3132
rect 612 3132 630 3150
rect 612 3150 630 3168
rect 612 3168 630 3186
rect 612 3186 630 3204
rect 612 3204 630 3222
rect 612 3222 630 3240
rect 612 3240 630 3258
rect 612 3258 630 3276
rect 612 3276 630 3294
rect 612 3294 630 3312
rect 612 3312 630 3330
rect 612 3330 630 3348
rect 612 3348 630 3366
rect 612 3366 630 3384
rect 612 3384 630 3402
rect 612 3402 630 3420
rect 612 3420 630 3438
rect 612 3438 630 3456
rect 612 3456 630 3474
rect 612 3474 630 3492
rect 612 3492 630 3510
rect 612 3510 630 3528
rect 612 3528 630 3546
rect 612 3546 630 3564
rect 612 3564 630 3582
rect 612 3582 630 3600
rect 612 3600 630 3618
rect 612 3618 630 3636
rect 612 3636 630 3654
rect 612 3654 630 3672
rect 612 3672 630 3690
rect 612 3690 630 3708
rect 612 3708 630 3726
rect 612 3726 630 3744
rect 612 3744 630 3762
rect 612 3762 630 3780
rect 612 3780 630 3798
rect 612 3798 630 3816
rect 612 3816 630 3834
rect 612 3834 630 3852
rect 612 3852 630 3870
rect 612 3870 630 3888
rect 612 3888 630 3906
rect 612 3906 630 3924
rect 612 3924 630 3942
rect 612 3942 630 3960
rect 612 3960 630 3978
rect 612 3978 630 3996
rect 612 3996 630 4014
rect 612 4014 630 4032
rect 612 4032 630 4050
rect 612 4050 630 4068
rect 612 4068 630 4086
rect 612 4086 630 4104
rect 612 4104 630 4122
rect 612 4122 630 4140
rect 612 4140 630 4158
rect 612 4158 630 4176
rect 612 4176 630 4194
rect 612 4194 630 4212
rect 612 4212 630 4230
rect 612 4230 630 4248
rect 612 4248 630 4266
rect 612 4266 630 4284
rect 612 4284 630 4302
rect 612 4302 630 4320
rect 612 4320 630 4338
rect 612 4338 630 4356
rect 612 4356 630 4374
rect 612 4374 630 4392
rect 612 4392 630 4410
rect 612 4410 630 4428
rect 612 4428 630 4446
rect 612 4446 630 4464
rect 612 4464 630 4482
rect 612 4482 630 4500
rect 612 4500 630 4518
rect 612 4518 630 4536
rect 612 4536 630 4554
rect 612 4554 630 4572
rect 612 4572 630 4590
rect 612 4590 630 4608
rect 612 4608 630 4626
rect 612 4626 630 4644
rect 612 4644 630 4662
rect 612 4662 630 4680
rect 612 4680 630 4698
rect 612 4698 630 4716
rect 612 4716 630 4734
rect 612 4734 630 4752
rect 612 4752 630 4770
rect 612 4770 630 4788
rect 612 4788 630 4806
rect 612 4806 630 4824
rect 612 4824 630 4842
rect 612 4842 630 4860
rect 612 4860 630 4878
rect 612 4878 630 4896
rect 612 4896 630 4914
rect 612 4914 630 4932
rect 612 4932 630 4950
rect 612 4950 630 4968
rect 612 4968 630 4986
rect 612 4986 630 5004
rect 612 5004 630 5022
rect 612 5022 630 5040
rect 612 5040 630 5058
rect 612 5058 630 5076
rect 612 5076 630 5094
rect 612 5094 630 5112
rect 612 5112 630 5130
rect 612 5130 630 5148
rect 612 5148 630 5166
rect 612 5166 630 5184
rect 612 5184 630 5202
rect 612 5202 630 5220
rect 612 5220 630 5238
rect 612 5238 630 5256
rect 612 5256 630 5274
rect 612 5274 630 5292
rect 612 5292 630 5310
rect 612 5310 630 5328
rect 612 5328 630 5346
rect 612 5346 630 5364
rect 612 5364 630 5382
rect 612 5382 630 5400
rect 612 5400 630 5418
rect 612 5418 630 5436
rect 612 5436 630 5454
rect 612 5454 630 5472
rect 612 5472 630 5490
rect 612 5490 630 5508
rect 612 5508 630 5526
rect 612 5526 630 5544
rect 612 5544 630 5562
rect 612 5562 630 5580
rect 612 5580 630 5598
rect 612 5598 630 5616
rect 612 5616 630 5634
rect 612 5634 630 5652
rect 612 5652 630 5670
rect 630 1584 648 1602
rect 630 1602 648 1620
rect 630 1620 648 1638
rect 630 1638 648 1656
rect 630 1656 648 1674
rect 630 1674 648 1692
rect 630 1692 648 1710
rect 630 1710 648 1728
rect 630 1728 648 1746
rect 630 1746 648 1764
rect 630 1764 648 1782
rect 630 1782 648 1800
rect 630 1800 648 1818
rect 630 1818 648 1836
rect 630 1836 648 1854
rect 630 1854 648 1872
rect 630 1872 648 1890
rect 630 1890 648 1908
rect 630 1908 648 1926
rect 630 1926 648 1944
rect 630 1944 648 1962
rect 630 1962 648 1980
rect 630 1980 648 1998
rect 630 1998 648 2016
rect 630 2016 648 2034
rect 630 2034 648 2052
rect 630 2052 648 2070
rect 630 2070 648 2088
rect 630 2088 648 2106
rect 630 2106 648 2124
rect 630 2124 648 2142
rect 630 2142 648 2160
rect 630 2160 648 2178
rect 630 2178 648 2196
rect 630 2196 648 2214
rect 630 2214 648 2232
rect 630 2232 648 2250
rect 630 2250 648 2268
rect 630 2268 648 2286
rect 630 2286 648 2304
rect 630 2304 648 2322
rect 630 2322 648 2340
rect 630 2340 648 2358
rect 630 2358 648 2376
rect 630 2376 648 2394
rect 630 2394 648 2412
rect 630 2412 648 2430
rect 630 2430 648 2448
rect 630 2448 648 2466
rect 630 2466 648 2484
rect 630 2484 648 2502
rect 630 2502 648 2520
rect 630 2520 648 2538
rect 630 2538 648 2556
rect 630 2556 648 2574
rect 630 2574 648 2592
rect 630 2592 648 2610
rect 630 2610 648 2628
rect 630 2628 648 2646
rect 630 2646 648 2664
rect 630 2664 648 2682
rect 630 2682 648 2700
rect 630 2700 648 2718
rect 630 2718 648 2736
rect 630 2736 648 2754
rect 630 2754 648 2772
rect 630 2772 648 2790
rect 630 2790 648 2808
rect 630 2808 648 2826
rect 630 2826 648 2844
rect 630 2844 648 2862
rect 630 2862 648 2880
rect 630 2880 648 2898
rect 630 2898 648 2916
rect 630 2916 648 2934
rect 630 2934 648 2952
rect 630 2952 648 2970
rect 630 2970 648 2988
rect 630 2988 648 3006
rect 630 3006 648 3024
rect 630 3024 648 3042
rect 630 3042 648 3060
rect 630 3060 648 3078
rect 630 3078 648 3096
rect 630 3096 648 3114
rect 630 3114 648 3132
rect 630 3132 648 3150
rect 630 3150 648 3168
rect 630 3168 648 3186
rect 630 3186 648 3204
rect 630 3204 648 3222
rect 630 3222 648 3240
rect 630 3240 648 3258
rect 630 3258 648 3276
rect 630 3276 648 3294
rect 630 3294 648 3312
rect 630 3312 648 3330
rect 630 3330 648 3348
rect 630 3348 648 3366
rect 630 3366 648 3384
rect 630 3384 648 3402
rect 630 3870 648 3888
rect 630 3888 648 3906
rect 630 3906 648 3924
rect 630 3924 648 3942
rect 630 3942 648 3960
rect 630 3960 648 3978
rect 630 3978 648 3996
rect 630 3996 648 4014
rect 630 4014 648 4032
rect 630 4032 648 4050
rect 630 4050 648 4068
rect 630 4068 648 4086
rect 630 4086 648 4104
rect 630 4104 648 4122
rect 630 4122 648 4140
rect 630 4140 648 4158
rect 630 4158 648 4176
rect 630 4176 648 4194
rect 630 4194 648 4212
rect 630 4212 648 4230
rect 630 4230 648 4248
rect 630 4248 648 4266
rect 630 4266 648 4284
rect 630 4284 648 4302
rect 630 4302 648 4320
rect 630 4320 648 4338
rect 630 4338 648 4356
rect 630 4356 648 4374
rect 630 4374 648 4392
rect 630 4392 648 4410
rect 630 4410 648 4428
rect 630 4428 648 4446
rect 630 4446 648 4464
rect 630 4464 648 4482
rect 630 4482 648 4500
rect 630 4500 648 4518
rect 630 4518 648 4536
rect 630 4536 648 4554
rect 630 4554 648 4572
rect 630 4572 648 4590
rect 630 4590 648 4608
rect 630 4608 648 4626
rect 630 4626 648 4644
rect 630 4644 648 4662
rect 630 4662 648 4680
rect 630 4680 648 4698
rect 630 4698 648 4716
rect 630 4716 648 4734
rect 630 4734 648 4752
rect 630 4752 648 4770
rect 630 4770 648 4788
rect 630 4788 648 4806
rect 630 4806 648 4824
rect 630 4824 648 4842
rect 630 4842 648 4860
rect 630 4860 648 4878
rect 630 4878 648 4896
rect 630 4896 648 4914
rect 630 4914 648 4932
rect 630 4932 648 4950
rect 630 4950 648 4968
rect 630 4968 648 4986
rect 630 4986 648 5004
rect 630 5004 648 5022
rect 630 5022 648 5040
rect 630 5040 648 5058
rect 630 5058 648 5076
rect 630 5076 648 5094
rect 630 5094 648 5112
rect 630 5112 648 5130
rect 630 5130 648 5148
rect 630 5148 648 5166
rect 630 5166 648 5184
rect 630 5184 648 5202
rect 630 5202 648 5220
rect 630 5220 648 5238
rect 630 5238 648 5256
rect 630 5256 648 5274
rect 630 5274 648 5292
rect 630 5292 648 5310
rect 630 5310 648 5328
rect 630 5328 648 5346
rect 630 5346 648 5364
rect 630 5364 648 5382
rect 630 5382 648 5400
rect 630 5400 648 5418
rect 630 5418 648 5436
rect 630 5436 648 5454
rect 630 5454 648 5472
rect 630 5472 648 5490
rect 630 5490 648 5508
rect 630 5508 648 5526
rect 630 5526 648 5544
rect 630 5544 648 5562
rect 630 5562 648 5580
rect 630 5580 648 5598
rect 630 5598 648 5616
rect 630 5616 648 5634
rect 630 5634 648 5652
rect 630 5652 648 5670
rect 630 5670 648 5688
rect 648 1548 666 1566
rect 648 1566 666 1584
rect 648 1584 666 1602
rect 648 1602 666 1620
rect 648 1620 666 1638
rect 648 1638 666 1656
rect 648 1656 666 1674
rect 648 1674 666 1692
rect 648 1692 666 1710
rect 648 1710 666 1728
rect 648 1728 666 1746
rect 648 1746 666 1764
rect 648 1764 666 1782
rect 648 1782 666 1800
rect 648 1800 666 1818
rect 648 1818 666 1836
rect 648 1836 666 1854
rect 648 1854 666 1872
rect 648 1872 666 1890
rect 648 1890 666 1908
rect 648 1908 666 1926
rect 648 1926 666 1944
rect 648 1944 666 1962
rect 648 1962 666 1980
rect 648 1980 666 1998
rect 648 1998 666 2016
rect 648 2016 666 2034
rect 648 2034 666 2052
rect 648 2052 666 2070
rect 648 2070 666 2088
rect 648 2088 666 2106
rect 648 2106 666 2124
rect 648 2124 666 2142
rect 648 2142 666 2160
rect 648 2160 666 2178
rect 648 2178 666 2196
rect 648 2196 666 2214
rect 648 2214 666 2232
rect 648 2232 666 2250
rect 648 2250 666 2268
rect 648 2268 666 2286
rect 648 2286 666 2304
rect 648 2304 666 2322
rect 648 2322 666 2340
rect 648 2340 666 2358
rect 648 2358 666 2376
rect 648 2376 666 2394
rect 648 2394 666 2412
rect 648 2412 666 2430
rect 648 2430 666 2448
rect 648 2448 666 2466
rect 648 2466 666 2484
rect 648 2484 666 2502
rect 648 2502 666 2520
rect 648 2520 666 2538
rect 648 2538 666 2556
rect 648 2556 666 2574
rect 648 2574 666 2592
rect 648 2592 666 2610
rect 648 2610 666 2628
rect 648 2628 666 2646
rect 648 2646 666 2664
rect 648 2664 666 2682
rect 648 2682 666 2700
rect 648 2700 666 2718
rect 648 2718 666 2736
rect 648 2736 666 2754
rect 648 2754 666 2772
rect 648 2772 666 2790
rect 648 2790 666 2808
rect 648 2808 666 2826
rect 648 2826 666 2844
rect 648 2844 666 2862
rect 648 2862 666 2880
rect 648 2880 666 2898
rect 648 2898 666 2916
rect 648 2916 666 2934
rect 648 2934 666 2952
rect 648 2952 666 2970
rect 648 2970 666 2988
rect 648 2988 666 3006
rect 648 3006 666 3024
rect 648 3024 666 3042
rect 648 3042 666 3060
rect 648 3060 666 3078
rect 648 3078 666 3096
rect 648 3096 666 3114
rect 648 3114 666 3132
rect 648 3132 666 3150
rect 648 3150 666 3168
rect 648 3168 666 3186
rect 648 3186 666 3204
rect 648 3204 666 3222
rect 648 4032 666 4050
rect 648 4050 666 4068
rect 648 4068 666 4086
rect 648 4086 666 4104
rect 648 4104 666 4122
rect 648 4122 666 4140
rect 648 4140 666 4158
rect 648 4158 666 4176
rect 648 4176 666 4194
rect 648 4194 666 4212
rect 648 4212 666 4230
rect 648 4230 666 4248
rect 648 4248 666 4266
rect 648 4266 666 4284
rect 648 4284 666 4302
rect 648 4302 666 4320
rect 648 4320 666 4338
rect 648 4338 666 4356
rect 648 4356 666 4374
rect 648 4374 666 4392
rect 648 4392 666 4410
rect 648 4410 666 4428
rect 648 4428 666 4446
rect 648 4446 666 4464
rect 648 4464 666 4482
rect 648 4482 666 4500
rect 648 4500 666 4518
rect 648 4518 666 4536
rect 648 4536 666 4554
rect 648 4554 666 4572
rect 648 4572 666 4590
rect 648 4590 666 4608
rect 648 4608 666 4626
rect 648 4626 666 4644
rect 648 4644 666 4662
rect 648 4662 666 4680
rect 648 4680 666 4698
rect 648 4698 666 4716
rect 648 4716 666 4734
rect 648 4734 666 4752
rect 648 4752 666 4770
rect 648 4770 666 4788
rect 648 4788 666 4806
rect 648 4806 666 4824
rect 648 4824 666 4842
rect 648 4842 666 4860
rect 648 4860 666 4878
rect 648 4878 666 4896
rect 648 4896 666 4914
rect 648 4914 666 4932
rect 648 4932 666 4950
rect 648 4950 666 4968
rect 648 4968 666 4986
rect 648 4986 666 5004
rect 648 5004 666 5022
rect 648 5022 666 5040
rect 648 5040 666 5058
rect 648 5058 666 5076
rect 648 5076 666 5094
rect 648 5094 666 5112
rect 648 5112 666 5130
rect 648 5130 666 5148
rect 648 5148 666 5166
rect 648 5166 666 5184
rect 648 5184 666 5202
rect 648 5202 666 5220
rect 648 5220 666 5238
rect 648 5238 666 5256
rect 648 5256 666 5274
rect 648 5274 666 5292
rect 648 5292 666 5310
rect 648 5310 666 5328
rect 648 5328 666 5346
rect 648 5346 666 5364
rect 648 5364 666 5382
rect 648 5382 666 5400
rect 648 5400 666 5418
rect 648 5418 666 5436
rect 648 5436 666 5454
rect 648 5454 666 5472
rect 648 5472 666 5490
rect 648 5490 666 5508
rect 648 5508 666 5526
rect 648 5526 666 5544
rect 648 5544 666 5562
rect 648 5562 666 5580
rect 648 5580 666 5598
rect 648 5598 666 5616
rect 648 5616 666 5634
rect 648 5634 666 5652
rect 648 5652 666 5670
rect 648 5670 666 5688
rect 648 5688 666 5706
rect 666 1530 684 1548
rect 666 1548 684 1566
rect 666 1566 684 1584
rect 666 1584 684 1602
rect 666 1602 684 1620
rect 666 1620 684 1638
rect 666 1638 684 1656
rect 666 1656 684 1674
rect 666 1674 684 1692
rect 666 1692 684 1710
rect 666 1710 684 1728
rect 666 1728 684 1746
rect 666 1746 684 1764
rect 666 1764 684 1782
rect 666 1782 684 1800
rect 666 1800 684 1818
rect 666 1818 684 1836
rect 666 1836 684 1854
rect 666 1854 684 1872
rect 666 1872 684 1890
rect 666 1890 684 1908
rect 666 1908 684 1926
rect 666 1926 684 1944
rect 666 1944 684 1962
rect 666 1962 684 1980
rect 666 1980 684 1998
rect 666 1998 684 2016
rect 666 2016 684 2034
rect 666 2034 684 2052
rect 666 2052 684 2070
rect 666 2070 684 2088
rect 666 2088 684 2106
rect 666 2106 684 2124
rect 666 2124 684 2142
rect 666 2142 684 2160
rect 666 2160 684 2178
rect 666 2178 684 2196
rect 666 2196 684 2214
rect 666 2214 684 2232
rect 666 2232 684 2250
rect 666 2250 684 2268
rect 666 2268 684 2286
rect 666 2286 684 2304
rect 666 2304 684 2322
rect 666 2322 684 2340
rect 666 2340 684 2358
rect 666 2358 684 2376
rect 666 2376 684 2394
rect 666 2394 684 2412
rect 666 2412 684 2430
rect 666 2430 684 2448
rect 666 2448 684 2466
rect 666 2466 684 2484
rect 666 2484 684 2502
rect 666 2502 684 2520
rect 666 2520 684 2538
rect 666 2538 684 2556
rect 666 2556 684 2574
rect 666 2574 684 2592
rect 666 2592 684 2610
rect 666 2610 684 2628
rect 666 2628 684 2646
rect 666 2646 684 2664
rect 666 2664 684 2682
rect 666 2682 684 2700
rect 666 2700 684 2718
rect 666 2718 684 2736
rect 666 2736 684 2754
rect 666 2754 684 2772
rect 666 2772 684 2790
rect 666 2790 684 2808
rect 666 2808 684 2826
rect 666 2826 684 2844
rect 666 2844 684 2862
rect 666 2862 684 2880
rect 666 2880 684 2898
rect 666 2898 684 2916
rect 666 2916 684 2934
rect 666 2934 684 2952
rect 666 2952 684 2970
rect 666 2970 684 2988
rect 666 2988 684 3006
rect 666 3006 684 3024
rect 666 3024 684 3042
rect 666 3042 684 3060
rect 666 3060 684 3078
rect 666 3078 684 3096
rect 666 3096 684 3114
rect 666 4158 684 4176
rect 666 4176 684 4194
rect 666 4194 684 4212
rect 666 4212 684 4230
rect 666 4230 684 4248
rect 666 4248 684 4266
rect 666 4266 684 4284
rect 666 4284 684 4302
rect 666 4302 684 4320
rect 666 4320 684 4338
rect 666 4338 684 4356
rect 666 4356 684 4374
rect 666 4374 684 4392
rect 666 4392 684 4410
rect 666 4410 684 4428
rect 666 4428 684 4446
rect 666 4446 684 4464
rect 666 4464 684 4482
rect 666 4482 684 4500
rect 666 4500 684 4518
rect 666 4518 684 4536
rect 666 4536 684 4554
rect 666 4554 684 4572
rect 666 4572 684 4590
rect 666 4590 684 4608
rect 666 4608 684 4626
rect 666 4626 684 4644
rect 666 4644 684 4662
rect 666 4662 684 4680
rect 666 4680 684 4698
rect 666 4698 684 4716
rect 666 4716 684 4734
rect 666 4734 684 4752
rect 666 4752 684 4770
rect 666 4770 684 4788
rect 666 4788 684 4806
rect 666 4806 684 4824
rect 666 4824 684 4842
rect 666 4842 684 4860
rect 666 4860 684 4878
rect 666 4878 684 4896
rect 666 4896 684 4914
rect 666 4914 684 4932
rect 666 4932 684 4950
rect 666 4950 684 4968
rect 666 4968 684 4986
rect 666 4986 684 5004
rect 666 5004 684 5022
rect 666 5022 684 5040
rect 666 5040 684 5058
rect 666 5058 684 5076
rect 666 5076 684 5094
rect 666 5094 684 5112
rect 666 5112 684 5130
rect 666 5130 684 5148
rect 666 5148 684 5166
rect 666 5166 684 5184
rect 666 5184 684 5202
rect 666 5202 684 5220
rect 666 5220 684 5238
rect 666 5238 684 5256
rect 666 5256 684 5274
rect 666 5274 684 5292
rect 666 5292 684 5310
rect 666 5310 684 5328
rect 666 5328 684 5346
rect 666 5346 684 5364
rect 666 5364 684 5382
rect 666 5382 684 5400
rect 666 5400 684 5418
rect 666 5418 684 5436
rect 666 5436 684 5454
rect 666 5454 684 5472
rect 666 5472 684 5490
rect 666 5490 684 5508
rect 666 5508 684 5526
rect 666 5526 684 5544
rect 666 5544 684 5562
rect 666 5562 684 5580
rect 666 5580 684 5598
rect 666 5598 684 5616
rect 666 5616 684 5634
rect 666 5634 684 5652
rect 666 5652 684 5670
rect 666 5670 684 5688
rect 666 5688 684 5706
rect 666 5706 684 5724
rect 666 5724 684 5742
rect 684 1512 702 1530
rect 684 1530 702 1548
rect 684 1548 702 1566
rect 684 1566 702 1584
rect 684 1584 702 1602
rect 684 1602 702 1620
rect 684 1620 702 1638
rect 684 1638 702 1656
rect 684 1656 702 1674
rect 684 1674 702 1692
rect 684 1692 702 1710
rect 684 1710 702 1728
rect 684 1728 702 1746
rect 684 1746 702 1764
rect 684 1764 702 1782
rect 684 1782 702 1800
rect 684 1800 702 1818
rect 684 1818 702 1836
rect 684 1836 702 1854
rect 684 1854 702 1872
rect 684 1872 702 1890
rect 684 1890 702 1908
rect 684 1908 702 1926
rect 684 1926 702 1944
rect 684 1944 702 1962
rect 684 1962 702 1980
rect 684 1980 702 1998
rect 684 1998 702 2016
rect 684 2016 702 2034
rect 684 2034 702 2052
rect 684 2052 702 2070
rect 684 2070 702 2088
rect 684 2088 702 2106
rect 684 2106 702 2124
rect 684 2124 702 2142
rect 684 2142 702 2160
rect 684 2160 702 2178
rect 684 2178 702 2196
rect 684 2196 702 2214
rect 684 2214 702 2232
rect 684 2232 702 2250
rect 684 2250 702 2268
rect 684 2268 702 2286
rect 684 2286 702 2304
rect 684 2304 702 2322
rect 684 2322 702 2340
rect 684 2340 702 2358
rect 684 2358 702 2376
rect 684 2376 702 2394
rect 684 2394 702 2412
rect 684 2412 702 2430
rect 684 2430 702 2448
rect 684 2448 702 2466
rect 684 2466 702 2484
rect 684 2484 702 2502
rect 684 2502 702 2520
rect 684 2520 702 2538
rect 684 2538 702 2556
rect 684 2556 702 2574
rect 684 2574 702 2592
rect 684 2592 702 2610
rect 684 2610 702 2628
rect 684 2628 702 2646
rect 684 2646 702 2664
rect 684 2664 702 2682
rect 684 2682 702 2700
rect 684 2700 702 2718
rect 684 2718 702 2736
rect 684 2736 702 2754
rect 684 2754 702 2772
rect 684 2772 702 2790
rect 684 2790 702 2808
rect 684 2808 702 2826
rect 684 2826 702 2844
rect 684 2844 702 2862
rect 684 2862 702 2880
rect 684 2880 702 2898
rect 684 2898 702 2916
rect 684 2916 702 2934
rect 684 2934 702 2952
rect 684 2952 702 2970
rect 684 2970 702 2988
rect 684 2988 702 3006
rect 684 3006 702 3024
rect 684 4248 702 4266
rect 684 4266 702 4284
rect 684 4284 702 4302
rect 684 4302 702 4320
rect 684 4320 702 4338
rect 684 4338 702 4356
rect 684 4356 702 4374
rect 684 4374 702 4392
rect 684 4392 702 4410
rect 684 4410 702 4428
rect 684 4428 702 4446
rect 684 4446 702 4464
rect 684 4464 702 4482
rect 684 4482 702 4500
rect 684 4500 702 4518
rect 684 4518 702 4536
rect 684 4536 702 4554
rect 684 4554 702 4572
rect 684 4572 702 4590
rect 684 4590 702 4608
rect 684 4608 702 4626
rect 684 4626 702 4644
rect 684 4644 702 4662
rect 684 4662 702 4680
rect 684 4680 702 4698
rect 684 4698 702 4716
rect 684 4716 702 4734
rect 684 4734 702 4752
rect 684 4752 702 4770
rect 684 4770 702 4788
rect 684 4788 702 4806
rect 684 4806 702 4824
rect 684 4824 702 4842
rect 684 4842 702 4860
rect 684 4860 702 4878
rect 684 4878 702 4896
rect 684 4896 702 4914
rect 684 4914 702 4932
rect 684 4932 702 4950
rect 684 4950 702 4968
rect 684 4968 702 4986
rect 684 4986 702 5004
rect 684 5004 702 5022
rect 684 5022 702 5040
rect 684 5040 702 5058
rect 684 5058 702 5076
rect 684 5076 702 5094
rect 684 5094 702 5112
rect 684 5112 702 5130
rect 684 5130 702 5148
rect 684 5148 702 5166
rect 684 5166 702 5184
rect 684 5184 702 5202
rect 684 5202 702 5220
rect 684 5220 702 5238
rect 684 5238 702 5256
rect 684 5256 702 5274
rect 684 5274 702 5292
rect 684 5292 702 5310
rect 684 5310 702 5328
rect 684 5328 702 5346
rect 684 5346 702 5364
rect 684 5364 702 5382
rect 684 5382 702 5400
rect 684 5400 702 5418
rect 684 5418 702 5436
rect 684 5436 702 5454
rect 684 5454 702 5472
rect 684 5472 702 5490
rect 684 5490 702 5508
rect 684 5508 702 5526
rect 684 5526 702 5544
rect 684 5544 702 5562
rect 684 5562 702 5580
rect 684 5580 702 5598
rect 684 5598 702 5616
rect 684 5616 702 5634
rect 684 5634 702 5652
rect 684 5652 702 5670
rect 684 5670 702 5688
rect 684 5688 702 5706
rect 684 5706 702 5724
rect 684 5724 702 5742
rect 684 5742 702 5760
rect 702 1476 720 1494
rect 702 1494 720 1512
rect 702 1512 720 1530
rect 702 1530 720 1548
rect 702 1548 720 1566
rect 702 1566 720 1584
rect 702 1584 720 1602
rect 702 1602 720 1620
rect 702 1620 720 1638
rect 702 1638 720 1656
rect 702 1656 720 1674
rect 702 1674 720 1692
rect 702 1692 720 1710
rect 702 1710 720 1728
rect 702 1728 720 1746
rect 702 1746 720 1764
rect 702 1764 720 1782
rect 702 1782 720 1800
rect 702 1800 720 1818
rect 702 1818 720 1836
rect 702 1836 720 1854
rect 702 1854 720 1872
rect 702 1872 720 1890
rect 702 1890 720 1908
rect 702 1908 720 1926
rect 702 1926 720 1944
rect 702 1944 720 1962
rect 702 1962 720 1980
rect 702 1980 720 1998
rect 702 1998 720 2016
rect 702 2016 720 2034
rect 702 2034 720 2052
rect 702 2052 720 2070
rect 702 2070 720 2088
rect 702 2088 720 2106
rect 702 2106 720 2124
rect 702 2124 720 2142
rect 702 2142 720 2160
rect 702 2160 720 2178
rect 702 2178 720 2196
rect 702 2196 720 2214
rect 702 2214 720 2232
rect 702 2232 720 2250
rect 702 2250 720 2268
rect 702 2268 720 2286
rect 702 2286 720 2304
rect 702 2304 720 2322
rect 702 2322 720 2340
rect 702 2340 720 2358
rect 702 2358 720 2376
rect 702 2376 720 2394
rect 702 2394 720 2412
rect 702 2412 720 2430
rect 702 2430 720 2448
rect 702 2448 720 2466
rect 702 2466 720 2484
rect 702 2484 720 2502
rect 702 2502 720 2520
rect 702 2520 720 2538
rect 702 2538 720 2556
rect 702 2556 720 2574
rect 702 2574 720 2592
rect 702 2592 720 2610
rect 702 2610 720 2628
rect 702 2628 720 2646
rect 702 2646 720 2664
rect 702 2664 720 2682
rect 702 2682 720 2700
rect 702 2700 720 2718
rect 702 2718 720 2736
rect 702 2736 720 2754
rect 702 2754 720 2772
rect 702 2772 720 2790
rect 702 2790 720 2808
rect 702 2808 720 2826
rect 702 2826 720 2844
rect 702 2844 720 2862
rect 702 2862 720 2880
rect 702 2880 720 2898
rect 702 2898 720 2916
rect 702 2916 720 2934
rect 702 4338 720 4356
rect 702 4356 720 4374
rect 702 4374 720 4392
rect 702 4392 720 4410
rect 702 4410 720 4428
rect 702 4428 720 4446
rect 702 4446 720 4464
rect 702 4464 720 4482
rect 702 4482 720 4500
rect 702 4500 720 4518
rect 702 4518 720 4536
rect 702 4536 720 4554
rect 702 4554 720 4572
rect 702 4572 720 4590
rect 702 4590 720 4608
rect 702 4608 720 4626
rect 702 4626 720 4644
rect 702 4644 720 4662
rect 702 4662 720 4680
rect 702 4680 720 4698
rect 702 4698 720 4716
rect 702 4716 720 4734
rect 702 4734 720 4752
rect 702 4752 720 4770
rect 702 4770 720 4788
rect 702 4788 720 4806
rect 702 4806 720 4824
rect 702 4824 720 4842
rect 702 4842 720 4860
rect 702 4860 720 4878
rect 702 4878 720 4896
rect 702 4896 720 4914
rect 702 4914 720 4932
rect 702 4932 720 4950
rect 702 4950 720 4968
rect 702 4968 720 4986
rect 702 4986 720 5004
rect 702 5004 720 5022
rect 702 5022 720 5040
rect 702 5040 720 5058
rect 702 5058 720 5076
rect 702 5076 720 5094
rect 702 5094 720 5112
rect 702 5112 720 5130
rect 702 5130 720 5148
rect 702 5148 720 5166
rect 702 5166 720 5184
rect 702 5184 720 5202
rect 702 5202 720 5220
rect 702 5220 720 5238
rect 702 5238 720 5256
rect 702 5256 720 5274
rect 702 5274 720 5292
rect 702 5292 720 5310
rect 702 5310 720 5328
rect 702 5328 720 5346
rect 702 5346 720 5364
rect 702 5364 720 5382
rect 702 5382 720 5400
rect 702 5400 720 5418
rect 702 5418 720 5436
rect 702 5436 720 5454
rect 702 5454 720 5472
rect 702 5472 720 5490
rect 702 5490 720 5508
rect 702 5508 720 5526
rect 702 5526 720 5544
rect 702 5544 720 5562
rect 702 5562 720 5580
rect 702 5580 720 5598
rect 702 5598 720 5616
rect 702 5616 720 5634
rect 702 5634 720 5652
rect 702 5652 720 5670
rect 702 5670 720 5688
rect 702 5688 720 5706
rect 702 5706 720 5724
rect 702 5724 720 5742
rect 702 5742 720 5760
rect 702 5760 720 5778
rect 702 5778 720 5796
rect 720 1458 738 1476
rect 720 1476 738 1494
rect 720 1494 738 1512
rect 720 1512 738 1530
rect 720 1530 738 1548
rect 720 1548 738 1566
rect 720 1566 738 1584
rect 720 1584 738 1602
rect 720 1602 738 1620
rect 720 1620 738 1638
rect 720 1638 738 1656
rect 720 1656 738 1674
rect 720 1674 738 1692
rect 720 1692 738 1710
rect 720 1710 738 1728
rect 720 1728 738 1746
rect 720 1746 738 1764
rect 720 1764 738 1782
rect 720 1782 738 1800
rect 720 1800 738 1818
rect 720 1818 738 1836
rect 720 1836 738 1854
rect 720 1854 738 1872
rect 720 1872 738 1890
rect 720 1890 738 1908
rect 720 1908 738 1926
rect 720 1926 738 1944
rect 720 1944 738 1962
rect 720 1962 738 1980
rect 720 1980 738 1998
rect 720 1998 738 2016
rect 720 2016 738 2034
rect 720 2034 738 2052
rect 720 2052 738 2070
rect 720 2070 738 2088
rect 720 2088 738 2106
rect 720 2106 738 2124
rect 720 2124 738 2142
rect 720 2142 738 2160
rect 720 2160 738 2178
rect 720 2178 738 2196
rect 720 2196 738 2214
rect 720 2214 738 2232
rect 720 2232 738 2250
rect 720 2250 738 2268
rect 720 2268 738 2286
rect 720 2286 738 2304
rect 720 2304 738 2322
rect 720 2322 738 2340
rect 720 2340 738 2358
rect 720 2358 738 2376
rect 720 2376 738 2394
rect 720 2394 738 2412
rect 720 2412 738 2430
rect 720 2430 738 2448
rect 720 2448 738 2466
rect 720 2466 738 2484
rect 720 2484 738 2502
rect 720 2502 738 2520
rect 720 2520 738 2538
rect 720 2538 738 2556
rect 720 2556 738 2574
rect 720 2574 738 2592
rect 720 2592 738 2610
rect 720 2610 738 2628
rect 720 2628 738 2646
rect 720 2646 738 2664
rect 720 2664 738 2682
rect 720 2682 738 2700
rect 720 2700 738 2718
rect 720 2718 738 2736
rect 720 2736 738 2754
rect 720 2754 738 2772
rect 720 2772 738 2790
rect 720 2790 738 2808
rect 720 2808 738 2826
rect 720 2826 738 2844
rect 720 2844 738 2862
rect 720 4410 738 4428
rect 720 4428 738 4446
rect 720 4446 738 4464
rect 720 4464 738 4482
rect 720 4482 738 4500
rect 720 4500 738 4518
rect 720 4518 738 4536
rect 720 4536 738 4554
rect 720 4554 738 4572
rect 720 4572 738 4590
rect 720 4590 738 4608
rect 720 4608 738 4626
rect 720 4626 738 4644
rect 720 4644 738 4662
rect 720 4662 738 4680
rect 720 4680 738 4698
rect 720 4698 738 4716
rect 720 4716 738 4734
rect 720 4734 738 4752
rect 720 4752 738 4770
rect 720 4770 738 4788
rect 720 4788 738 4806
rect 720 4806 738 4824
rect 720 4824 738 4842
rect 720 4842 738 4860
rect 720 4860 738 4878
rect 720 4878 738 4896
rect 720 4896 738 4914
rect 720 4914 738 4932
rect 720 4932 738 4950
rect 720 4950 738 4968
rect 720 4968 738 4986
rect 720 4986 738 5004
rect 720 5004 738 5022
rect 720 5022 738 5040
rect 720 5040 738 5058
rect 720 5058 738 5076
rect 720 5076 738 5094
rect 720 5094 738 5112
rect 720 5112 738 5130
rect 720 5130 738 5148
rect 720 5148 738 5166
rect 720 5166 738 5184
rect 720 5184 738 5202
rect 720 5202 738 5220
rect 720 5220 738 5238
rect 720 5238 738 5256
rect 720 5256 738 5274
rect 720 5274 738 5292
rect 720 5292 738 5310
rect 720 5310 738 5328
rect 720 5328 738 5346
rect 720 5346 738 5364
rect 720 5364 738 5382
rect 720 5382 738 5400
rect 720 5400 738 5418
rect 720 5418 738 5436
rect 720 5436 738 5454
rect 720 5454 738 5472
rect 720 5472 738 5490
rect 720 5490 738 5508
rect 720 5508 738 5526
rect 720 5526 738 5544
rect 720 5544 738 5562
rect 720 5562 738 5580
rect 720 5580 738 5598
rect 720 5598 738 5616
rect 720 5616 738 5634
rect 720 5634 738 5652
rect 720 5652 738 5670
rect 720 5670 738 5688
rect 720 5688 738 5706
rect 720 5706 738 5724
rect 720 5724 738 5742
rect 720 5742 738 5760
rect 720 5760 738 5778
rect 720 5778 738 5796
rect 720 5796 738 5814
rect 738 1440 756 1458
rect 738 1458 756 1476
rect 738 1476 756 1494
rect 738 1494 756 1512
rect 738 1512 756 1530
rect 738 1530 756 1548
rect 738 1548 756 1566
rect 738 1566 756 1584
rect 738 1584 756 1602
rect 738 1602 756 1620
rect 738 1620 756 1638
rect 738 1638 756 1656
rect 738 1656 756 1674
rect 738 1674 756 1692
rect 738 1692 756 1710
rect 738 1710 756 1728
rect 738 1728 756 1746
rect 738 1746 756 1764
rect 738 1764 756 1782
rect 738 1782 756 1800
rect 738 1800 756 1818
rect 738 1818 756 1836
rect 738 1836 756 1854
rect 738 1854 756 1872
rect 738 1872 756 1890
rect 738 1890 756 1908
rect 738 1908 756 1926
rect 738 1926 756 1944
rect 738 1944 756 1962
rect 738 1962 756 1980
rect 738 1980 756 1998
rect 738 1998 756 2016
rect 738 2016 756 2034
rect 738 2034 756 2052
rect 738 2052 756 2070
rect 738 2070 756 2088
rect 738 2088 756 2106
rect 738 2106 756 2124
rect 738 2124 756 2142
rect 738 2142 756 2160
rect 738 2160 756 2178
rect 738 2178 756 2196
rect 738 2196 756 2214
rect 738 2214 756 2232
rect 738 2232 756 2250
rect 738 2250 756 2268
rect 738 2268 756 2286
rect 738 2286 756 2304
rect 738 2304 756 2322
rect 738 2322 756 2340
rect 738 2340 756 2358
rect 738 2358 756 2376
rect 738 2376 756 2394
rect 738 2394 756 2412
rect 738 2412 756 2430
rect 738 2430 756 2448
rect 738 2448 756 2466
rect 738 2466 756 2484
rect 738 2484 756 2502
rect 738 2502 756 2520
rect 738 2520 756 2538
rect 738 2538 756 2556
rect 738 2556 756 2574
rect 738 2574 756 2592
rect 738 2592 756 2610
rect 738 2610 756 2628
rect 738 2628 756 2646
rect 738 2646 756 2664
rect 738 2664 756 2682
rect 738 2682 756 2700
rect 738 2700 756 2718
rect 738 2718 756 2736
rect 738 2736 756 2754
rect 738 2754 756 2772
rect 738 2772 756 2790
rect 738 2790 756 2808
rect 738 4464 756 4482
rect 738 4482 756 4500
rect 738 4500 756 4518
rect 738 4518 756 4536
rect 738 4536 756 4554
rect 738 4554 756 4572
rect 738 4572 756 4590
rect 738 4590 756 4608
rect 738 4608 756 4626
rect 738 4626 756 4644
rect 738 4644 756 4662
rect 738 4662 756 4680
rect 738 4680 756 4698
rect 738 4698 756 4716
rect 738 4716 756 4734
rect 738 4734 756 4752
rect 738 4752 756 4770
rect 738 4770 756 4788
rect 738 4788 756 4806
rect 738 4806 756 4824
rect 738 4824 756 4842
rect 738 4842 756 4860
rect 738 4860 756 4878
rect 738 4878 756 4896
rect 738 4896 756 4914
rect 738 4914 756 4932
rect 738 4932 756 4950
rect 738 4950 756 4968
rect 738 4968 756 4986
rect 738 4986 756 5004
rect 738 5004 756 5022
rect 738 5022 756 5040
rect 738 5040 756 5058
rect 738 5058 756 5076
rect 738 5076 756 5094
rect 738 5094 756 5112
rect 738 5112 756 5130
rect 738 5130 756 5148
rect 738 5148 756 5166
rect 738 5166 756 5184
rect 738 5184 756 5202
rect 738 5202 756 5220
rect 738 5220 756 5238
rect 738 5238 756 5256
rect 738 5256 756 5274
rect 738 5274 756 5292
rect 738 5292 756 5310
rect 738 5310 756 5328
rect 738 5328 756 5346
rect 738 5346 756 5364
rect 738 5364 756 5382
rect 738 5382 756 5400
rect 738 5400 756 5418
rect 738 5418 756 5436
rect 738 5436 756 5454
rect 738 5454 756 5472
rect 738 5472 756 5490
rect 738 5490 756 5508
rect 738 5508 756 5526
rect 738 5526 756 5544
rect 738 5544 756 5562
rect 738 5562 756 5580
rect 738 5580 756 5598
rect 738 5598 756 5616
rect 738 5616 756 5634
rect 738 5634 756 5652
rect 738 5652 756 5670
rect 738 5670 756 5688
rect 738 5688 756 5706
rect 738 5706 756 5724
rect 738 5724 756 5742
rect 738 5742 756 5760
rect 738 5760 756 5778
rect 738 5778 756 5796
rect 738 5796 756 5814
rect 738 5814 756 5832
rect 756 1404 774 1422
rect 756 1422 774 1440
rect 756 1440 774 1458
rect 756 1458 774 1476
rect 756 1476 774 1494
rect 756 1494 774 1512
rect 756 1512 774 1530
rect 756 1530 774 1548
rect 756 1548 774 1566
rect 756 1566 774 1584
rect 756 1584 774 1602
rect 756 1602 774 1620
rect 756 1620 774 1638
rect 756 1638 774 1656
rect 756 1656 774 1674
rect 756 1674 774 1692
rect 756 1692 774 1710
rect 756 1710 774 1728
rect 756 1728 774 1746
rect 756 1746 774 1764
rect 756 1764 774 1782
rect 756 1782 774 1800
rect 756 1800 774 1818
rect 756 1818 774 1836
rect 756 1836 774 1854
rect 756 1854 774 1872
rect 756 1872 774 1890
rect 756 1890 774 1908
rect 756 1908 774 1926
rect 756 1926 774 1944
rect 756 1944 774 1962
rect 756 1962 774 1980
rect 756 1980 774 1998
rect 756 1998 774 2016
rect 756 2016 774 2034
rect 756 2034 774 2052
rect 756 2052 774 2070
rect 756 2070 774 2088
rect 756 2088 774 2106
rect 756 2106 774 2124
rect 756 2124 774 2142
rect 756 2142 774 2160
rect 756 2160 774 2178
rect 756 2178 774 2196
rect 756 2196 774 2214
rect 756 2214 774 2232
rect 756 2232 774 2250
rect 756 2250 774 2268
rect 756 2268 774 2286
rect 756 2286 774 2304
rect 756 2304 774 2322
rect 756 2322 774 2340
rect 756 2340 774 2358
rect 756 2358 774 2376
rect 756 2376 774 2394
rect 756 2394 774 2412
rect 756 2412 774 2430
rect 756 2430 774 2448
rect 756 2448 774 2466
rect 756 2466 774 2484
rect 756 2484 774 2502
rect 756 2502 774 2520
rect 756 2520 774 2538
rect 756 2538 774 2556
rect 756 2556 774 2574
rect 756 2574 774 2592
rect 756 2592 774 2610
rect 756 2610 774 2628
rect 756 2628 774 2646
rect 756 2646 774 2664
rect 756 2664 774 2682
rect 756 2682 774 2700
rect 756 2700 774 2718
rect 756 2718 774 2736
rect 756 4536 774 4554
rect 756 4554 774 4572
rect 756 4572 774 4590
rect 756 4590 774 4608
rect 756 4608 774 4626
rect 756 4626 774 4644
rect 756 4644 774 4662
rect 756 4662 774 4680
rect 756 4680 774 4698
rect 756 4698 774 4716
rect 756 4716 774 4734
rect 756 4734 774 4752
rect 756 4752 774 4770
rect 756 4770 774 4788
rect 756 4788 774 4806
rect 756 4806 774 4824
rect 756 4824 774 4842
rect 756 4842 774 4860
rect 756 4860 774 4878
rect 756 4878 774 4896
rect 756 4896 774 4914
rect 756 4914 774 4932
rect 756 4932 774 4950
rect 756 4950 774 4968
rect 756 4968 774 4986
rect 756 4986 774 5004
rect 756 5004 774 5022
rect 756 5022 774 5040
rect 756 5040 774 5058
rect 756 5058 774 5076
rect 756 5076 774 5094
rect 756 5094 774 5112
rect 756 5112 774 5130
rect 756 5130 774 5148
rect 756 5148 774 5166
rect 756 5166 774 5184
rect 756 5184 774 5202
rect 756 5202 774 5220
rect 756 5220 774 5238
rect 756 5238 774 5256
rect 756 5256 774 5274
rect 756 5274 774 5292
rect 756 5292 774 5310
rect 756 5310 774 5328
rect 756 5328 774 5346
rect 756 5346 774 5364
rect 756 5364 774 5382
rect 756 5382 774 5400
rect 756 5400 774 5418
rect 756 5418 774 5436
rect 756 5436 774 5454
rect 756 5454 774 5472
rect 756 5472 774 5490
rect 756 5490 774 5508
rect 756 5508 774 5526
rect 756 5526 774 5544
rect 756 5544 774 5562
rect 756 5562 774 5580
rect 756 5580 774 5598
rect 756 5598 774 5616
rect 756 5616 774 5634
rect 756 5634 774 5652
rect 756 5652 774 5670
rect 756 5670 774 5688
rect 756 5688 774 5706
rect 756 5706 774 5724
rect 756 5724 774 5742
rect 756 5742 774 5760
rect 756 5760 774 5778
rect 756 5778 774 5796
rect 756 5796 774 5814
rect 756 5814 774 5832
rect 756 5832 774 5850
rect 756 5850 774 5868
rect 774 1386 792 1404
rect 774 1404 792 1422
rect 774 1422 792 1440
rect 774 1440 792 1458
rect 774 1458 792 1476
rect 774 1476 792 1494
rect 774 1494 792 1512
rect 774 1512 792 1530
rect 774 1530 792 1548
rect 774 1548 792 1566
rect 774 1566 792 1584
rect 774 1584 792 1602
rect 774 1602 792 1620
rect 774 1620 792 1638
rect 774 1638 792 1656
rect 774 1656 792 1674
rect 774 1674 792 1692
rect 774 1692 792 1710
rect 774 1710 792 1728
rect 774 1728 792 1746
rect 774 1746 792 1764
rect 774 1764 792 1782
rect 774 1782 792 1800
rect 774 1800 792 1818
rect 774 1818 792 1836
rect 774 1836 792 1854
rect 774 1854 792 1872
rect 774 1872 792 1890
rect 774 1890 792 1908
rect 774 1908 792 1926
rect 774 1926 792 1944
rect 774 1944 792 1962
rect 774 1962 792 1980
rect 774 1980 792 1998
rect 774 1998 792 2016
rect 774 2016 792 2034
rect 774 2034 792 2052
rect 774 2052 792 2070
rect 774 2070 792 2088
rect 774 2088 792 2106
rect 774 2106 792 2124
rect 774 2124 792 2142
rect 774 2142 792 2160
rect 774 2160 792 2178
rect 774 2178 792 2196
rect 774 2196 792 2214
rect 774 2214 792 2232
rect 774 2232 792 2250
rect 774 2250 792 2268
rect 774 2268 792 2286
rect 774 2286 792 2304
rect 774 2304 792 2322
rect 774 2322 792 2340
rect 774 2340 792 2358
rect 774 2358 792 2376
rect 774 2376 792 2394
rect 774 2394 792 2412
rect 774 2412 792 2430
rect 774 2430 792 2448
rect 774 2448 792 2466
rect 774 2466 792 2484
rect 774 2484 792 2502
rect 774 2502 792 2520
rect 774 2520 792 2538
rect 774 2538 792 2556
rect 774 2556 792 2574
rect 774 2574 792 2592
rect 774 2592 792 2610
rect 774 2610 792 2628
rect 774 2628 792 2646
rect 774 2646 792 2664
rect 774 2664 792 2682
rect 774 4590 792 4608
rect 774 4608 792 4626
rect 774 4626 792 4644
rect 774 4644 792 4662
rect 774 4662 792 4680
rect 774 4680 792 4698
rect 774 4698 792 4716
rect 774 4716 792 4734
rect 774 4734 792 4752
rect 774 4752 792 4770
rect 774 4770 792 4788
rect 774 4788 792 4806
rect 774 4806 792 4824
rect 774 4824 792 4842
rect 774 4842 792 4860
rect 774 4860 792 4878
rect 774 4878 792 4896
rect 774 4896 792 4914
rect 774 4914 792 4932
rect 774 4932 792 4950
rect 774 4950 792 4968
rect 774 4968 792 4986
rect 774 4986 792 5004
rect 774 5004 792 5022
rect 774 5022 792 5040
rect 774 5040 792 5058
rect 774 5058 792 5076
rect 774 5076 792 5094
rect 774 5094 792 5112
rect 774 5112 792 5130
rect 774 5130 792 5148
rect 774 5148 792 5166
rect 774 5166 792 5184
rect 774 5184 792 5202
rect 774 5202 792 5220
rect 774 5220 792 5238
rect 774 5238 792 5256
rect 774 5256 792 5274
rect 774 5274 792 5292
rect 774 5292 792 5310
rect 774 5310 792 5328
rect 774 5328 792 5346
rect 774 5346 792 5364
rect 774 5364 792 5382
rect 774 5382 792 5400
rect 774 5400 792 5418
rect 774 5418 792 5436
rect 774 5436 792 5454
rect 774 5454 792 5472
rect 774 5472 792 5490
rect 774 5490 792 5508
rect 774 5508 792 5526
rect 774 5526 792 5544
rect 774 5544 792 5562
rect 774 5562 792 5580
rect 774 5580 792 5598
rect 774 5598 792 5616
rect 774 5616 792 5634
rect 774 5634 792 5652
rect 774 5652 792 5670
rect 774 5670 792 5688
rect 774 5688 792 5706
rect 774 5706 792 5724
rect 774 5724 792 5742
rect 774 5742 792 5760
rect 774 5760 792 5778
rect 774 5778 792 5796
rect 774 5796 792 5814
rect 774 5814 792 5832
rect 774 5832 792 5850
rect 774 5850 792 5868
rect 774 5868 792 5886
rect 792 1368 810 1386
rect 792 1386 810 1404
rect 792 1404 810 1422
rect 792 1422 810 1440
rect 792 1440 810 1458
rect 792 1458 810 1476
rect 792 1476 810 1494
rect 792 1494 810 1512
rect 792 1512 810 1530
rect 792 1530 810 1548
rect 792 1548 810 1566
rect 792 1566 810 1584
rect 792 1584 810 1602
rect 792 1602 810 1620
rect 792 1620 810 1638
rect 792 1638 810 1656
rect 792 1656 810 1674
rect 792 1674 810 1692
rect 792 1692 810 1710
rect 792 1710 810 1728
rect 792 1728 810 1746
rect 792 1746 810 1764
rect 792 1764 810 1782
rect 792 1782 810 1800
rect 792 1800 810 1818
rect 792 1818 810 1836
rect 792 1836 810 1854
rect 792 1854 810 1872
rect 792 1872 810 1890
rect 792 1890 810 1908
rect 792 1908 810 1926
rect 792 1926 810 1944
rect 792 1944 810 1962
rect 792 1962 810 1980
rect 792 1980 810 1998
rect 792 1998 810 2016
rect 792 2016 810 2034
rect 792 2034 810 2052
rect 792 2052 810 2070
rect 792 2070 810 2088
rect 792 2088 810 2106
rect 792 2106 810 2124
rect 792 2124 810 2142
rect 792 2142 810 2160
rect 792 2160 810 2178
rect 792 2178 810 2196
rect 792 2196 810 2214
rect 792 2214 810 2232
rect 792 2232 810 2250
rect 792 2250 810 2268
rect 792 2268 810 2286
rect 792 2286 810 2304
rect 792 2304 810 2322
rect 792 2322 810 2340
rect 792 2340 810 2358
rect 792 2358 810 2376
rect 792 2376 810 2394
rect 792 2394 810 2412
rect 792 2412 810 2430
rect 792 2430 810 2448
rect 792 2448 810 2466
rect 792 2466 810 2484
rect 792 2484 810 2502
rect 792 2502 810 2520
rect 792 2520 810 2538
rect 792 2538 810 2556
rect 792 2556 810 2574
rect 792 2574 810 2592
rect 792 2592 810 2610
rect 792 2610 810 2628
rect 792 4644 810 4662
rect 792 4662 810 4680
rect 792 4680 810 4698
rect 792 4698 810 4716
rect 792 4716 810 4734
rect 792 4734 810 4752
rect 792 4752 810 4770
rect 792 4770 810 4788
rect 792 4788 810 4806
rect 792 4806 810 4824
rect 792 4824 810 4842
rect 792 4842 810 4860
rect 792 4860 810 4878
rect 792 4878 810 4896
rect 792 4896 810 4914
rect 792 4914 810 4932
rect 792 4932 810 4950
rect 792 4950 810 4968
rect 792 4968 810 4986
rect 792 4986 810 5004
rect 792 5004 810 5022
rect 792 5022 810 5040
rect 792 5040 810 5058
rect 792 5058 810 5076
rect 792 5076 810 5094
rect 792 5094 810 5112
rect 792 5112 810 5130
rect 792 5130 810 5148
rect 792 5148 810 5166
rect 792 5166 810 5184
rect 792 5184 810 5202
rect 792 5202 810 5220
rect 792 5220 810 5238
rect 792 5238 810 5256
rect 792 5256 810 5274
rect 792 5274 810 5292
rect 792 5292 810 5310
rect 792 5310 810 5328
rect 792 5328 810 5346
rect 792 5346 810 5364
rect 792 5364 810 5382
rect 792 5382 810 5400
rect 792 5400 810 5418
rect 792 5418 810 5436
rect 792 5436 810 5454
rect 792 5454 810 5472
rect 792 5472 810 5490
rect 792 5490 810 5508
rect 792 5508 810 5526
rect 792 5526 810 5544
rect 792 5544 810 5562
rect 792 5562 810 5580
rect 792 5580 810 5598
rect 792 5598 810 5616
rect 792 5616 810 5634
rect 792 5634 810 5652
rect 792 5652 810 5670
rect 792 5670 810 5688
rect 792 5688 810 5706
rect 792 5706 810 5724
rect 792 5724 810 5742
rect 792 5742 810 5760
rect 792 5760 810 5778
rect 792 5778 810 5796
rect 792 5796 810 5814
rect 792 5814 810 5832
rect 792 5832 810 5850
rect 792 5850 810 5868
rect 792 5868 810 5886
rect 792 5886 810 5904
rect 810 1332 828 1350
rect 810 1350 828 1368
rect 810 1368 828 1386
rect 810 1386 828 1404
rect 810 1404 828 1422
rect 810 1422 828 1440
rect 810 1440 828 1458
rect 810 1458 828 1476
rect 810 1476 828 1494
rect 810 1494 828 1512
rect 810 1512 828 1530
rect 810 1530 828 1548
rect 810 1548 828 1566
rect 810 1566 828 1584
rect 810 1584 828 1602
rect 810 1602 828 1620
rect 810 1620 828 1638
rect 810 1638 828 1656
rect 810 1656 828 1674
rect 810 1674 828 1692
rect 810 1692 828 1710
rect 810 1710 828 1728
rect 810 1728 828 1746
rect 810 1746 828 1764
rect 810 1764 828 1782
rect 810 1782 828 1800
rect 810 1800 828 1818
rect 810 1818 828 1836
rect 810 1836 828 1854
rect 810 1854 828 1872
rect 810 1872 828 1890
rect 810 1890 828 1908
rect 810 1908 828 1926
rect 810 1926 828 1944
rect 810 1944 828 1962
rect 810 1962 828 1980
rect 810 1980 828 1998
rect 810 1998 828 2016
rect 810 2016 828 2034
rect 810 2034 828 2052
rect 810 2052 828 2070
rect 810 2070 828 2088
rect 810 2088 828 2106
rect 810 2106 828 2124
rect 810 2124 828 2142
rect 810 2142 828 2160
rect 810 2160 828 2178
rect 810 2178 828 2196
rect 810 2196 828 2214
rect 810 2214 828 2232
rect 810 2232 828 2250
rect 810 2250 828 2268
rect 810 2268 828 2286
rect 810 2286 828 2304
rect 810 2304 828 2322
rect 810 2322 828 2340
rect 810 2340 828 2358
rect 810 2358 828 2376
rect 810 2376 828 2394
rect 810 2394 828 2412
rect 810 2412 828 2430
rect 810 2430 828 2448
rect 810 2448 828 2466
rect 810 2466 828 2484
rect 810 2484 828 2502
rect 810 2502 828 2520
rect 810 2520 828 2538
rect 810 2538 828 2556
rect 810 2556 828 2574
rect 810 2574 828 2592
rect 810 4680 828 4698
rect 810 4698 828 4716
rect 810 4716 828 4734
rect 810 4734 828 4752
rect 810 4752 828 4770
rect 810 4770 828 4788
rect 810 4788 828 4806
rect 810 4806 828 4824
rect 810 4824 828 4842
rect 810 4842 828 4860
rect 810 4860 828 4878
rect 810 4878 828 4896
rect 810 4896 828 4914
rect 810 4914 828 4932
rect 810 4932 828 4950
rect 810 4950 828 4968
rect 810 4968 828 4986
rect 810 4986 828 5004
rect 810 5004 828 5022
rect 810 5022 828 5040
rect 810 5040 828 5058
rect 810 5058 828 5076
rect 810 5076 828 5094
rect 810 5094 828 5112
rect 810 5112 828 5130
rect 810 5130 828 5148
rect 810 5148 828 5166
rect 810 5166 828 5184
rect 810 5184 828 5202
rect 810 5202 828 5220
rect 810 5220 828 5238
rect 810 5238 828 5256
rect 810 5256 828 5274
rect 810 5274 828 5292
rect 810 5292 828 5310
rect 810 5310 828 5328
rect 810 5328 828 5346
rect 810 5346 828 5364
rect 810 5364 828 5382
rect 810 5382 828 5400
rect 810 5400 828 5418
rect 810 5418 828 5436
rect 810 5436 828 5454
rect 810 5454 828 5472
rect 810 5472 828 5490
rect 810 5490 828 5508
rect 810 5508 828 5526
rect 810 5526 828 5544
rect 810 5544 828 5562
rect 810 5562 828 5580
rect 810 5580 828 5598
rect 810 5598 828 5616
rect 810 5616 828 5634
rect 810 5634 828 5652
rect 810 5652 828 5670
rect 810 5670 828 5688
rect 810 5688 828 5706
rect 810 5706 828 5724
rect 810 5724 828 5742
rect 810 5742 828 5760
rect 810 5760 828 5778
rect 810 5778 828 5796
rect 810 5796 828 5814
rect 810 5814 828 5832
rect 810 5832 828 5850
rect 810 5850 828 5868
rect 810 5868 828 5886
rect 810 5886 828 5904
rect 810 5904 828 5922
rect 828 1314 846 1332
rect 828 1332 846 1350
rect 828 1350 846 1368
rect 828 1368 846 1386
rect 828 1386 846 1404
rect 828 1404 846 1422
rect 828 1422 846 1440
rect 828 1440 846 1458
rect 828 1458 846 1476
rect 828 1476 846 1494
rect 828 1494 846 1512
rect 828 1512 846 1530
rect 828 1530 846 1548
rect 828 1548 846 1566
rect 828 1566 846 1584
rect 828 1584 846 1602
rect 828 1602 846 1620
rect 828 1620 846 1638
rect 828 1638 846 1656
rect 828 1656 846 1674
rect 828 1674 846 1692
rect 828 1692 846 1710
rect 828 1710 846 1728
rect 828 1728 846 1746
rect 828 1746 846 1764
rect 828 1764 846 1782
rect 828 1782 846 1800
rect 828 1800 846 1818
rect 828 1818 846 1836
rect 828 1836 846 1854
rect 828 1854 846 1872
rect 828 1872 846 1890
rect 828 1890 846 1908
rect 828 1908 846 1926
rect 828 1926 846 1944
rect 828 1944 846 1962
rect 828 1962 846 1980
rect 828 1980 846 1998
rect 828 1998 846 2016
rect 828 2016 846 2034
rect 828 2034 846 2052
rect 828 2052 846 2070
rect 828 2070 846 2088
rect 828 2088 846 2106
rect 828 2106 846 2124
rect 828 2124 846 2142
rect 828 2142 846 2160
rect 828 2160 846 2178
rect 828 2178 846 2196
rect 828 2196 846 2214
rect 828 2214 846 2232
rect 828 2232 846 2250
rect 828 2250 846 2268
rect 828 2268 846 2286
rect 828 2286 846 2304
rect 828 2304 846 2322
rect 828 2322 846 2340
rect 828 2340 846 2358
rect 828 2358 846 2376
rect 828 2376 846 2394
rect 828 2394 846 2412
rect 828 2412 846 2430
rect 828 2430 846 2448
rect 828 2448 846 2466
rect 828 2466 846 2484
rect 828 2484 846 2502
rect 828 2502 846 2520
rect 828 2520 846 2538
rect 828 4734 846 4752
rect 828 4752 846 4770
rect 828 4770 846 4788
rect 828 4788 846 4806
rect 828 4806 846 4824
rect 828 4824 846 4842
rect 828 4842 846 4860
rect 828 4860 846 4878
rect 828 4878 846 4896
rect 828 4896 846 4914
rect 828 4914 846 4932
rect 828 4932 846 4950
rect 828 4950 846 4968
rect 828 4968 846 4986
rect 828 4986 846 5004
rect 828 5004 846 5022
rect 828 5022 846 5040
rect 828 5040 846 5058
rect 828 5058 846 5076
rect 828 5076 846 5094
rect 828 5094 846 5112
rect 828 5112 846 5130
rect 828 5130 846 5148
rect 828 5148 846 5166
rect 828 5166 846 5184
rect 828 5184 846 5202
rect 828 5202 846 5220
rect 828 5220 846 5238
rect 828 5238 846 5256
rect 828 5256 846 5274
rect 828 5274 846 5292
rect 828 5292 846 5310
rect 828 5310 846 5328
rect 828 5328 846 5346
rect 828 5346 846 5364
rect 828 5364 846 5382
rect 828 5382 846 5400
rect 828 5400 846 5418
rect 828 5418 846 5436
rect 828 5436 846 5454
rect 828 5454 846 5472
rect 828 5472 846 5490
rect 828 5490 846 5508
rect 828 5508 846 5526
rect 828 5526 846 5544
rect 828 5544 846 5562
rect 828 5562 846 5580
rect 828 5580 846 5598
rect 828 5598 846 5616
rect 828 5616 846 5634
rect 828 5634 846 5652
rect 828 5652 846 5670
rect 828 5670 846 5688
rect 828 5688 846 5706
rect 828 5706 846 5724
rect 828 5724 846 5742
rect 828 5742 846 5760
rect 828 5760 846 5778
rect 828 5778 846 5796
rect 828 5796 846 5814
rect 828 5814 846 5832
rect 828 5832 846 5850
rect 828 5850 846 5868
rect 828 5868 846 5886
rect 828 5886 846 5904
rect 828 5904 846 5922
rect 828 5922 846 5940
rect 828 5940 846 5958
rect 846 1296 864 1314
rect 846 1314 864 1332
rect 846 1332 864 1350
rect 846 1350 864 1368
rect 846 1368 864 1386
rect 846 1386 864 1404
rect 846 1404 864 1422
rect 846 1422 864 1440
rect 846 1440 864 1458
rect 846 1458 864 1476
rect 846 1476 864 1494
rect 846 1494 864 1512
rect 846 1512 864 1530
rect 846 1530 864 1548
rect 846 1548 864 1566
rect 846 1566 864 1584
rect 846 1584 864 1602
rect 846 1602 864 1620
rect 846 1620 864 1638
rect 846 1638 864 1656
rect 846 1656 864 1674
rect 846 1674 864 1692
rect 846 1692 864 1710
rect 846 1710 864 1728
rect 846 1728 864 1746
rect 846 1746 864 1764
rect 846 1764 864 1782
rect 846 1782 864 1800
rect 846 1800 864 1818
rect 846 1818 864 1836
rect 846 1836 864 1854
rect 846 1854 864 1872
rect 846 1872 864 1890
rect 846 1890 864 1908
rect 846 1908 864 1926
rect 846 1926 864 1944
rect 846 1944 864 1962
rect 846 1962 864 1980
rect 846 1980 864 1998
rect 846 1998 864 2016
rect 846 2016 864 2034
rect 846 2034 864 2052
rect 846 2052 864 2070
rect 846 2070 864 2088
rect 846 2088 864 2106
rect 846 2106 864 2124
rect 846 2124 864 2142
rect 846 2142 864 2160
rect 846 2160 864 2178
rect 846 2178 864 2196
rect 846 2196 864 2214
rect 846 2214 864 2232
rect 846 2232 864 2250
rect 846 2250 864 2268
rect 846 2268 864 2286
rect 846 2286 864 2304
rect 846 2304 864 2322
rect 846 2322 864 2340
rect 846 2340 864 2358
rect 846 2358 864 2376
rect 846 2376 864 2394
rect 846 2394 864 2412
rect 846 2412 864 2430
rect 846 2430 864 2448
rect 846 2448 864 2466
rect 846 2466 864 2484
rect 846 4788 864 4806
rect 846 4806 864 4824
rect 846 4824 864 4842
rect 846 4842 864 4860
rect 846 4860 864 4878
rect 846 4878 864 4896
rect 846 4896 864 4914
rect 846 4914 864 4932
rect 846 4932 864 4950
rect 846 4950 864 4968
rect 846 4968 864 4986
rect 846 4986 864 5004
rect 846 5004 864 5022
rect 846 5022 864 5040
rect 846 5040 864 5058
rect 846 5058 864 5076
rect 846 5076 864 5094
rect 846 5094 864 5112
rect 846 5112 864 5130
rect 846 5130 864 5148
rect 846 5148 864 5166
rect 846 5166 864 5184
rect 846 5184 864 5202
rect 846 5202 864 5220
rect 846 5220 864 5238
rect 846 5238 864 5256
rect 846 5256 864 5274
rect 846 5274 864 5292
rect 846 5292 864 5310
rect 846 5310 864 5328
rect 846 5328 864 5346
rect 846 5346 864 5364
rect 846 5364 864 5382
rect 846 5382 864 5400
rect 846 5400 864 5418
rect 846 5418 864 5436
rect 846 5436 864 5454
rect 846 5454 864 5472
rect 846 5472 864 5490
rect 846 5490 864 5508
rect 846 5508 864 5526
rect 846 5526 864 5544
rect 846 5544 864 5562
rect 846 5562 864 5580
rect 846 5580 864 5598
rect 846 5598 864 5616
rect 846 5616 864 5634
rect 846 5634 864 5652
rect 846 5652 864 5670
rect 846 5670 864 5688
rect 846 5688 864 5706
rect 846 5706 864 5724
rect 846 5724 864 5742
rect 846 5742 864 5760
rect 846 5760 864 5778
rect 846 5778 864 5796
rect 846 5796 864 5814
rect 846 5814 864 5832
rect 846 5832 864 5850
rect 846 5850 864 5868
rect 846 5868 864 5886
rect 846 5886 864 5904
rect 846 5904 864 5922
rect 846 5922 864 5940
rect 846 5940 864 5958
rect 846 5958 864 5976
rect 864 1278 882 1296
rect 864 1296 882 1314
rect 864 1314 882 1332
rect 864 1332 882 1350
rect 864 1350 882 1368
rect 864 1368 882 1386
rect 864 1386 882 1404
rect 864 1404 882 1422
rect 864 1422 882 1440
rect 864 1440 882 1458
rect 864 1458 882 1476
rect 864 1476 882 1494
rect 864 1494 882 1512
rect 864 1512 882 1530
rect 864 1530 882 1548
rect 864 1548 882 1566
rect 864 1566 882 1584
rect 864 1584 882 1602
rect 864 1602 882 1620
rect 864 1620 882 1638
rect 864 1638 882 1656
rect 864 1656 882 1674
rect 864 1674 882 1692
rect 864 1692 882 1710
rect 864 1710 882 1728
rect 864 1728 882 1746
rect 864 1746 882 1764
rect 864 1764 882 1782
rect 864 1782 882 1800
rect 864 1800 882 1818
rect 864 1818 882 1836
rect 864 1836 882 1854
rect 864 1854 882 1872
rect 864 1872 882 1890
rect 864 1890 882 1908
rect 864 1908 882 1926
rect 864 1926 882 1944
rect 864 1944 882 1962
rect 864 1962 882 1980
rect 864 1980 882 1998
rect 864 1998 882 2016
rect 864 2016 882 2034
rect 864 2034 882 2052
rect 864 2052 882 2070
rect 864 2070 882 2088
rect 864 2088 882 2106
rect 864 2106 882 2124
rect 864 2124 882 2142
rect 864 2142 882 2160
rect 864 2160 882 2178
rect 864 2178 882 2196
rect 864 2196 882 2214
rect 864 2214 882 2232
rect 864 2232 882 2250
rect 864 2250 882 2268
rect 864 2268 882 2286
rect 864 2286 882 2304
rect 864 2304 882 2322
rect 864 2322 882 2340
rect 864 2340 882 2358
rect 864 2358 882 2376
rect 864 2376 882 2394
rect 864 2394 882 2412
rect 864 2412 882 2430
rect 864 2430 882 2448
rect 864 4824 882 4842
rect 864 4842 882 4860
rect 864 4860 882 4878
rect 864 4878 882 4896
rect 864 4896 882 4914
rect 864 4914 882 4932
rect 864 4932 882 4950
rect 864 4950 882 4968
rect 864 4968 882 4986
rect 864 4986 882 5004
rect 864 5004 882 5022
rect 864 5022 882 5040
rect 864 5040 882 5058
rect 864 5058 882 5076
rect 864 5076 882 5094
rect 864 5094 882 5112
rect 864 5112 882 5130
rect 864 5130 882 5148
rect 864 5148 882 5166
rect 864 5166 882 5184
rect 864 5184 882 5202
rect 864 5202 882 5220
rect 864 5220 882 5238
rect 864 5238 882 5256
rect 864 5256 882 5274
rect 864 5274 882 5292
rect 864 5292 882 5310
rect 864 5310 882 5328
rect 864 5328 882 5346
rect 864 5346 882 5364
rect 864 5364 882 5382
rect 864 5382 882 5400
rect 864 5400 882 5418
rect 864 5418 882 5436
rect 864 5436 882 5454
rect 864 5454 882 5472
rect 864 5472 882 5490
rect 864 5490 882 5508
rect 864 5508 882 5526
rect 864 5526 882 5544
rect 864 5544 882 5562
rect 864 5562 882 5580
rect 864 5580 882 5598
rect 864 5598 882 5616
rect 864 5616 882 5634
rect 864 5634 882 5652
rect 864 5652 882 5670
rect 864 5670 882 5688
rect 864 5688 882 5706
rect 864 5706 882 5724
rect 864 5724 882 5742
rect 864 5742 882 5760
rect 864 5760 882 5778
rect 864 5778 882 5796
rect 864 5796 882 5814
rect 864 5814 882 5832
rect 864 5832 882 5850
rect 864 5850 882 5868
rect 864 5868 882 5886
rect 864 5886 882 5904
rect 864 5904 882 5922
rect 864 5922 882 5940
rect 864 5940 882 5958
rect 864 5958 882 5976
rect 864 5976 882 5994
rect 882 1260 900 1278
rect 882 1278 900 1296
rect 882 1296 900 1314
rect 882 1314 900 1332
rect 882 1332 900 1350
rect 882 1350 900 1368
rect 882 1368 900 1386
rect 882 1386 900 1404
rect 882 1404 900 1422
rect 882 1422 900 1440
rect 882 1440 900 1458
rect 882 1458 900 1476
rect 882 1476 900 1494
rect 882 1494 900 1512
rect 882 1512 900 1530
rect 882 1530 900 1548
rect 882 1548 900 1566
rect 882 1566 900 1584
rect 882 1584 900 1602
rect 882 1602 900 1620
rect 882 1620 900 1638
rect 882 1638 900 1656
rect 882 1656 900 1674
rect 882 1674 900 1692
rect 882 1692 900 1710
rect 882 1710 900 1728
rect 882 1728 900 1746
rect 882 1746 900 1764
rect 882 1764 900 1782
rect 882 1782 900 1800
rect 882 1800 900 1818
rect 882 1818 900 1836
rect 882 1836 900 1854
rect 882 1854 900 1872
rect 882 1872 900 1890
rect 882 1890 900 1908
rect 882 1908 900 1926
rect 882 1926 900 1944
rect 882 1944 900 1962
rect 882 1962 900 1980
rect 882 1980 900 1998
rect 882 1998 900 2016
rect 882 2016 900 2034
rect 882 2034 900 2052
rect 882 2052 900 2070
rect 882 2070 900 2088
rect 882 2088 900 2106
rect 882 2106 900 2124
rect 882 2124 900 2142
rect 882 2142 900 2160
rect 882 2160 900 2178
rect 882 2178 900 2196
rect 882 2196 900 2214
rect 882 2214 900 2232
rect 882 2232 900 2250
rect 882 2250 900 2268
rect 882 2268 900 2286
rect 882 2286 900 2304
rect 882 2304 900 2322
rect 882 2322 900 2340
rect 882 2340 900 2358
rect 882 2358 900 2376
rect 882 2376 900 2394
rect 882 2394 900 2412
rect 882 4860 900 4878
rect 882 4878 900 4896
rect 882 4896 900 4914
rect 882 4914 900 4932
rect 882 4932 900 4950
rect 882 4950 900 4968
rect 882 4968 900 4986
rect 882 4986 900 5004
rect 882 5004 900 5022
rect 882 5022 900 5040
rect 882 5040 900 5058
rect 882 5058 900 5076
rect 882 5076 900 5094
rect 882 5094 900 5112
rect 882 5112 900 5130
rect 882 5130 900 5148
rect 882 5148 900 5166
rect 882 5166 900 5184
rect 882 5184 900 5202
rect 882 5202 900 5220
rect 882 5220 900 5238
rect 882 5238 900 5256
rect 882 5256 900 5274
rect 882 5274 900 5292
rect 882 5292 900 5310
rect 882 5310 900 5328
rect 882 5328 900 5346
rect 882 5346 900 5364
rect 882 5364 900 5382
rect 882 5382 900 5400
rect 882 5400 900 5418
rect 882 5418 900 5436
rect 882 5436 900 5454
rect 882 5454 900 5472
rect 882 5472 900 5490
rect 882 5490 900 5508
rect 882 5508 900 5526
rect 882 5526 900 5544
rect 882 5544 900 5562
rect 882 5562 900 5580
rect 882 5580 900 5598
rect 882 5598 900 5616
rect 882 5616 900 5634
rect 882 5634 900 5652
rect 882 5652 900 5670
rect 882 5670 900 5688
rect 882 5688 900 5706
rect 882 5706 900 5724
rect 882 5724 900 5742
rect 882 5742 900 5760
rect 882 5760 900 5778
rect 882 5778 900 5796
rect 882 5796 900 5814
rect 882 5814 900 5832
rect 882 5832 900 5850
rect 882 5850 900 5868
rect 882 5868 900 5886
rect 882 5886 900 5904
rect 882 5904 900 5922
rect 882 5922 900 5940
rect 882 5940 900 5958
rect 882 5958 900 5976
rect 882 5976 900 5994
rect 882 5994 900 6012
rect 900 1242 918 1260
rect 900 1260 918 1278
rect 900 1278 918 1296
rect 900 1296 918 1314
rect 900 1314 918 1332
rect 900 1332 918 1350
rect 900 1350 918 1368
rect 900 1368 918 1386
rect 900 1386 918 1404
rect 900 1404 918 1422
rect 900 1422 918 1440
rect 900 1440 918 1458
rect 900 1458 918 1476
rect 900 1476 918 1494
rect 900 1494 918 1512
rect 900 1512 918 1530
rect 900 1530 918 1548
rect 900 1548 918 1566
rect 900 1566 918 1584
rect 900 1584 918 1602
rect 900 1602 918 1620
rect 900 1620 918 1638
rect 900 1638 918 1656
rect 900 1656 918 1674
rect 900 1674 918 1692
rect 900 1692 918 1710
rect 900 1710 918 1728
rect 900 1728 918 1746
rect 900 1746 918 1764
rect 900 1764 918 1782
rect 900 1782 918 1800
rect 900 1800 918 1818
rect 900 1818 918 1836
rect 900 1836 918 1854
rect 900 1854 918 1872
rect 900 1872 918 1890
rect 900 1890 918 1908
rect 900 1908 918 1926
rect 900 1926 918 1944
rect 900 1944 918 1962
rect 900 1962 918 1980
rect 900 1980 918 1998
rect 900 1998 918 2016
rect 900 2016 918 2034
rect 900 2034 918 2052
rect 900 2052 918 2070
rect 900 2070 918 2088
rect 900 2088 918 2106
rect 900 2106 918 2124
rect 900 2124 918 2142
rect 900 2142 918 2160
rect 900 2160 918 2178
rect 900 2178 918 2196
rect 900 2196 918 2214
rect 900 2214 918 2232
rect 900 2232 918 2250
rect 900 2250 918 2268
rect 900 2268 918 2286
rect 900 2286 918 2304
rect 900 2304 918 2322
rect 900 2322 918 2340
rect 900 2340 918 2358
rect 900 2358 918 2376
rect 900 4896 918 4914
rect 900 4914 918 4932
rect 900 4932 918 4950
rect 900 4950 918 4968
rect 900 4968 918 4986
rect 900 4986 918 5004
rect 900 5004 918 5022
rect 900 5022 918 5040
rect 900 5040 918 5058
rect 900 5058 918 5076
rect 900 5076 918 5094
rect 900 5094 918 5112
rect 900 5112 918 5130
rect 900 5130 918 5148
rect 900 5148 918 5166
rect 900 5166 918 5184
rect 900 5184 918 5202
rect 900 5202 918 5220
rect 900 5220 918 5238
rect 900 5238 918 5256
rect 900 5256 918 5274
rect 900 5274 918 5292
rect 900 5292 918 5310
rect 900 5310 918 5328
rect 900 5328 918 5346
rect 900 5346 918 5364
rect 900 5364 918 5382
rect 900 5382 918 5400
rect 900 5400 918 5418
rect 900 5418 918 5436
rect 900 5436 918 5454
rect 900 5454 918 5472
rect 900 5472 918 5490
rect 900 5490 918 5508
rect 900 5508 918 5526
rect 900 5526 918 5544
rect 900 5544 918 5562
rect 900 5562 918 5580
rect 900 5580 918 5598
rect 900 5598 918 5616
rect 900 5616 918 5634
rect 900 5634 918 5652
rect 900 5652 918 5670
rect 900 5670 918 5688
rect 900 5688 918 5706
rect 900 5706 918 5724
rect 900 5724 918 5742
rect 900 5742 918 5760
rect 900 5760 918 5778
rect 900 5778 918 5796
rect 900 5796 918 5814
rect 900 5814 918 5832
rect 900 5832 918 5850
rect 900 5850 918 5868
rect 900 5868 918 5886
rect 900 5886 918 5904
rect 900 5904 918 5922
rect 900 5922 918 5940
rect 900 5940 918 5958
rect 900 5958 918 5976
rect 900 5976 918 5994
rect 900 5994 918 6012
rect 900 6012 918 6030
rect 918 1206 936 1224
rect 918 1224 936 1242
rect 918 1242 936 1260
rect 918 1260 936 1278
rect 918 1278 936 1296
rect 918 1296 936 1314
rect 918 1314 936 1332
rect 918 1332 936 1350
rect 918 1350 936 1368
rect 918 1368 936 1386
rect 918 1386 936 1404
rect 918 1404 936 1422
rect 918 1422 936 1440
rect 918 1440 936 1458
rect 918 1458 936 1476
rect 918 1476 936 1494
rect 918 1494 936 1512
rect 918 1512 936 1530
rect 918 1530 936 1548
rect 918 1548 936 1566
rect 918 1566 936 1584
rect 918 1584 936 1602
rect 918 1602 936 1620
rect 918 1620 936 1638
rect 918 1638 936 1656
rect 918 1656 936 1674
rect 918 1674 936 1692
rect 918 1692 936 1710
rect 918 1710 936 1728
rect 918 1728 936 1746
rect 918 1746 936 1764
rect 918 1764 936 1782
rect 918 1782 936 1800
rect 918 1800 936 1818
rect 918 1818 936 1836
rect 918 1836 936 1854
rect 918 1854 936 1872
rect 918 1872 936 1890
rect 918 1890 936 1908
rect 918 1908 936 1926
rect 918 1926 936 1944
rect 918 1944 936 1962
rect 918 1962 936 1980
rect 918 1980 936 1998
rect 918 1998 936 2016
rect 918 2016 936 2034
rect 918 2034 936 2052
rect 918 2052 936 2070
rect 918 2070 936 2088
rect 918 2088 936 2106
rect 918 2106 936 2124
rect 918 2124 936 2142
rect 918 2142 936 2160
rect 918 2160 936 2178
rect 918 2178 936 2196
rect 918 2196 936 2214
rect 918 2214 936 2232
rect 918 2232 936 2250
rect 918 2250 936 2268
rect 918 2268 936 2286
rect 918 2286 936 2304
rect 918 2304 936 2322
rect 918 4932 936 4950
rect 918 4950 936 4968
rect 918 4968 936 4986
rect 918 4986 936 5004
rect 918 5004 936 5022
rect 918 5022 936 5040
rect 918 5040 936 5058
rect 918 5058 936 5076
rect 918 5076 936 5094
rect 918 5094 936 5112
rect 918 5112 936 5130
rect 918 5130 936 5148
rect 918 5148 936 5166
rect 918 5166 936 5184
rect 918 5184 936 5202
rect 918 5202 936 5220
rect 918 5220 936 5238
rect 918 5238 936 5256
rect 918 5256 936 5274
rect 918 5274 936 5292
rect 918 5292 936 5310
rect 918 5310 936 5328
rect 918 5328 936 5346
rect 918 5346 936 5364
rect 918 5364 936 5382
rect 918 5382 936 5400
rect 918 5400 936 5418
rect 918 5418 936 5436
rect 918 5436 936 5454
rect 918 5454 936 5472
rect 918 5472 936 5490
rect 918 5490 936 5508
rect 918 5508 936 5526
rect 918 5526 936 5544
rect 918 5544 936 5562
rect 918 5562 936 5580
rect 918 5580 936 5598
rect 918 5598 936 5616
rect 918 5616 936 5634
rect 918 5634 936 5652
rect 918 5652 936 5670
rect 918 5670 936 5688
rect 918 5688 936 5706
rect 918 5706 936 5724
rect 918 5724 936 5742
rect 918 5742 936 5760
rect 918 5760 936 5778
rect 918 5778 936 5796
rect 918 5796 936 5814
rect 918 5814 936 5832
rect 918 5832 936 5850
rect 918 5850 936 5868
rect 918 5868 936 5886
rect 918 5886 936 5904
rect 918 5904 936 5922
rect 918 5922 936 5940
rect 918 5940 936 5958
rect 918 5958 936 5976
rect 918 5976 936 5994
rect 918 5994 936 6012
rect 918 6012 936 6030
rect 918 6030 936 6048
rect 936 1188 954 1206
rect 936 1206 954 1224
rect 936 1224 954 1242
rect 936 1242 954 1260
rect 936 1260 954 1278
rect 936 1278 954 1296
rect 936 1296 954 1314
rect 936 1314 954 1332
rect 936 1332 954 1350
rect 936 1350 954 1368
rect 936 1368 954 1386
rect 936 1386 954 1404
rect 936 1404 954 1422
rect 936 1422 954 1440
rect 936 1440 954 1458
rect 936 1458 954 1476
rect 936 1476 954 1494
rect 936 1494 954 1512
rect 936 1512 954 1530
rect 936 1530 954 1548
rect 936 1548 954 1566
rect 936 1566 954 1584
rect 936 1584 954 1602
rect 936 1602 954 1620
rect 936 1620 954 1638
rect 936 1638 954 1656
rect 936 1656 954 1674
rect 936 1674 954 1692
rect 936 1692 954 1710
rect 936 1710 954 1728
rect 936 1728 954 1746
rect 936 1746 954 1764
rect 936 1764 954 1782
rect 936 1782 954 1800
rect 936 1800 954 1818
rect 936 1818 954 1836
rect 936 1836 954 1854
rect 936 1854 954 1872
rect 936 1872 954 1890
rect 936 1890 954 1908
rect 936 1908 954 1926
rect 936 1926 954 1944
rect 936 1944 954 1962
rect 936 1962 954 1980
rect 936 1980 954 1998
rect 936 1998 954 2016
rect 936 2016 954 2034
rect 936 2034 954 2052
rect 936 2052 954 2070
rect 936 2070 954 2088
rect 936 2088 954 2106
rect 936 2106 954 2124
rect 936 2124 954 2142
rect 936 2142 954 2160
rect 936 2160 954 2178
rect 936 2178 954 2196
rect 936 2196 954 2214
rect 936 2214 954 2232
rect 936 2232 954 2250
rect 936 2250 954 2268
rect 936 2268 954 2286
rect 936 4968 954 4986
rect 936 4986 954 5004
rect 936 5004 954 5022
rect 936 5022 954 5040
rect 936 5040 954 5058
rect 936 5058 954 5076
rect 936 5076 954 5094
rect 936 5094 954 5112
rect 936 5112 954 5130
rect 936 5130 954 5148
rect 936 5148 954 5166
rect 936 5166 954 5184
rect 936 5184 954 5202
rect 936 5202 954 5220
rect 936 5220 954 5238
rect 936 5238 954 5256
rect 936 5256 954 5274
rect 936 5274 954 5292
rect 936 5292 954 5310
rect 936 5310 954 5328
rect 936 5328 954 5346
rect 936 5346 954 5364
rect 936 5364 954 5382
rect 936 5382 954 5400
rect 936 5400 954 5418
rect 936 5418 954 5436
rect 936 5436 954 5454
rect 936 5454 954 5472
rect 936 5472 954 5490
rect 936 5490 954 5508
rect 936 5508 954 5526
rect 936 5526 954 5544
rect 936 5544 954 5562
rect 936 5562 954 5580
rect 936 5580 954 5598
rect 936 5598 954 5616
rect 936 5616 954 5634
rect 936 5634 954 5652
rect 936 5652 954 5670
rect 936 5670 954 5688
rect 936 5688 954 5706
rect 936 5706 954 5724
rect 936 5724 954 5742
rect 936 5742 954 5760
rect 936 5760 954 5778
rect 936 5778 954 5796
rect 936 5796 954 5814
rect 936 5814 954 5832
rect 936 5832 954 5850
rect 936 5850 954 5868
rect 936 5868 954 5886
rect 936 5886 954 5904
rect 936 5904 954 5922
rect 936 5922 954 5940
rect 936 5940 954 5958
rect 936 5958 954 5976
rect 936 5976 954 5994
rect 936 5994 954 6012
rect 936 6012 954 6030
rect 936 6030 954 6048
rect 936 6048 954 6066
rect 936 6066 954 6084
rect 954 1170 972 1188
rect 954 1188 972 1206
rect 954 1206 972 1224
rect 954 1224 972 1242
rect 954 1242 972 1260
rect 954 1260 972 1278
rect 954 1278 972 1296
rect 954 1296 972 1314
rect 954 1314 972 1332
rect 954 1332 972 1350
rect 954 1350 972 1368
rect 954 1368 972 1386
rect 954 1386 972 1404
rect 954 1404 972 1422
rect 954 1422 972 1440
rect 954 1440 972 1458
rect 954 1458 972 1476
rect 954 1476 972 1494
rect 954 1494 972 1512
rect 954 1512 972 1530
rect 954 1530 972 1548
rect 954 1548 972 1566
rect 954 1566 972 1584
rect 954 1584 972 1602
rect 954 1602 972 1620
rect 954 1620 972 1638
rect 954 1638 972 1656
rect 954 1656 972 1674
rect 954 1674 972 1692
rect 954 1692 972 1710
rect 954 1710 972 1728
rect 954 1728 972 1746
rect 954 1746 972 1764
rect 954 1764 972 1782
rect 954 1782 972 1800
rect 954 1800 972 1818
rect 954 1818 972 1836
rect 954 1836 972 1854
rect 954 1854 972 1872
rect 954 1872 972 1890
rect 954 1890 972 1908
rect 954 1908 972 1926
rect 954 1926 972 1944
rect 954 1944 972 1962
rect 954 1962 972 1980
rect 954 1980 972 1998
rect 954 1998 972 2016
rect 954 2016 972 2034
rect 954 2034 972 2052
rect 954 2052 972 2070
rect 954 2070 972 2088
rect 954 2088 972 2106
rect 954 2106 972 2124
rect 954 2124 972 2142
rect 954 2142 972 2160
rect 954 2160 972 2178
rect 954 2178 972 2196
rect 954 2196 972 2214
rect 954 2214 972 2232
rect 954 2232 972 2250
rect 954 5004 972 5022
rect 954 5022 972 5040
rect 954 5040 972 5058
rect 954 5058 972 5076
rect 954 5076 972 5094
rect 954 5094 972 5112
rect 954 5112 972 5130
rect 954 5130 972 5148
rect 954 5148 972 5166
rect 954 5166 972 5184
rect 954 5184 972 5202
rect 954 5202 972 5220
rect 954 5220 972 5238
rect 954 5238 972 5256
rect 954 5256 972 5274
rect 954 5274 972 5292
rect 954 5292 972 5310
rect 954 5310 972 5328
rect 954 5328 972 5346
rect 954 5346 972 5364
rect 954 5364 972 5382
rect 954 5382 972 5400
rect 954 5400 972 5418
rect 954 5418 972 5436
rect 954 5436 972 5454
rect 954 5454 972 5472
rect 954 5472 972 5490
rect 954 5490 972 5508
rect 954 5508 972 5526
rect 954 5526 972 5544
rect 954 5544 972 5562
rect 954 5562 972 5580
rect 954 5580 972 5598
rect 954 5598 972 5616
rect 954 5616 972 5634
rect 954 5634 972 5652
rect 954 5652 972 5670
rect 954 5670 972 5688
rect 954 5688 972 5706
rect 954 5706 972 5724
rect 954 5724 972 5742
rect 954 5742 972 5760
rect 954 5760 972 5778
rect 954 5778 972 5796
rect 954 5796 972 5814
rect 954 5814 972 5832
rect 954 5832 972 5850
rect 954 5850 972 5868
rect 954 5868 972 5886
rect 954 5886 972 5904
rect 954 5904 972 5922
rect 954 5922 972 5940
rect 954 5940 972 5958
rect 954 5958 972 5976
rect 954 5976 972 5994
rect 954 5994 972 6012
rect 954 6012 972 6030
rect 954 6030 972 6048
rect 954 6048 972 6066
rect 954 6066 972 6084
rect 954 6084 972 6102
rect 972 1152 990 1170
rect 972 1170 990 1188
rect 972 1188 990 1206
rect 972 1206 990 1224
rect 972 1224 990 1242
rect 972 1242 990 1260
rect 972 1260 990 1278
rect 972 1278 990 1296
rect 972 1296 990 1314
rect 972 1314 990 1332
rect 972 1332 990 1350
rect 972 1350 990 1368
rect 972 1368 990 1386
rect 972 1386 990 1404
rect 972 1404 990 1422
rect 972 1422 990 1440
rect 972 1440 990 1458
rect 972 1458 990 1476
rect 972 1476 990 1494
rect 972 1494 990 1512
rect 972 1512 990 1530
rect 972 1530 990 1548
rect 972 1548 990 1566
rect 972 1566 990 1584
rect 972 1584 990 1602
rect 972 1602 990 1620
rect 972 1620 990 1638
rect 972 1638 990 1656
rect 972 1656 990 1674
rect 972 1674 990 1692
rect 972 1692 990 1710
rect 972 1710 990 1728
rect 972 1728 990 1746
rect 972 1746 990 1764
rect 972 1764 990 1782
rect 972 1782 990 1800
rect 972 1800 990 1818
rect 972 1818 990 1836
rect 972 1836 990 1854
rect 972 1854 990 1872
rect 972 1872 990 1890
rect 972 1890 990 1908
rect 972 1908 990 1926
rect 972 1926 990 1944
rect 972 1944 990 1962
rect 972 1962 990 1980
rect 972 1980 990 1998
rect 972 1998 990 2016
rect 972 2016 990 2034
rect 972 2034 990 2052
rect 972 2052 990 2070
rect 972 2070 990 2088
rect 972 2088 990 2106
rect 972 2106 990 2124
rect 972 2124 990 2142
rect 972 2142 990 2160
rect 972 2160 990 2178
rect 972 2178 990 2196
rect 972 2196 990 2214
rect 972 5040 990 5058
rect 972 5058 990 5076
rect 972 5076 990 5094
rect 972 5094 990 5112
rect 972 5112 990 5130
rect 972 5130 990 5148
rect 972 5148 990 5166
rect 972 5166 990 5184
rect 972 5184 990 5202
rect 972 5202 990 5220
rect 972 5220 990 5238
rect 972 5238 990 5256
rect 972 5256 990 5274
rect 972 5274 990 5292
rect 972 5292 990 5310
rect 972 5310 990 5328
rect 972 5328 990 5346
rect 972 5346 990 5364
rect 972 5364 990 5382
rect 972 5382 990 5400
rect 972 5400 990 5418
rect 972 5418 990 5436
rect 972 5436 990 5454
rect 972 5454 990 5472
rect 972 5472 990 5490
rect 972 5490 990 5508
rect 972 5508 990 5526
rect 972 5526 990 5544
rect 972 5544 990 5562
rect 972 5562 990 5580
rect 972 5580 990 5598
rect 972 5598 990 5616
rect 972 5616 990 5634
rect 972 5634 990 5652
rect 972 5652 990 5670
rect 972 5670 990 5688
rect 972 5688 990 5706
rect 972 5706 990 5724
rect 972 5724 990 5742
rect 972 5742 990 5760
rect 972 5760 990 5778
rect 972 5778 990 5796
rect 972 5796 990 5814
rect 972 5814 990 5832
rect 972 5832 990 5850
rect 972 5850 990 5868
rect 972 5868 990 5886
rect 972 5886 990 5904
rect 972 5904 990 5922
rect 972 5922 990 5940
rect 972 5940 990 5958
rect 972 5958 990 5976
rect 972 5976 990 5994
rect 972 5994 990 6012
rect 972 6012 990 6030
rect 972 6030 990 6048
rect 972 6048 990 6066
rect 972 6066 990 6084
rect 972 6084 990 6102
rect 972 6102 990 6120
rect 990 1134 1008 1152
rect 990 1152 1008 1170
rect 990 1170 1008 1188
rect 990 1188 1008 1206
rect 990 1206 1008 1224
rect 990 1224 1008 1242
rect 990 1242 1008 1260
rect 990 1260 1008 1278
rect 990 1278 1008 1296
rect 990 1296 1008 1314
rect 990 1314 1008 1332
rect 990 1332 1008 1350
rect 990 1350 1008 1368
rect 990 1368 1008 1386
rect 990 1386 1008 1404
rect 990 1404 1008 1422
rect 990 1422 1008 1440
rect 990 1440 1008 1458
rect 990 1458 1008 1476
rect 990 1476 1008 1494
rect 990 1494 1008 1512
rect 990 1512 1008 1530
rect 990 1530 1008 1548
rect 990 1548 1008 1566
rect 990 1566 1008 1584
rect 990 1584 1008 1602
rect 990 1602 1008 1620
rect 990 1620 1008 1638
rect 990 1638 1008 1656
rect 990 1656 1008 1674
rect 990 1674 1008 1692
rect 990 1692 1008 1710
rect 990 1710 1008 1728
rect 990 1728 1008 1746
rect 990 1746 1008 1764
rect 990 1764 1008 1782
rect 990 1782 1008 1800
rect 990 1800 1008 1818
rect 990 1818 1008 1836
rect 990 1836 1008 1854
rect 990 1854 1008 1872
rect 990 1872 1008 1890
rect 990 1890 1008 1908
rect 990 1908 1008 1926
rect 990 1926 1008 1944
rect 990 1944 1008 1962
rect 990 1962 1008 1980
rect 990 1980 1008 1998
rect 990 1998 1008 2016
rect 990 2016 1008 2034
rect 990 2034 1008 2052
rect 990 2052 1008 2070
rect 990 2070 1008 2088
rect 990 2088 1008 2106
rect 990 2106 1008 2124
rect 990 2124 1008 2142
rect 990 2142 1008 2160
rect 990 2160 1008 2178
rect 990 2178 1008 2196
rect 990 5076 1008 5094
rect 990 5094 1008 5112
rect 990 5112 1008 5130
rect 990 5130 1008 5148
rect 990 5148 1008 5166
rect 990 5166 1008 5184
rect 990 5184 1008 5202
rect 990 5202 1008 5220
rect 990 5220 1008 5238
rect 990 5238 1008 5256
rect 990 5256 1008 5274
rect 990 5274 1008 5292
rect 990 5292 1008 5310
rect 990 5310 1008 5328
rect 990 5328 1008 5346
rect 990 5346 1008 5364
rect 990 5364 1008 5382
rect 990 5382 1008 5400
rect 990 5400 1008 5418
rect 990 5418 1008 5436
rect 990 5436 1008 5454
rect 990 5454 1008 5472
rect 990 5472 1008 5490
rect 990 5490 1008 5508
rect 990 5508 1008 5526
rect 990 5526 1008 5544
rect 990 5544 1008 5562
rect 990 5562 1008 5580
rect 990 5580 1008 5598
rect 990 5598 1008 5616
rect 990 5616 1008 5634
rect 990 5634 1008 5652
rect 990 5652 1008 5670
rect 990 5670 1008 5688
rect 990 5688 1008 5706
rect 990 5706 1008 5724
rect 990 5724 1008 5742
rect 990 5742 1008 5760
rect 990 5760 1008 5778
rect 990 5778 1008 5796
rect 990 5796 1008 5814
rect 990 5814 1008 5832
rect 990 5832 1008 5850
rect 990 5850 1008 5868
rect 990 5868 1008 5886
rect 990 5886 1008 5904
rect 990 5904 1008 5922
rect 990 5922 1008 5940
rect 990 5940 1008 5958
rect 990 5958 1008 5976
rect 990 5976 1008 5994
rect 990 5994 1008 6012
rect 990 6012 1008 6030
rect 990 6030 1008 6048
rect 990 6048 1008 6066
rect 990 6066 1008 6084
rect 990 6084 1008 6102
rect 990 6102 1008 6120
rect 990 6120 1008 6138
rect 1008 1116 1026 1134
rect 1008 1134 1026 1152
rect 1008 1152 1026 1170
rect 1008 1170 1026 1188
rect 1008 1188 1026 1206
rect 1008 1206 1026 1224
rect 1008 1224 1026 1242
rect 1008 1242 1026 1260
rect 1008 1260 1026 1278
rect 1008 1278 1026 1296
rect 1008 1296 1026 1314
rect 1008 1314 1026 1332
rect 1008 1332 1026 1350
rect 1008 1350 1026 1368
rect 1008 1368 1026 1386
rect 1008 1386 1026 1404
rect 1008 1404 1026 1422
rect 1008 1422 1026 1440
rect 1008 1440 1026 1458
rect 1008 1458 1026 1476
rect 1008 1476 1026 1494
rect 1008 1494 1026 1512
rect 1008 1512 1026 1530
rect 1008 1530 1026 1548
rect 1008 1548 1026 1566
rect 1008 1566 1026 1584
rect 1008 1584 1026 1602
rect 1008 1602 1026 1620
rect 1008 1620 1026 1638
rect 1008 1638 1026 1656
rect 1008 1656 1026 1674
rect 1008 1674 1026 1692
rect 1008 1692 1026 1710
rect 1008 1710 1026 1728
rect 1008 1728 1026 1746
rect 1008 1746 1026 1764
rect 1008 1764 1026 1782
rect 1008 1782 1026 1800
rect 1008 1800 1026 1818
rect 1008 1818 1026 1836
rect 1008 1836 1026 1854
rect 1008 1854 1026 1872
rect 1008 1872 1026 1890
rect 1008 1890 1026 1908
rect 1008 1908 1026 1926
rect 1008 1926 1026 1944
rect 1008 1944 1026 1962
rect 1008 1962 1026 1980
rect 1008 1980 1026 1998
rect 1008 1998 1026 2016
rect 1008 2016 1026 2034
rect 1008 2034 1026 2052
rect 1008 2052 1026 2070
rect 1008 2070 1026 2088
rect 1008 2088 1026 2106
rect 1008 2106 1026 2124
rect 1008 2124 1026 2142
rect 1008 2142 1026 2160
rect 1008 5112 1026 5130
rect 1008 5130 1026 5148
rect 1008 5148 1026 5166
rect 1008 5166 1026 5184
rect 1008 5184 1026 5202
rect 1008 5202 1026 5220
rect 1008 5220 1026 5238
rect 1008 5238 1026 5256
rect 1008 5256 1026 5274
rect 1008 5274 1026 5292
rect 1008 5292 1026 5310
rect 1008 5310 1026 5328
rect 1008 5328 1026 5346
rect 1008 5346 1026 5364
rect 1008 5364 1026 5382
rect 1008 5382 1026 5400
rect 1008 5400 1026 5418
rect 1008 5418 1026 5436
rect 1008 5436 1026 5454
rect 1008 5454 1026 5472
rect 1008 5472 1026 5490
rect 1008 5490 1026 5508
rect 1008 5508 1026 5526
rect 1008 5526 1026 5544
rect 1008 5544 1026 5562
rect 1008 5562 1026 5580
rect 1008 5580 1026 5598
rect 1008 5598 1026 5616
rect 1008 5616 1026 5634
rect 1008 5634 1026 5652
rect 1008 5652 1026 5670
rect 1008 5670 1026 5688
rect 1008 5688 1026 5706
rect 1008 5706 1026 5724
rect 1008 5724 1026 5742
rect 1008 5742 1026 5760
rect 1008 5760 1026 5778
rect 1008 5778 1026 5796
rect 1008 5796 1026 5814
rect 1008 5814 1026 5832
rect 1008 5832 1026 5850
rect 1008 5850 1026 5868
rect 1008 5868 1026 5886
rect 1008 5886 1026 5904
rect 1008 5904 1026 5922
rect 1008 5922 1026 5940
rect 1008 5940 1026 5958
rect 1008 5958 1026 5976
rect 1008 5976 1026 5994
rect 1008 5994 1026 6012
rect 1008 6012 1026 6030
rect 1008 6030 1026 6048
rect 1008 6048 1026 6066
rect 1008 6066 1026 6084
rect 1008 6084 1026 6102
rect 1008 6102 1026 6120
rect 1008 6120 1026 6138
rect 1008 6138 1026 6156
rect 1026 1098 1044 1116
rect 1026 1116 1044 1134
rect 1026 1134 1044 1152
rect 1026 1152 1044 1170
rect 1026 1170 1044 1188
rect 1026 1188 1044 1206
rect 1026 1206 1044 1224
rect 1026 1224 1044 1242
rect 1026 1242 1044 1260
rect 1026 1260 1044 1278
rect 1026 1278 1044 1296
rect 1026 1296 1044 1314
rect 1026 1314 1044 1332
rect 1026 1332 1044 1350
rect 1026 1350 1044 1368
rect 1026 1368 1044 1386
rect 1026 1386 1044 1404
rect 1026 1404 1044 1422
rect 1026 1422 1044 1440
rect 1026 1440 1044 1458
rect 1026 1458 1044 1476
rect 1026 1476 1044 1494
rect 1026 1494 1044 1512
rect 1026 1512 1044 1530
rect 1026 1530 1044 1548
rect 1026 1548 1044 1566
rect 1026 1566 1044 1584
rect 1026 1584 1044 1602
rect 1026 1602 1044 1620
rect 1026 1620 1044 1638
rect 1026 1638 1044 1656
rect 1026 1656 1044 1674
rect 1026 1674 1044 1692
rect 1026 1692 1044 1710
rect 1026 1710 1044 1728
rect 1026 1728 1044 1746
rect 1026 1746 1044 1764
rect 1026 1764 1044 1782
rect 1026 1782 1044 1800
rect 1026 1800 1044 1818
rect 1026 1818 1044 1836
rect 1026 1836 1044 1854
rect 1026 1854 1044 1872
rect 1026 1872 1044 1890
rect 1026 1890 1044 1908
rect 1026 1908 1044 1926
rect 1026 1926 1044 1944
rect 1026 1944 1044 1962
rect 1026 1962 1044 1980
rect 1026 1980 1044 1998
rect 1026 1998 1044 2016
rect 1026 2016 1044 2034
rect 1026 2034 1044 2052
rect 1026 2052 1044 2070
rect 1026 2070 1044 2088
rect 1026 2088 1044 2106
rect 1026 2106 1044 2124
rect 1026 5148 1044 5166
rect 1026 5166 1044 5184
rect 1026 5184 1044 5202
rect 1026 5202 1044 5220
rect 1026 5220 1044 5238
rect 1026 5238 1044 5256
rect 1026 5256 1044 5274
rect 1026 5274 1044 5292
rect 1026 5292 1044 5310
rect 1026 5310 1044 5328
rect 1026 5328 1044 5346
rect 1026 5346 1044 5364
rect 1026 5364 1044 5382
rect 1026 5382 1044 5400
rect 1026 5400 1044 5418
rect 1026 5418 1044 5436
rect 1026 5436 1044 5454
rect 1026 5454 1044 5472
rect 1026 5472 1044 5490
rect 1026 5490 1044 5508
rect 1026 5508 1044 5526
rect 1026 5526 1044 5544
rect 1026 5544 1044 5562
rect 1026 5562 1044 5580
rect 1026 5580 1044 5598
rect 1026 5598 1044 5616
rect 1026 5616 1044 5634
rect 1026 5634 1044 5652
rect 1026 5652 1044 5670
rect 1026 5670 1044 5688
rect 1026 5688 1044 5706
rect 1026 5706 1044 5724
rect 1026 5724 1044 5742
rect 1026 5742 1044 5760
rect 1026 5760 1044 5778
rect 1026 5778 1044 5796
rect 1026 5796 1044 5814
rect 1026 5814 1044 5832
rect 1026 5832 1044 5850
rect 1026 5850 1044 5868
rect 1026 5868 1044 5886
rect 1026 5886 1044 5904
rect 1026 5904 1044 5922
rect 1026 5922 1044 5940
rect 1026 5940 1044 5958
rect 1026 5958 1044 5976
rect 1026 5976 1044 5994
rect 1026 5994 1044 6012
rect 1026 6012 1044 6030
rect 1026 6030 1044 6048
rect 1026 6048 1044 6066
rect 1026 6066 1044 6084
rect 1026 6084 1044 6102
rect 1026 6102 1044 6120
rect 1026 6120 1044 6138
rect 1026 6138 1044 6156
rect 1026 6156 1044 6174
rect 1044 1080 1062 1098
rect 1044 1098 1062 1116
rect 1044 1116 1062 1134
rect 1044 1134 1062 1152
rect 1044 1152 1062 1170
rect 1044 1170 1062 1188
rect 1044 1188 1062 1206
rect 1044 1206 1062 1224
rect 1044 1224 1062 1242
rect 1044 1242 1062 1260
rect 1044 1260 1062 1278
rect 1044 1278 1062 1296
rect 1044 1296 1062 1314
rect 1044 1314 1062 1332
rect 1044 1332 1062 1350
rect 1044 1350 1062 1368
rect 1044 1368 1062 1386
rect 1044 1386 1062 1404
rect 1044 1404 1062 1422
rect 1044 1422 1062 1440
rect 1044 1440 1062 1458
rect 1044 1458 1062 1476
rect 1044 1476 1062 1494
rect 1044 1494 1062 1512
rect 1044 1512 1062 1530
rect 1044 1530 1062 1548
rect 1044 1548 1062 1566
rect 1044 1566 1062 1584
rect 1044 1584 1062 1602
rect 1044 1602 1062 1620
rect 1044 1620 1062 1638
rect 1044 1638 1062 1656
rect 1044 1656 1062 1674
rect 1044 1674 1062 1692
rect 1044 1692 1062 1710
rect 1044 1710 1062 1728
rect 1044 1728 1062 1746
rect 1044 1746 1062 1764
rect 1044 1764 1062 1782
rect 1044 1782 1062 1800
rect 1044 1800 1062 1818
rect 1044 1818 1062 1836
rect 1044 1836 1062 1854
rect 1044 1854 1062 1872
rect 1044 1872 1062 1890
rect 1044 1890 1062 1908
rect 1044 1908 1062 1926
rect 1044 1926 1062 1944
rect 1044 1944 1062 1962
rect 1044 1962 1062 1980
rect 1044 1980 1062 1998
rect 1044 1998 1062 2016
rect 1044 2016 1062 2034
rect 1044 2034 1062 2052
rect 1044 2052 1062 2070
rect 1044 2070 1062 2088
rect 1044 5184 1062 5202
rect 1044 5202 1062 5220
rect 1044 5220 1062 5238
rect 1044 5238 1062 5256
rect 1044 5256 1062 5274
rect 1044 5274 1062 5292
rect 1044 5292 1062 5310
rect 1044 5310 1062 5328
rect 1044 5328 1062 5346
rect 1044 5346 1062 5364
rect 1044 5364 1062 5382
rect 1044 5382 1062 5400
rect 1044 5400 1062 5418
rect 1044 5418 1062 5436
rect 1044 5436 1062 5454
rect 1044 5454 1062 5472
rect 1044 5472 1062 5490
rect 1044 5490 1062 5508
rect 1044 5508 1062 5526
rect 1044 5526 1062 5544
rect 1044 5544 1062 5562
rect 1044 5562 1062 5580
rect 1044 5580 1062 5598
rect 1044 5598 1062 5616
rect 1044 5616 1062 5634
rect 1044 5634 1062 5652
rect 1044 5652 1062 5670
rect 1044 5670 1062 5688
rect 1044 5688 1062 5706
rect 1044 5706 1062 5724
rect 1044 5724 1062 5742
rect 1044 5742 1062 5760
rect 1044 5760 1062 5778
rect 1044 5778 1062 5796
rect 1044 5796 1062 5814
rect 1044 5814 1062 5832
rect 1044 5832 1062 5850
rect 1044 5850 1062 5868
rect 1044 5868 1062 5886
rect 1044 5886 1062 5904
rect 1044 5904 1062 5922
rect 1044 5922 1062 5940
rect 1044 5940 1062 5958
rect 1044 5958 1062 5976
rect 1044 5976 1062 5994
rect 1044 5994 1062 6012
rect 1044 6012 1062 6030
rect 1044 6030 1062 6048
rect 1044 6048 1062 6066
rect 1044 6066 1062 6084
rect 1044 6084 1062 6102
rect 1044 6102 1062 6120
rect 1044 6120 1062 6138
rect 1044 6138 1062 6156
rect 1044 6156 1062 6174
rect 1044 6174 1062 6192
rect 1062 1062 1080 1080
rect 1062 1080 1080 1098
rect 1062 1098 1080 1116
rect 1062 1116 1080 1134
rect 1062 1134 1080 1152
rect 1062 1152 1080 1170
rect 1062 1170 1080 1188
rect 1062 1188 1080 1206
rect 1062 1206 1080 1224
rect 1062 1224 1080 1242
rect 1062 1242 1080 1260
rect 1062 1260 1080 1278
rect 1062 1278 1080 1296
rect 1062 1296 1080 1314
rect 1062 1314 1080 1332
rect 1062 1332 1080 1350
rect 1062 1350 1080 1368
rect 1062 1368 1080 1386
rect 1062 1386 1080 1404
rect 1062 1404 1080 1422
rect 1062 1422 1080 1440
rect 1062 1440 1080 1458
rect 1062 1458 1080 1476
rect 1062 1476 1080 1494
rect 1062 1494 1080 1512
rect 1062 1512 1080 1530
rect 1062 1530 1080 1548
rect 1062 1548 1080 1566
rect 1062 1566 1080 1584
rect 1062 1584 1080 1602
rect 1062 1602 1080 1620
rect 1062 1620 1080 1638
rect 1062 1638 1080 1656
rect 1062 1656 1080 1674
rect 1062 1674 1080 1692
rect 1062 1692 1080 1710
rect 1062 1710 1080 1728
rect 1062 1728 1080 1746
rect 1062 1746 1080 1764
rect 1062 1764 1080 1782
rect 1062 1782 1080 1800
rect 1062 1800 1080 1818
rect 1062 1818 1080 1836
rect 1062 1836 1080 1854
rect 1062 1854 1080 1872
rect 1062 1872 1080 1890
rect 1062 1890 1080 1908
rect 1062 1908 1080 1926
rect 1062 1926 1080 1944
rect 1062 1944 1080 1962
rect 1062 1962 1080 1980
rect 1062 1980 1080 1998
rect 1062 1998 1080 2016
rect 1062 2016 1080 2034
rect 1062 2034 1080 2052
rect 1062 2052 1080 2070
rect 1062 5202 1080 5220
rect 1062 5220 1080 5238
rect 1062 5238 1080 5256
rect 1062 5256 1080 5274
rect 1062 5274 1080 5292
rect 1062 5292 1080 5310
rect 1062 5310 1080 5328
rect 1062 5328 1080 5346
rect 1062 5346 1080 5364
rect 1062 5364 1080 5382
rect 1062 5382 1080 5400
rect 1062 5400 1080 5418
rect 1062 5418 1080 5436
rect 1062 5436 1080 5454
rect 1062 5454 1080 5472
rect 1062 5472 1080 5490
rect 1062 5490 1080 5508
rect 1062 5508 1080 5526
rect 1062 5526 1080 5544
rect 1062 5544 1080 5562
rect 1062 5562 1080 5580
rect 1062 5580 1080 5598
rect 1062 5598 1080 5616
rect 1062 5616 1080 5634
rect 1062 5634 1080 5652
rect 1062 5652 1080 5670
rect 1062 5670 1080 5688
rect 1062 5688 1080 5706
rect 1062 5706 1080 5724
rect 1062 5724 1080 5742
rect 1062 5742 1080 5760
rect 1062 5760 1080 5778
rect 1062 5778 1080 5796
rect 1062 5796 1080 5814
rect 1062 5814 1080 5832
rect 1062 5832 1080 5850
rect 1062 5850 1080 5868
rect 1062 5868 1080 5886
rect 1062 5886 1080 5904
rect 1062 5904 1080 5922
rect 1062 5922 1080 5940
rect 1062 5940 1080 5958
rect 1062 5958 1080 5976
rect 1062 5976 1080 5994
rect 1062 5994 1080 6012
rect 1062 6012 1080 6030
rect 1062 6030 1080 6048
rect 1062 6048 1080 6066
rect 1062 6066 1080 6084
rect 1062 6084 1080 6102
rect 1062 6102 1080 6120
rect 1062 6120 1080 6138
rect 1062 6138 1080 6156
rect 1062 6156 1080 6174
rect 1062 6174 1080 6192
rect 1062 6192 1080 6210
rect 1080 1044 1098 1062
rect 1080 1062 1098 1080
rect 1080 1080 1098 1098
rect 1080 1098 1098 1116
rect 1080 1116 1098 1134
rect 1080 1134 1098 1152
rect 1080 1152 1098 1170
rect 1080 1170 1098 1188
rect 1080 1188 1098 1206
rect 1080 1206 1098 1224
rect 1080 1224 1098 1242
rect 1080 1242 1098 1260
rect 1080 1260 1098 1278
rect 1080 1278 1098 1296
rect 1080 1296 1098 1314
rect 1080 1314 1098 1332
rect 1080 1332 1098 1350
rect 1080 1350 1098 1368
rect 1080 1368 1098 1386
rect 1080 1386 1098 1404
rect 1080 1404 1098 1422
rect 1080 1422 1098 1440
rect 1080 1440 1098 1458
rect 1080 1458 1098 1476
rect 1080 1476 1098 1494
rect 1080 1494 1098 1512
rect 1080 1512 1098 1530
rect 1080 1530 1098 1548
rect 1080 1548 1098 1566
rect 1080 1566 1098 1584
rect 1080 1584 1098 1602
rect 1080 1602 1098 1620
rect 1080 1620 1098 1638
rect 1080 1638 1098 1656
rect 1080 1656 1098 1674
rect 1080 1674 1098 1692
rect 1080 1692 1098 1710
rect 1080 1710 1098 1728
rect 1080 1728 1098 1746
rect 1080 1746 1098 1764
rect 1080 1764 1098 1782
rect 1080 1782 1098 1800
rect 1080 1800 1098 1818
rect 1080 1818 1098 1836
rect 1080 1836 1098 1854
rect 1080 1854 1098 1872
rect 1080 1872 1098 1890
rect 1080 1890 1098 1908
rect 1080 1908 1098 1926
rect 1080 1926 1098 1944
rect 1080 1944 1098 1962
rect 1080 1962 1098 1980
rect 1080 1980 1098 1998
rect 1080 1998 1098 2016
rect 1080 2016 1098 2034
rect 1080 5238 1098 5256
rect 1080 5256 1098 5274
rect 1080 5274 1098 5292
rect 1080 5292 1098 5310
rect 1080 5310 1098 5328
rect 1080 5328 1098 5346
rect 1080 5346 1098 5364
rect 1080 5364 1098 5382
rect 1080 5382 1098 5400
rect 1080 5400 1098 5418
rect 1080 5418 1098 5436
rect 1080 5436 1098 5454
rect 1080 5454 1098 5472
rect 1080 5472 1098 5490
rect 1080 5490 1098 5508
rect 1080 5508 1098 5526
rect 1080 5526 1098 5544
rect 1080 5544 1098 5562
rect 1080 5562 1098 5580
rect 1080 5580 1098 5598
rect 1080 5598 1098 5616
rect 1080 5616 1098 5634
rect 1080 5634 1098 5652
rect 1080 5652 1098 5670
rect 1080 5670 1098 5688
rect 1080 5688 1098 5706
rect 1080 5706 1098 5724
rect 1080 5724 1098 5742
rect 1080 5742 1098 5760
rect 1080 5760 1098 5778
rect 1080 5778 1098 5796
rect 1080 5796 1098 5814
rect 1080 5814 1098 5832
rect 1080 5832 1098 5850
rect 1080 5850 1098 5868
rect 1080 5868 1098 5886
rect 1080 5886 1098 5904
rect 1080 5904 1098 5922
rect 1080 5922 1098 5940
rect 1080 5940 1098 5958
rect 1080 5958 1098 5976
rect 1080 5976 1098 5994
rect 1080 5994 1098 6012
rect 1080 6012 1098 6030
rect 1080 6030 1098 6048
rect 1080 6048 1098 6066
rect 1080 6066 1098 6084
rect 1080 6084 1098 6102
rect 1080 6102 1098 6120
rect 1080 6120 1098 6138
rect 1080 6138 1098 6156
rect 1080 6156 1098 6174
rect 1080 6174 1098 6192
rect 1080 6192 1098 6210
rect 1080 6210 1098 6228
rect 1098 1026 1116 1044
rect 1098 1044 1116 1062
rect 1098 1062 1116 1080
rect 1098 1080 1116 1098
rect 1098 1098 1116 1116
rect 1098 1116 1116 1134
rect 1098 1134 1116 1152
rect 1098 1152 1116 1170
rect 1098 1170 1116 1188
rect 1098 1188 1116 1206
rect 1098 1206 1116 1224
rect 1098 1224 1116 1242
rect 1098 1242 1116 1260
rect 1098 1260 1116 1278
rect 1098 1278 1116 1296
rect 1098 1296 1116 1314
rect 1098 1314 1116 1332
rect 1098 1332 1116 1350
rect 1098 1350 1116 1368
rect 1098 1368 1116 1386
rect 1098 1386 1116 1404
rect 1098 1404 1116 1422
rect 1098 1422 1116 1440
rect 1098 1440 1116 1458
rect 1098 1458 1116 1476
rect 1098 1476 1116 1494
rect 1098 1494 1116 1512
rect 1098 1512 1116 1530
rect 1098 1530 1116 1548
rect 1098 1548 1116 1566
rect 1098 1566 1116 1584
rect 1098 1584 1116 1602
rect 1098 1602 1116 1620
rect 1098 1620 1116 1638
rect 1098 1638 1116 1656
rect 1098 1656 1116 1674
rect 1098 1674 1116 1692
rect 1098 1692 1116 1710
rect 1098 1710 1116 1728
rect 1098 1728 1116 1746
rect 1098 1746 1116 1764
rect 1098 1764 1116 1782
rect 1098 1782 1116 1800
rect 1098 1800 1116 1818
rect 1098 1818 1116 1836
rect 1098 1836 1116 1854
rect 1098 1854 1116 1872
rect 1098 1872 1116 1890
rect 1098 1890 1116 1908
rect 1098 1908 1116 1926
rect 1098 1926 1116 1944
rect 1098 1944 1116 1962
rect 1098 1962 1116 1980
rect 1098 1980 1116 1998
rect 1098 1998 1116 2016
rect 1098 5256 1116 5274
rect 1098 5274 1116 5292
rect 1098 5292 1116 5310
rect 1098 5310 1116 5328
rect 1098 5328 1116 5346
rect 1098 5346 1116 5364
rect 1098 5364 1116 5382
rect 1098 5382 1116 5400
rect 1098 5400 1116 5418
rect 1098 5418 1116 5436
rect 1098 5436 1116 5454
rect 1098 5454 1116 5472
rect 1098 5472 1116 5490
rect 1098 5490 1116 5508
rect 1098 5508 1116 5526
rect 1098 5526 1116 5544
rect 1098 5544 1116 5562
rect 1098 5562 1116 5580
rect 1098 5580 1116 5598
rect 1098 5598 1116 5616
rect 1098 5616 1116 5634
rect 1098 5634 1116 5652
rect 1098 5652 1116 5670
rect 1098 5670 1116 5688
rect 1098 5688 1116 5706
rect 1098 5706 1116 5724
rect 1098 5724 1116 5742
rect 1098 5742 1116 5760
rect 1098 5760 1116 5778
rect 1098 5778 1116 5796
rect 1098 5796 1116 5814
rect 1098 5814 1116 5832
rect 1098 5832 1116 5850
rect 1098 5850 1116 5868
rect 1098 5868 1116 5886
rect 1098 5886 1116 5904
rect 1098 5904 1116 5922
rect 1098 5922 1116 5940
rect 1098 5940 1116 5958
rect 1098 5958 1116 5976
rect 1098 5976 1116 5994
rect 1098 5994 1116 6012
rect 1098 6012 1116 6030
rect 1098 6030 1116 6048
rect 1098 6048 1116 6066
rect 1098 6066 1116 6084
rect 1098 6084 1116 6102
rect 1098 6102 1116 6120
rect 1098 6120 1116 6138
rect 1098 6138 1116 6156
rect 1098 6156 1116 6174
rect 1098 6174 1116 6192
rect 1098 6192 1116 6210
rect 1098 6210 1116 6228
rect 1098 6228 1116 6246
rect 1116 1008 1134 1026
rect 1116 1026 1134 1044
rect 1116 1044 1134 1062
rect 1116 1062 1134 1080
rect 1116 1080 1134 1098
rect 1116 1098 1134 1116
rect 1116 1116 1134 1134
rect 1116 1134 1134 1152
rect 1116 1152 1134 1170
rect 1116 1170 1134 1188
rect 1116 1188 1134 1206
rect 1116 1206 1134 1224
rect 1116 1224 1134 1242
rect 1116 1242 1134 1260
rect 1116 1260 1134 1278
rect 1116 1278 1134 1296
rect 1116 1296 1134 1314
rect 1116 1314 1134 1332
rect 1116 1332 1134 1350
rect 1116 1350 1134 1368
rect 1116 1368 1134 1386
rect 1116 1386 1134 1404
rect 1116 1404 1134 1422
rect 1116 1422 1134 1440
rect 1116 1440 1134 1458
rect 1116 1458 1134 1476
rect 1116 1476 1134 1494
rect 1116 1494 1134 1512
rect 1116 1512 1134 1530
rect 1116 1530 1134 1548
rect 1116 1548 1134 1566
rect 1116 1566 1134 1584
rect 1116 1584 1134 1602
rect 1116 1602 1134 1620
rect 1116 1620 1134 1638
rect 1116 1638 1134 1656
rect 1116 1656 1134 1674
rect 1116 1674 1134 1692
rect 1116 1692 1134 1710
rect 1116 1710 1134 1728
rect 1116 1728 1134 1746
rect 1116 1746 1134 1764
rect 1116 1764 1134 1782
rect 1116 1782 1134 1800
rect 1116 1800 1134 1818
rect 1116 1818 1134 1836
rect 1116 1836 1134 1854
rect 1116 1854 1134 1872
rect 1116 1872 1134 1890
rect 1116 1890 1134 1908
rect 1116 1908 1134 1926
rect 1116 1926 1134 1944
rect 1116 1944 1134 1962
rect 1116 1962 1134 1980
rect 1116 5292 1134 5310
rect 1116 5310 1134 5328
rect 1116 5328 1134 5346
rect 1116 5346 1134 5364
rect 1116 5364 1134 5382
rect 1116 5382 1134 5400
rect 1116 5400 1134 5418
rect 1116 5418 1134 5436
rect 1116 5436 1134 5454
rect 1116 5454 1134 5472
rect 1116 5472 1134 5490
rect 1116 5490 1134 5508
rect 1116 5508 1134 5526
rect 1116 5526 1134 5544
rect 1116 5544 1134 5562
rect 1116 5562 1134 5580
rect 1116 5580 1134 5598
rect 1116 5598 1134 5616
rect 1116 5616 1134 5634
rect 1116 5634 1134 5652
rect 1116 5652 1134 5670
rect 1116 5670 1134 5688
rect 1116 5688 1134 5706
rect 1116 5706 1134 5724
rect 1116 5724 1134 5742
rect 1116 5742 1134 5760
rect 1116 5760 1134 5778
rect 1116 5778 1134 5796
rect 1116 5796 1134 5814
rect 1116 5814 1134 5832
rect 1116 5832 1134 5850
rect 1116 5850 1134 5868
rect 1116 5868 1134 5886
rect 1116 5886 1134 5904
rect 1116 5904 1134 5922
rect 1116 5922 1134 5940
rect 1116 5940 1134 5958
rect 1116 5958 1134 5976
rect 1116 5976 1134 5994
rect 1116 5994 1134 6012
rect 1116 6012 1134 6030
rect 1116 6030 1134 6048
rect 1116 6048 1134 6066
rect 1116 6066 1134 6084
rect 1116 6084 1134 6102
rect 1116 6102 1134 6120
rect 1116 6120 1134 6138
rect 1116 6138 1134 6156
rect 1116 6156 1134 6174
rect 1116 6174 1134 6192
rect 1116 6192 1134 6210
rect 1116 6210 1134 6228
rect 1116 6228 1134 6246
rect 1116 6246 1134 6264
rect 1134 990 1152 1008
rect 1134 1008 1152 1026
rect 1134 1026 1152 1044
rect 1134 1044 1152 1062
rect 1134 1062 1152 1080
rect 1134 1080 1152 1098
rect 1134 1098 1152 1116
rect 1134 1116 1152 1134
rect 1134 1134 1152 1152
rect 1134 1152 1152 1170
rect 1134 1170 1152 1188
rect 1134 1188 1152 1206
rect 1134 1206 1152 1224
rect 1134 1224 1152 1242
rect 1134 1242 1152 1260
rect 1134 1260 1152 1278
rect 1134 1278 1152 1296
rect 1134 1296 1152 1314
rect 1134 1314 1152 1332
rect 1134 1332 1152 1350
rect 1134 1350 1152 1368
rect 1134 1368 1152 1386
rect 1134 1386 1152 1404
rect 1134 1404 1152 1422
rect 1134 1422 1152 1440
rect 1134 1440 1152 1458
rect 1134 1458 1152 1476
rect 1134 1476 1152 1494
rect 1134 1494 1152 1512
rect 1134 1512 1152 1530
rect 1134 1530 1152 1548
rect 1134 1548 1152 1566
rect 1134 1566 1152 1584
rect 1134 1584 1152 1602
rect 1134 1602 1152 1620
rect 1134 1620 1152 1638
rect 1134 1638 1152 1656
rect 1134 1656 1152 1674
rect 1134 1674 1152 1692
rect 1134 1692 1152 1710
rect 1134 1710 1152 1728
rect 1134 1728 1152 1746
rect 1134 1746 1152 1764
rect 1134 1764 1152 1782
rect 1134 1782 1152 1800
rect 1134 1800 1152 1818
rect 1134 1818 1152 1836
rect 1134 1836 1152 1854
rect 1134 1854 1152 1872
rect 1134 1872 1152 1890
rect 1134 1890 1152 1908
rect 1134 1908 1152 1926
rect 1134 1926 1152 1944
rect 1134 5310 1152 5328
rect 1134 5328 1152 5346
rect 1134 5346 1152 5364
rect 1134 5364 1152 5382
rect 1134 5382 1152 5400
rect 1134 5400 1152 5418
rect 1134 5418 1152 5436
rect 1134 5436 1152 5454
rect 1134 5454 1152 5472
rect 1134 5472 1152 5490
rect 1134 5490 1152 5508
rect 1134 5508 1152 5526
rect 1134 5526 1152 5544
rect 1134 5544 1152 5562
rect 1134 5562 1152 5580
rect 1134 5580 1152 5598
rect 1134 5598 1152 5616
rect 1134 5616 1152 5634
rect 1134 5634 1152 5652
rect 1134 5652 1152 5670
rect 1134 5670 1152 5688
rect 1134 5688 1152 5706
rect 1134 5706 1152 5724
rect 1134 5724 1152 5742
rect 1134 5742 1152 5760
rect 1134 5760 1152 5778
rect 1134 5778 1152 5796
rect 1134 5796 1152 5814
rect 1134 5814 1152 5832
rect 1134 5832 1152 5850
rect 1134 5850 1152 5868
rect 1134 5868 1152 5886
rect 1134 5886 1152 5904
rect 1134 5904 1152 5922
rect 1134 5922 1152 5940
rect 1134 5940 1152 5958
rect 1134 5958 1152 5976
rect 1134 5976 1152 5994
rect 1134 5994 1152 6012
rect 1134 6012 1152 6030
rect 1134 6030 1152 6048
rect 1134 6048 1152 6066
rect 1134 6066 1152 6084
rect 1134 6084 1152 6102
rect 1134 6102 1152 6120
rect 1134 6120 1152 6138
rect 1134 6138 1152 6156
rect 1134 6156 1152 6174
rect 1134 6174 1152 6192
rect 1134 6192 1152 6210
rect 1134 6210 1152 6228
rect 1134 6228 1152 6246
rect 1134 6246 1152 6264
rect 1134 6264 1152 6282
rect 1152 972 1170 990
rect 1152 990 1170 1008
rect 1152 1008 1170 1026
rect 1152 1026 1170 1044
rect 1152 1044 1170 1062
rect 1152 1062 1170 1080
rect 1152 1080 1170 1098
rect 1152 1098 1170 1116
rect 1152 1116 1170 1134
rect 1152 1134 1170 1152
rect 1152 1152 1170 1170
rect 1152 1170 1170 1188
rect 1152 1188 1170 1206
rect 1152 1206 1170 1224
rect 1152 1224 1170 1242
rect 1152 1242 1170 1260
rect 1152 1260 1170 1278
rect 1152 1278 1170 1296
rect 1152 1296 1170 1314
rect 1152 1314 1170 1332
rect 1152 1332 1170 1350
rect 1152 1350 1170 1368
rect 1152 1368 1170 1386
rect 1152 1386 1170 1404
rect 1152 1404 1170 1422
rect 1152 1422 1170 1440
rect 1152 1440 1170 1458
rect 1152 1458 1170 1476
rect 1152 1476 1170 1494
rect 1152 1494 1170 1512
rect 1152 1512 1170 1530
rect 1152 1530 1170 1548
rect 1152 1548 1170 1566
rect 1152 1566 1170 1584
rect 1152 1584 1170 1602
rect 1152 1602 1170 1620
rect 1152 1620 1170 1638
rect 1152 1638 1170 1656
rect 1152 1656 1170 1674
rect 1152 1674 1170 1692
rect 1152 1692 1170 1710
rect 1152 1710 1170 1728
rect 1152 1728 1170 1746
rect 1152 1746 1170 1764
rect 1152 1764 1170 1782
rect 1152 1782 1170 1800
rect 1152 1800 1170 1818
rect 1152 1818 1170 1836
rect 1152 1836 1170 1854
rect 1152 1854 1170 1872
rect 1152 1872 1170 1890
rect 1152 1890 1170 1908
rect 1152 1908 1170 1926
rect 1152 5346 1170 5364
rect 1152 5364 1170 5382
rect 1152 5382 1170 5400
rect 1152 5400 1170 5418
rect 1152 5418 1170 5436
rect 1152 5436 1170 5454
rect 1152 5454 1170 5472
rect 1152 5472 1170 5490
rect 1152 5490 1170 5508
rect 1152 5508 1170 5526
rect 1152 5526 1170 5544
rect 1152 5544 1170 5562
rect 1152 5562 1170 5580
rect 1152 5580 1170 5598
rect 1152 5598 1170 5616
rect 1152 5616 1170 5634
rect 1152 5634 1170 5652
rect 1152 5652 1170 5670
rect 1152 5670 1170 5688
rect 1152 5688 1170 5706
rect 1152 5706 1170 5724
rect 1152 5724 1170 5742
rect 1152 5742 1170 5760
rect 1152 5760 1170 5778
rect 1152 5778 1170 5796
rect 1152 5796 1170 5814
rect 1152 5814 1170 5832
rect 1152 5832 1170 5850
rect 1152 5850 1170 5868
rect 1152 5868 1170 5886
rect 1152 5886 1170 5904
rect 1152 5904 1170 5922
rect 1152 5922 1170 5940
rect 1152 5940 1170 5958
rect 1152 5958 1170 5976
rect 1152 5976 1170 5994
rect 1152 5994 1170 6012
rect 1152 6012 1170 6030
rect 1152 6030 1170 6048
rect 1152 6048 1170 6066
rect 1152 6066 1170 6084
rect 1152 6084 1170 6102
rect 1152 6102 1170 6120
rect 1152 6120 1170 6138
rect 1152 6138 1170 6156
rect 1152 6156 1170 6174
rect 1152 6174 1170 6192
rect 1152 6192 1170 6210
rect 1152 6210 1170 6228
rect 1152 6228 1170 6246
rect 1152 6246 1170 6264
rect 1152 6264 1170 6282
rect 1152 6282 1170 6300
rect 1170 954 1188 972
rect 1170 972 1188 990
rect 1170 990 1188 1008
rect 1170 1008 1188 1026
rect 1170 1026 1188 1044
rect 1170 1044 1188 1062
rect 1170 1062 1188 1080
rect 1170 1080 1188 1098
rect 1170 1098 1188 1116
rect 1170 1116 1188 1134
rect 1170 1134 1188 1152
rect 1170 1152 1188 1170
rect 1170 1170 1188 1188
rect 1170 1188 1188 1206
rect 1170 1206 1188 1224
rect 1170 1224 1188 1242
rect 1170 1242 1188 1260
rect 1170 1260 1188 1278
rect 1170 1278 1188 1296
rect 1170 1296 1188 1314
rect 1170 1314 1188 1332
rect 1170 1332 1188 1350
rect 1170 1350 1188 1368
rect 1170 1368 1188 1386
rect 1170 1386 1188 1404
rect 1170 1404 1188 1422
rect 1170 1422 1188 1440
rect 1170 1440 1188 1458
rect 1170 1458 1188 1476
rect 1170 1476 1188 1494
rect 1170 1494 1188 1512
rect 1170 1512 1188 1530
rect 1170 1530 1188 1548
rect 1170 1548 1188 1566
rect 1170 1566 1188 1584
rect 1170 1584 1188 1602
rect 1170 1602 1188 1620
rect 1170 1620 1188 1638
rect 1170 1638 1188 1656
rect 1170 1656 1188 1674
rect 1170 1674 1188 1692
rect 1170 1692 1188 1710
rect 1170 1710 1188 1728
rect 1170 1728 1188 1746
rect 1170 1746 1188 1764
rect 1170 1764 1188 1782
rect 1170 1782 1188 1800
rect 1170 1800 1188 1818
rect 1170 1818 1188 1836
rect 1170 1836 1188 1854
rect 1170 1854 1188 1872
rect 1170 1872 1188 1890
rect 1170 1890 1188 1908
rect 1170 5364 1188 5382
rect 1170 5382 1188 5400
rect 1170 5400 1188 5418
rect 1170 5418 1188 5436
rect 1170 5436 1188 5454
rect 1170 5454 1188 5472
rect 1170 5472 1188 5490
rect 1170 5490 1188 5508
rect 1170 5508 1188 5526
rect 1170 5526 1188 5544
rect 1170 5544 1188 5562
rect 1170 5562 1188 5580
rect 1170 5580 1188 5598
rect 1170 5598 1188 5616
rect 1170 5616 1188 5634
rect 1170 5634 1188 5652
rect 1170 5652 1188 5670
rect 1170 5670 1188 5688
rect 1170 5688 1188 5706
rect 1170 5706 1188 5724
rect 1170 5724 1188 5742
rect 1170 5742 1188 5760
rect 1170 5760 1188 5778
rect 1170 5778 1188 5796
rect 1170 5796 1188 5814
rect 1170 5814 1188 5832
rect 1170 5832 1188 5850
rect 1170 5850 1188 5868
rect 1170 5868 1188 5886
rect 1170 5886 1188 5904
rect 1170 5904 1188 5922
rect 1170 5922 1188 5940
rect 1170 5940 1188 5958
rect 1170 5958 1188 5976
rect 1170 5976 1188 5994
rect 1170 5994 1188 6012
rect 1170 6012 1188 6030
rect 1170 6030 1188 6048
rect 1170 6048 1188 6066
rect 1170 6066 1188 6084
rect 1170 6084 1188 6102
rect 1170 6102 1188 6120
rect 1170 6120 1188 6138
rect 1170 6138 1188 6156
rect 1170 6156 1188 6174
rect 1170 6174 1188 6192
rect 1170 6192 1188 6210
rect 1170 6210 1188 6228
rect 1170 6228 1188 6246
rect 1170 6246 1188 6264
rect 1170 6264 1188 6282
rect 1170 6282 1188 6300
rect 1170 6300 1188 6318
rect 1188 936 1206 954
rect 1188 954 1206 972
rect 1188 972 1206 990
rect 1188 990 1206 1008
rect 1188 1008 1206 1026
rect 1188 1026 1206 1044
rect 1188 1044 1206 1062
rect 1188 1062 1206 1080
rect 1188 1080 1206 1098
rect 1188 1098 1206 1116
rect 1188 1116 1206 1134
rect 1188 1134 1206 1152
rect 1188 1152 1206 1170
rect 1188 1170 1206 1188
rect 1188 1188 1206 1206
rect 1188 1206 1206 1224
rect 1188 1224 1206 1242
rect 1188 1242 1206 1260
rect 1188 1260 1206 1278
rect 1188 1278 1206 1296
rect 1188 1296 1206 1314
rect 1188 1314 1206 1332
rect 1188 1332 1206 1350
rect 1188 1350 1206 1368
rect 1188 1368 1206 1386
rect 1188 1386 1206 1404
rect 1188 1404 1206 1422
rect 1188 1422 1206 1440
rect 1188 1440 1206 1458
rect 1188 1458 1206 1476
rect 1188 1476 1206 1494
rect 1188 1494 1206 1512
rect 1188 1512 1206 1530
rect 1188 1530 1206 1548
rect 1188 1548 1206 1566
rect 1188 1566 1206 1584
rect 1188 1584 1206 1602
rect 1188 1602 1206 1620
rect 1188 1620 1206 1638
rect 1188 1638 1206 1656
rect 1188 1656 1206 1674
rect 1188 1674 1206 1692
rect 1188 1692 1206 1710
rect 1188 1710 1206 1728
rect 1188 1728 1206 1746
rect 1188 1746 1206 1764
rect 1188 1764 1206 1782
rect 1188 1782 1206 1800
rect 1188 1800 1206 1818
rect 1188 1818 1206 1836
rect 1188 1836 1206 1854
rect 1188 1854 1206 1872
rect 1188 5400 1206 5418
rect 1188 5418 1206 5436
rect 1188 5436 1206 5454
rect 1188 5454 1206 5472
rect 1188 5472 1206 5490
rect 1188 5490 1206 5508
rect 1188 5508 1206 5526
rect 1188 5526 1206 5544
rect 1188 5544 1206 5562
rect 1188 5562 1206 5580
rect 1188 5580 1206 5598
rect 1188 5598 1206 5616
rect 1188 5616 1206 5634
rect 1188 5634 1206 5652
rect 1188 5652 1206 5670
rect 1188 5670 1206 5688
rect 1188 5688 1206 5706
rect 1188 5706 1206 5724
rect 1188 5724 1206 5742
rect 1188 5742 1206 5760
rect 1188 5760 1206 5778
rect 1188 5778 1206 5796
rect 1188 5796 1206 5814
rect 1188 5814 1206 5832
rect 1188 5832 1206 5850
rect 1188 5850 1206 5868
rect 1188 5868 1206 5886
rect 1188 5886 1206 5904
rect 1188 5904 1206 5922
rect 1188 5922 1206 5940
rect 1188 5940 1206 5958
rect 1188 5958 1206 5976
rect 1188 5976 1206 5994
rect 1188 5994 1206 6012
rect 1188 6012 1206 6030
rect 1188 6030 1206 6048
rect 1188 6048 1206 6066
rect 1188 6066 1206 6084
rect 1188 6084 1206 6102
rect 1188 6102 1206 6120
rect 1188 6120 1206 6138
rect 1188 6138 1206 6156
rect 1188 6156 1206 6174
rect 1188 6174 1206 6192
rect 1188 6192 1206 6210
rect 1188 6210 1206 6228
rect 1188 6228 1206 6246
rect 1188 6246 1206 6264
rect 1188 6264 1206 6282
rect 1188 6282 1206 6300
rect 1188 6300 1206 6318
rect 1188 6318 1206 6336
rect 1206 918 1224 936
rect 1206 936 1224 954
rect 1206 954 1224 972
rect 1206 972 1224 990
rect 1206 990 1224 1008
rect 1206 1008 1224 1026
rect 1206 1026 1224 1044
rect 1206 1044 1224 1062
rect 1206 1062 1224 1080
rect 1206 1080 1224 1098
rect 1206 1098 1224 1116
rect 1206 1116 1224 1134
rect 1206 1134 1224 1152
rect 1206 1152 1224 1170
rect 1206 1170 1224 1188
rect 1206 1188 1224 1206
rect 1206 1206 1224 1224
rect 1206 1224 1224 1242
rect 1206 1242 1224 1260
rect 1206 1260 1224 1278
rect 1206 1278 1224 1296
rect 1206 1296 1224 1314
rect 1206 1314 1224 1332
rect 1206 1332 1224 1350
rect 1206 1350 1224 1368
rect 1206 1368 1224 1386
rect 1206 1386 1224 1404
rect 1206 1404 1224 1422
rect 1206 1422 1224 1440
rect 1206 1440 1224 1458
rect 1206 1458 1224 1476
rect 1206 1476 1224 1494
rect 1206 1494 1224 1512
rect 1206 1512 1224 1530
rect 1206 1530 1224 1548
rect 1206 1548 1224 1566
rect 1206 1566 1224 1584
rect 1206 1584 1224 1602
rect 1206 1602 1224 1620
rect 1206 1620 1224 1638
rect 1206 1638 1224 1656
rect 1206 1656 1224 1674
rect 1206 1674 1224 1692
rect 1206 1692 1224 1710
rect 1206 1710 1224 1728
rect 1206 1728 1224 1746
rect 1206 1746 1224 1764
rect 1206 1764 1224 1782
rect 1206 1782 1224 1800
rect 1206 1800 1224 1818
rect 1206 1818 1224 1836
rect 1206 1836 1224 1854
rect 1206 5418 1224 5436
rect 1206 5436 1224 5454
rect 1206 5454 1224 5472
rect 1206 5472 1224 5490
rect 1206 5490 1224 5508
rect 1206 5508 1224 5526
rect 1206 5526 1224 5544
rect 1206 5544 1224 5562
rect 1206 5562 1224 5580
rect 1206 5580 1224 5598
rect 1206 5598 1224 5616
rect 1206 5616 1224 5634
rect 1206 5634 1224 5652
rect 1206 5652 1224 5670
rect 1206 5670 1224 5688
rect 1206 5688 1224 5706
rect 1206 5706 1224 5724
rect 1206 5724 1224 5742
rect 1206 5742 1224 5760
rect 1206 5760 1224 5778
rect 1206 5778 1224 5796
rect 1206 5796 1224 5814
rect 1206 5814 1224 5832
rect 1206 5832 1224 5850
rect 1206 5850 1224 5868
rect 1206 5868 1224 5886
rect 1206 5886 1224 5904
rect 1206 5904 1224 5922
rect 1206 5922 1224 5940
rect 1206 5940 1224 5958
rect 1206 5958 1224 5976
rect 1206 5976 1224 5994
rect 1206 5994 1224 6012
rect 1206 6012 1224 6030
rect 1206 6030 1224 6048
rect 1206 6048 1224 6066
rect 1206 6066 1224 6084
rect 1206 6084 1224 6102
rect 1206 6102 1224 6120
rect 1206 6120 1224 6138
rect 1206 6138 1224 6156
rect 1206 6156 1224 6174
rect 1206 6174 1224 6192
rect 1206 6192 1224 6210
rect 1206 6210 1224 6228
rect 1206 6228 1224 6246
rect 1206 6246 1224 6264
rect 1206 6264 1224 6282
rect 1206 6282 1224 6300
rect 1206 6300 1224 6318
rect 1206 6318 1224 6336
rect 1206 6336 1224 6354
rect 1224 900 1242 918
rect 1224 918 1242 936
rect 1224 936 1242 954
rect 1224 954 1242 972
rect 1224 972 1242 990
rect 1224 990 1242 1008
rect 1224 1008 1242 1026
rect 1224 1026 1242 1044
rect 1224 1044 1242 1062
rect 1224 1062 1242 1080
rect 1224 1080 1242 1098
rect 1224 1098 1242 1116
rect 1224 1116 1242 1134
rect 1224 1134 1242 1152
rect 1224 1152 1242 1170
rect 1224 1170 1242 1188
rect 1224 1188 1242 1206
rect 1224 1206 1242 1224
rect 1224 1224 1242 1242
rect 1224 1242 1242 1260
rect 1224 1260 1242 1278
rect 1224 1278 1242 1296
rect 1224 1296 1242 1314
rect 1224 1314 1242 1332
rect 1224 1332 1242 1350
rect 1224 1350 1242 1368
rect 1224 1368 1242 1386
rect 1224 1386 1242 1404
rect 1224 1404 1242 1422
rect 1224 1422 1242 1440
rect 1224 1440 1242 1458
rect 1224 1458 1242 1476
rect 1224 1476 1242 1494
rect 1224 1494 1242 1512
rect 1224 1512 1242 1530
rect 1224 1530 1242 1548
rect 1224 1548 1242 1566
rect 1224 1566 1242 1584
rect 1224 1584 1242 1602
rect 1224 1602 1242 1620
rect 1224 1620 1242 1638
rect 1224 1638 1242 1656
rect 1224 1656 1242 1674
rect 1224 1674 1242 1692
rect 1224 1692 1242 1710
rect 1224 1710 1242 1728
rect 1224 1728 1242 1746
rect 1224 1746 1242 1764
rect 1224 1764 1242 1782
rect 1224 1782 1242 1800
rect 1224 1800 1242 1818
rect 1224 5436 1242 5454
rect 1224 5454 1242 5472
rect 1224 5472 1242 5490
rect 1224 5490 1242 5508
rect 1224 5508 1242 5526
rect 1224 5526 1242 5544
rect 1224 5544 1242 5562
rect 1224 5562 1242 5580
rect 1224 5580 1242 5598
rect 1224 5598 1242 5616
rect 1224 5616 1242 5634
rect 1224 5634 1242 5652
rect 1224 5652 1242 5670
rect 1224 5670 1242 5688
rect 1224 5688 1242 5706
rect 1224 5706 1242 5724
rect 1224 5724 1242 5742
rect 1224 5742 1242 5760
rect 1224 5760 1242 5778
rect 1224 5778 1242 5796
rect 1224 5796 1242 5814
rect 1224 5814 1242 5832
rect 1224 5832 1242 5850
rect 1224 5850 1242 5868
rect 1224 5868 1242 5886
rect 1224 5886 1242 5904
rect 1224 5904 1242 5922
rect 1224 5922 1242 5940
rect 1224 5940 1242 5958
rect 1224 5958 1242 5976
rect 1224 5976 1242 5994
rect 1224 5994 1242 6012
rect 1224 6012 1242 6030
rect 1224 6030 1242 6048
rect 1224 6048 1242 6066
rect 1224 6066 1242 6084
rect 1224 6084 1242 6102
rect 1224 6102 1242 6120
rect 1224 6120 1242 6138
rect 1224 6138 1242 6156
rect 1224 6156 1242 6174
rect 1224 6174 1242 6192
rect 1224 6192 1242 6210
rect 1224 6210 1242 6228
rect 1224 6228 1242 6246
rect 1224 6246 1242 6264
rect 1224 6264 1242 6282
rect 1224 6282 1242 6300
rect 1224 6300 1242 6318
rect 1224 6318 1242 6336
rect 1224 6336 1242 6354
rect 1242 900 1260 918
rect 1242 918 1260 936
rect 1242 936 1260 954
rect 1242 954 1260 972
rect 1242 972 1260 990
rect 1242 990 1260 1008
rect 1242 1008 1260 1026
rect 1242 1026 1260 1044
rect 1242 1044 1260 1062
rect 1242 1062 1260 1080
rect 1242 1080 1260 1098
rect 1242 1098 1260 1116
rect 1242 1116 1260 1134
rect 1242 1134 1260 1152
rect 1242 1152 1260 1170
rect 1242 1170 1260 1188
rect 1242 1188 1260 1206
rect 1242 1206 1260 1224
rect 1242 1224 1260 1242
rect 1242 1242 1260 1260
rect 1242 1260 1260 1278
rect 1242 1278 1260 1296
rect 1242 1296 1260 1314
rect 1242 1314 1260 1332
rect 1242 1332 1260 1350
rect 1242 1350 1260 1368
rect 1242 1368 1260 1386
rect 1242 1386 1260 1404
rect 1242 1404 1260 1422
rect 1242 1422 1260 1440
rect 1242 1440 1260 1458
rect 1242 1458 1260 1476
rect 1242 1476 1260 1494
rect 1242 1494 1260 1512
rect 1242 1512 1260 1530
rect 1242 1530 1260 1548
rect 1242 1548 1260 1566
rect 1242 1566 1260 1584
rect 1242 1584 1260 1602
rect 1242 1602 1260 1620
rect 1242 1620 1260 1638
rect 1242 1638 1260 1656
rect 1242 1656 1260 1674
rect 1242 1674 1260 1692
rect 1242 1692 1260 1710
rect 1242 1710 1260 1728
rect 1242 1728 1260 1746
rect 1242 1746 1260 1764
rect 1242 1764 1260 1782
rect 1242 1782 1260 1800
rect 1242 5472 1260 5490
rect 1242 5490 1260 5508
rect 1242 5508 1260 5526
rect 1242 5526 1260 5544
rect 1242 5544 1260 5562
rect 1242 5562 1260 5580
rect 1242 5580 1260 5598
rect 1242 5598 1260 5616
rect 1242 5616 1260 5634
rect 1242 5634 1260 5652
rect 1242 5652 1260 5670
rect 1242 5670 1260 5688
rect 1242 5688 1260 5706
rect 1242 5706 1260 5724
rect 1242 5724 1260 5742
rect 1242 5742 1260 5760
rect 1242 5760 1260 5778
rect 1242 5778 1260 5796
rect 1242 5796 1260 5814
rect 1242 5814 1260 5832
rect 1242 5832 1260 5850
rect 1242 5850 1260 5868
rect 1242 5868 1260 5886
rect 1242 5886 1260 5904
rect 1242 5904 1260 5922
rect 1242 5922 1260 5940
rect 1242 5940 1260 5958
rect 1242 5958 1260 5976
rect 1242 5976 1260 5994
rect 1242 5994 1260 6012
rect 1242 6012 1260 6030
rect 1242 6030 1260 6048
rect 1242 6048 1260 6066
rect 1242 6066 1260 6084
rect 1242 6084 1260 6102
rect 1242 6102 1260 6120
rect 1242 6120 1260 6138
rect 1242 6138 1260 6156
rect 1242 6156 1260 6174
rect 1242 6174 1260 6192
rect 1242 6192 1260 6210
rect 1242 6210 1260 6228
rect 1242 6228 1260 6246
rect 1242 6246 1260 6264
rect 1242 6264 1260 6282
rect 1242 6282 1260 6300
rect 1242 6300 1260 6318
rect 1242 6318 1260 6336
rect 1242 6336 1260 6354
rect 1242 6354 1260 6372
rect 1260 882 1278 900
rect 1260 900 1278 918
rect 1260 918 1278 936
rect 1260 936 1278 954
rect 1260 954 1278 972
rect 1260 972 1278 990
rect 1260 990 1278 1008
rect 1260 1008 1278 1026
rect 1260 1026 1278 1044
rect 1260 1044 1278 1062
rect 1260 1062 1278 1080
rect 1260 1080 1278 1098
rect 1260 1098 1278 1116
rect 1260 1116 1278 1134
rect 1260 1134 1278 1152
rect 1260 1152 1278 1170
rect 1260 1170 1278 1188
rect 1260 1188 1278 1206
rect 1260 1206 1278 1224
rect 1260 1224 1278 1242
rect 1260 1242 1278 1260
rect 1260 1260 1278 1278
rect 1260 1278 1278 1296
rect 1260 1296 1278 1314
rect 1260 1314 1278 1332
rect 1260 1332 1278 1350
rect 1260 1350 1278 1368
rect 1260 1368 1278 1386
rect 1260 1386 1278 1404
rect 1260 1404 1278 1422
rect 1260 1422 1278 1440
rect 1260 1440 1278 1458
rect 1260 1458 1278 1476
rect 1260 1476 1278 1494
rect 1260 1494 1278 1512
rect 1260 1512 1278 1530
rect 1260 1530 1278 1548
rect 1260 1548 1278 1566
rect 1260 1566 1278 1584
rect 1260 1584 1278 1602
rect 1260 1602 1278 1620
rect 1260 1620 1278 1638
rect 1260 1638 1278 1656
rect 1260 1656 1278 1674
rect 1260 1674 1278 1692
rect 1260 1692 1278 1710
rect 1260 1710 1278 1728
rect 1260 1728 1278 1746
rect 1260 1746 1278 1764
rect 1260 1764 1278 1782
rect 1260 5490 1278 5508
rect 1260 5508 1278 5526
rect 1260 5526 1278 5544
rect 1260 5544 1278 5562
rect 1260 5562 1278 5580
rect 1260 5580 1278 5598
rect 1260 5598 1278 5616
rect 1260 5616 1278 5634
rect 1260 5634 1278 5652
rect 1260 5652 1278 5670
rect 1260 5670 1278 5688
rect 1260 5688 1278 5706
rect 1260 5706 1278 5724
rect 1260 5724 1278 5742
rect 1260 5742 1278 5760
rect 1260 5760 1278 5778
rect 1260 5778 1278 5796
rect 1260 5796 1278 5814
rect 1260 5814 1278 5832
rect 1260 5832 1278 5850
rect 1260 5850 1278 5868
rect 1260 5868 1278 5886
rect 1260 5886 1278 5904
rect 1260 5904 1278 5922
rect 1260 5922 1278 5940
rect 1260 5940 1278 5958
rect 1260 5958 1278 5976
rect 1260 5976 1278 5994
rect 1260 5994 1278 6012
rect 1260 6012 1278 6030
rect 1260 6030 1278 6048
rect 1260 6048 1278 6066
rect 1260 6066 1278 6084
rect 1260 6084 1278 6102
rect 1260 6102 1278 6120
rect 1260 6120 1278 6138
rect 1260 6138 1278 6156
rect 1260 6156 1278 6174
rect 1260 6174 1278 6192
rect 1260 6192 1278 6210
rect 1260 6210 1278 6228
rect 1260 6228 1278 6246
rect 1260 6246 1278 6264
rect 1260 6264 1278 6282
rect 1260 6282 1278 6300
rect 1260 6300 1278 6318
rect 1260 6318 1278 6336
rect 1260 6336 1278 6354
rect 1260 6354 1278 6372
rect 1260 6372 1278 6390
rect 1278 864 1296 882
rect 1278 882 1296 900
rect 1278 900 1296 918
rect 1278 918 1296 936
rect 1278 936 1296 954
rect 1278 954 1296 972
rect 1278 972 1296 990
rect 1278 990 1296 1008
rect 1278 1008 1296 1026
rect 1278 1026 1296 1044
rect 1278 1044 1296 1062
rect 1278 1062 1296 1080
rect 1278 1080 1296 1098
rect 1278 1098 1296 1116
rect 1278 1116 1296 1134
rect 1278 1134 1296 1152
rect 1278 1152 1296 1170
rect 1278 1170 1296 1188
rect 1278 1188 1296 1206
rect 1278 1206 1296 1224
rect 1278 1224 1296 1242
rect 1278 1242 1296 1260
rect 1278 1260 1296 1278
rect 1278 1278 1296 1296
rect 1278 1296 1296 1314
rect 1278 1314 1296 1332
rect 1278 1332 1296 1350
rect 1278 1350 1296 1368
rect 1278 1368 1296 1386
rect 1278 1386 1296 1404
rect 1278 1404 1296 1422
rect 1278 1422 1296 1440
rect 1278 1440 1296 1458
rect 1278 1458 1296 1476
rect 1278 1476 1296 1494
rect 1278 1494 1296 1512
rect 1278 1512 1296 1530
rect 1278 1530 1296 1548
rect 1278 1548 1296 1566
rect 1278 1566 1296 1584
rect 1278 1584 1296 1602
rect 1278 1602 1296 1620
rect 1278 1620 1296 1638
rect 1278 1638 1296 1656
rect 1278 1656 1296 1674
rect 1278 1674 1296 1692
rect 1278 1692 1296 1710
rect 1278 1710 1296 1728
rect 1278 1728 1296 1746
rect 1278 1746 1296 1764
rect 1278 5508 1296 5526
rect 1278 5526 1296 5544
rect 1278 5544 1296 5562
rect 1278 5562 1296 5580
rect 1278 5580 1296 5598
rect 1278 5598 1296 5616
rect 1278 5616 1296 5634
rect 1278 5634 1296 5652
rect 1278 5652 1296 5670
rect 1278 5670 1296 5688
rect 1278 5688 1296 5706
rect 1278 5706 1296 5724
rect 1278 5724 1296 5742
rect 1278 5742 1296 5760
rect 1278 5760 1296 5778
rect 1278 5778 1296 5796
rect 1278 5796 1296 5814
rect 1278 5814 1296 5832
rect 1278 5832 1296 5850
rect 1278 5850 1296 5868
rect 1278 5868 1296 5886
rect 1278 5886 1296 5904
rect 1278 5904 1296 5922
rect 1278 5922 1296 5940
rect 1278 5940 1296 5958
rect 1278 5958 1296 5976
rect 1278 5976 1296 5994
rect 1278 5994 1296 6012
rect 1278 6012 1296 6030
rect 1278 6030 1296 6048
rect 1278 6048 1296 6066
rect 1278 6066 1296 6084
rect 1278 6084 1296 6102
rect 1278 6102 1296 6120
rect 1278 6120 1296 6138
rect 1278 6138 1296 6156
rect 1278 6156 1296 6174
rect 1278 6174 1296 6192
rect 1278 6192 1296 6210
rect 1278 6210 1296 6228
rect 1278 6228 1296 6246
rect 1278 6246 1296 6264
rect 1278 6264 1296 6282
rect 1278 6282 1296 6300
rect 1278 6300 1296 6318
rect 1278 6318 1296 6336
rect 1278 6336 1296 6354
rect 1278 6354 1296 6372
rect 1278 6372 1296 6390
rect 1278 6390 1296 6408
rect 1296 846 1314 864
rect 1296 864 1314 882
rect 1296 882 1314 900
rect 1296 900 1314 918
rect 1296 918 1314 936
rect 1296 936 1314 954
rect 1296 954 1314 972
rect 1296 972 1314 990
rect 1296 990 1314 1008
rect 1296 1008 1314 1026
rect 1296 1026 1314 1044
rect 1296 1044 1314 1062
rect 1296 1062 1314 1080
rect 1296 1080 1314 1098
rect 1296 1098 1314 1116
rect 1296 1116 1314 1134
rect 1296 1134 1314 1152
rect 1296 1152 1314 1170
rect 1296 1170 1314 1188
rect 1296 1188 1314 1206
rect 1296 1206 1314 1224
rect 1296 1224 1314 1242
rect 1296 1242 1314 1260
rect 1296 1260 1314 1278
rect 1296 1278 1314 1296
rect 1296 1296 1314 1314
rect 1296 1314 1314 1332
rect 1296 1332 1314 1350
rect 1296 1350 1314 1368
rect 1296 1368 1314 1386
rect 1296 1386 1314 1404
rect 1296 1404 1314 1422
rect 1296 1422 1314 1440
rect 1296 1440 1314 1458
rect 1296 1458 1314 1476
rect 1296 1476 1314 1494
rect 1296 1494 1314 1512
rect 1296 1512 1314 1530
rect 1296 1530 1314 1548
rect 1296 1548 1314 1566
rect 1296 1566 1314 1584
rect 1296 1584 1314 1602
rect 1296 1602 1314 1620
rect 1296 1620 1314 1638
rect 1296 1638 1314 1656
rect 1296 1656 1314 1674
rect 1296 1674 1314 1692
rect 1296 1692 1314 1710
rect 1296 1710 1314 1728
rect 1296 5544 1314 5562
rect 1296 5562 1314 5580
rect 1296 5580 1314 5598
rect 1296 5598 1314 5616
rect 1296 5616 1314 5634
rect 1296 5634 1314 5652
rect 1296 5652 1314 5670
rect 1296 5670 1314 5688
rect 1296 5688 1314 5706
rect 1296 5706 1314 5724
rect 1296 5724 1314 5742
rect 1296 5742 1314 5760
rect 1296 5760 1314 5778
rect 1296 5778 1314 5796
rect 1296 5796 1314 5814
rect 1296 5814 1314 5832
rect 1296 5832 1314 5850
rect 1296 5850 1314 5868
rect 1296 5868 1314 5886
rect 1296 5886 1314 5904
rect 1296 5904 1314 5922
rect 1296 5922 1314 5940
rect 1296 5940 1314 5958
rect 1296 5958 1314 5976
rect 1296 5976 1314 5994
rect 1296 5994 1314 6012
rect 1296 6012 1314 6030
rect 1296 6030 1314 6048
rect 1296 6048 1314 6066
rect 1296 6066 1314 6084
rect 1296 6084 1314 6102
rect 1296 6102 1314 6120
rect 1296 6120 1314 6138
rect 1296 6138 1314 6156
rect 1296 6156 1314 6174
rect 1296 6174 1314 6192
rect 1296 6192 1314 6210
rect 1296 6210 1314 6228
rect 1296 6228 1314 6246
rect 1296 6246 1314 6264
rect 1296 6264 1314 6282
rect 1296 6282 1314 6300
rect 1296 6300 1314 6318
rect 1296 6318 1314 6336
rect 1296 6336 1314 6354
rect 1296 6354 1314 6372
rect 1296 6372 1314 6390
rect 1296 6390 1314 6408
rect 1296 6408 1314 6426
rect 1314 828 1332 846
rect 1314 846 1332 864
rect 1314 864 1332 882
rect 1314 882 1332 900
rect 1314 900 1332 918
rect 1314 918 1332 936
rect 1314 936 1332 954
rect 1314 954 1332 972
rect 1314 972 1332 990
rect 1314 990 1332 1008
rect 1314 1008 1332 1026
rect 1314 1026 1332 1044
rect 1314 1044 1332 1062
rect 1314 1062 1332 1080
rect 1314 1080 1332 1098
rect 1314 1098 1332 1116
rect 1314 1116 1332 1134
rect 1314 1134 1332 1152
rect 1314 1152 1332 1170
rect 1314 1170 1332 1188
rect 1314 1188 1332 1206
rect 1314 1206 1332 1224
rect 1314 1224 1332 1242
rect 1314 1242 1332 1260
rect 1314 1260 1332 1278
rect 1314 1278 1332 1296
rect 1314 1296 1332 1314
rect 1314 1314 1332 1332
rect 1314 1332 1332 1350
rect 1314 1350 1332 1368
rect 1314 1368 1332 1386
rect 1314 1386 1332 1404
rect 1314 1404 1332 1422
rect 1314 1422 1332 1440
rect 1314 1440 1332 1458
rect 1314 1458 1332 1476
rect 1314 1476 1332 1494
rect 1314 1494 1332 1512
rect 1314 1512 1332 1530
rect 1314 1530 1332 1548
rect 1314 1548 1332 1566
rect 1314 1566 1332 1584
rect 1314 1584 1332 1602
rect 1314 1602 1332 1620
rect 1314 1620 1332 1638
rect 1314 1638 1332 1656
rect 1314 1656 1332 1674
rect 1314 1674 1332 1692
rect 1314 1692 1332 1710
rect 1314 5562 1332 5580
rect 1314 5580 1332 5598
rect 1314 5598 1332 5616
rect 1314 5616 1332 5634
rect 1314 5634 1332 5652
rect 1314 5652 1332 5670
rect 1314 5670 1332 5688
rect 1314 5688 1332 5706
rect 1314 5706 1332 5724
rect 1314 5724 1332 5742
rect 1314 5742 1332 5760
rect 1314 5760 1332 5778
rect 1314 5778 1332 5796
rect 1314 5796 1332 5814
rect 1314 5814 1332 5832
rect 1314 5832 1332 5850
rect 1314 5850 1332 5868
rect 1314 5868 1332 5886
rect 1314 5886 1332 5904
rect 1314 5904 1332 5922
rect 1314 5922 1332 5940
rect 1314 5940 1332 5958
rect 1314 5958 1332 5976
rect 1314 5976 1332 5994
rect 1314 5994 1332 6012
rect 1314 6012 1332 6030
rect 1314 6030 1332 6048
rect 1314 6048 1332 6066
rect 1314 6066 1332 6084
rect 1314 6084 1332 6102
rect 1314 6102 1332 6120
rect 1314 6120 1332 6138
rect 1314 6138 1332 6156
rect 1314 6156 1332 6174
rect 1314 6174 1332 6192
rect 1314 6192 1332 6210
rect 1314 6210 1332 6228
rect 1314 6228 1332 6246
rect 1314 6246 1332 6264
rect 1314 6264 1332 6282
rect 1314 6282 1332 6300
rect 1314 6300 1332 6318
rect 1314 6318 1332 6336
rect 1314 6336 1332 6354
rect 1314 6354 1332 6372
rect 1314 6372 1332 6390
rect 1314 6390 1332 6408
rect 1314 6408 1332 6426
rect 1314 6426 1332 6444
rect 1332 810 1350 828
rect 1332 828 1350 846
rect 1332 846 1350 864
rect 1332 864 1350 882
rect 1332 882 1350 900
rect 1332 900 1350 918
rect 1332 918 1350 936
rect 1332 936 1350 954
rect 1332 954 1350 972
rect 1332 972 1350 990
rect 1332 990 1350 1008
rect 1332 1008 1350 1026
rect 1332 1026 1350 1044
rect 1332 1044 1350 1062
rect 1332 1062 1350 1080
rect 1332 1080 1350 1098
rect 1332 1098 1350 1116
rect 1332 1116 1350 1134
rect 1332 1134 1350 1152
rect 1332 1152 1350 1170
rect 1332 1170 1350 1188
rect 1332 1188 1350 1206
rect 1332 1206 1350 1224
rect 1332 1224 1350 1242
rect 1332 1242 1350 1260
rect 1332 1260 1350 1278
rect 1332 1278 1350 1296
rect 1332 1296 1350 1314
rect 1332 1314 1350 1332
rect 1332 1332 1350 1350
rect 1332 1350 1350 1368
rect 1332 1368 1350 1386
rect 1332 1386 1350 1404
rect 1332 1404 1350 1422
rect 1332 1422 1350 1440
rect 1332 1440 1350 1458
rect 1332 1458 1350 1476
rect 1332 1476 1350 1494
rect 1332 1494 1350 1512
rect 1332 1512 1350 1530
rect 1332 1530 1350 1548
rect 1332 1548 1350 1566
rect 1332 1566 1350 1584
rect 1332 1584 1350 1602
rect 1332 1602 1350 1620
rect 1332 1620 1350 1638
rect 1332 1638 1350 1656
rect 1332 1656 1350 1674
rect 1332 1674 1350 1692
rect 1332 5580 1350 5598
rect 1332 5598 1350 5616
rect 1332 5616 1350 5634
rect 1332 5634 1350 5652
rect 1332 5652 1350 5670
rect 1332 5670 1350 5688
rect 1332 5688 1350 5706
rect 1332 5706 1350 5724
rect 1332 5724 1350 5742
rect 1332 5742 1350 5760
rect 1332 5760 1350 5778
rect 1332 5778 1350 5796
rect 1332 5796 1350 5814
rect 1332 5814 1350 5832
rect 1332 5832 1350 5850
rect 1332 5850 1350 5868
rect 1332 5868 1350 5886
rect 1332 5886 1350 5904
rect 1332 5904 1350 5922
rect 1332 5922 1350 5940
rect 1332 5940 1350 5958
rect 1332 5958 1350 5976
rect 1332 5976 1350 5994
rect 1332 5994 1350 6012
rect 1332 6012 1350 6030
rect 1332 6030 1350 6048
rect 1332 6048 1350 6066
rect 1332 6066 1350 6084
rect 1332 6084 1350 6102
rect 1332 6102 1350 6120
rect 1332 6120 1350 6138
rect 1332 6138 1350 6156
rect 1332 6156 1350 6174
rect 1332 6174 1350 6192
rect 1332 6192 1350 6210
rect 1332 6210 1350 6228
rect 1332 6228 1350 6246
rect 1332 6246 1350 6264
rect 1332 6264 1350 6282
rect 1332 6282 1350 6300
rect 1332 6300 1350 6318
rect 1332 6318 1350 6336
rect 1332 6336 1350 6354
rect 1332 6354 1350 6372
rect 1332 6372 1350 6390
rect 1332 6390 1350 6408
rect 1332 6408 1350 6426
rect 1332 6426 1350 6444
rect 1332 6444 1350 6462
rect 1350 810 1368 828
rect 1350 828 1368 846
rect 1350 846 1368 864
rect 1350 864 1368 882
rect 1350 882 1368 900
rect 1350 900 1368 918
rect 1350 918 1368 936
rect 1350 936 1368 954
rect 1350 954 1368 972
rect 1350 972 1368 990
rect 1350 990 1368 1008
rect 1350 1008 1368 1026
rect 1350 1026 1368 1044
rect 1350 1044 1368 1062
rect 1350 1062 1368 1080
rect 1350 1080 1368 1098
rect 1350 1098 1368 1116
rect 1350 1116 1368 1134
rect 1350 1134 1368 1152
rect 1350 1152 1368 1170
rect 1350 1170 1368 1188
rect 1350 1188 1368 1206
rect 1350 1206 1368 1224
rect 1350 1224 1368 1242
rect 1350 1242 1368 1260
rect 1350 1260 1368 1278
rect 1350 1278 1368 1296
rect 1350 1296 1368 1314
rect 1350 1314 1368 1332
rect 1350 1332 1368 1350
rect 1350 1350 1368 1368
rect 1350 1368 1368 1386
rect 1350 1386 1368 1404
rect 1350 1404 1368 1422
rect 1350 1422 1368 1440
rect 1350 1440 1368 1458
rect 1350 1458 1368 1476
rect 1350 1476 1368 1494
rect 1350 1494 1368 1512
rect 1350 1512 1368 1530
rect 1350 1530 1368 1548
rect 1350 1548 1368 1566
rect 1350 1566 1368 1584
rect 1350 1584 1368 1602
rect 1350 1602 1368 1620
rect 1350 1620 1368 1638
rect 1350 1638 1368 1656
rect 1350 1656 1368 1674
rect 1350 5598 1368 5616
rect 1350 5616 1368 5634
rect 1350 5634 1368 5652
rect 1350 5652 1368 5670
rect 1350 5670 1368 5688
rect 1350 5688 1368 5706
rect 1350 5706 1368 5724
rect 1350 5724 1368 5742
rect 1350 5742 1368 5760
rect 1350 5760 1368 5778
rect 1350 5778 1368 5796
rect 1350 5796 1368 5814
rect 1350 5814 1368 5832
rect 1350 5832 1368 5850
rect 1350 5850 1368 5868
rect 1350 5868 1368 5886
rect 1350 5886 1368 5904
rect 1350 5904 1368 5922
rect 1350 5922 1368 5940
rect 1350 5940 1368 5958
rect 1350 5958 1368 5976
rect 1350 5976 1368 5994
rect 1350 5994 1368 6012
rect 1350 6012 1368 6030
rect 1350 6030 1368 6048
rect 1350 6048 1368 6066
rect 1350 6066 1368 6084
rect 1350 6084 1368 6102
rect 1350 6102 1368 6120
rect 1350 6120 1368 6138
rect 1350 6138 1368 6156
rect 1350 6156 1368 6174
rect 1350 6174 1368 6192
rect 1350 6192 1368 6210
rect 1350 6210 1368 6228
rect 1350 6228 1368 6246
rect 1350 6246 1368 6264
rect 1350 6264 1368 6282
rect 1350 6282 1368 6300
rect 1350 6300 1368 6318
rect 1350 6318 1368 6336
rect 1350 6336 1368 6354
rect 1350 6354 1368 6372
rect 1350 6372 1368 6390
rect 1350 6390 1368 6408
rect 1350 6408 1368 6426
rect 1350 6426 1368 6444
rect 1350 6444 1368 6462
rect 1368 792 1386 810
rect 1368 810 1386 828
rect 1368 828 1386 846
rect 1368 846 1386 864
rect 1368 864 1386 882
rect 1368 882 1386 900
rect 1368 900 1386 918
rect 1368 918 1386 936
rect 1368 936 1386 954
rect 1368 954 1386 972
rect 1368 972 1386 990
rect 1368 990 1386 1008
rect 1368 1008 1386 1026
rect 1368 1026 1386 1044
rect 1368 1044 1386 1062
rect 1368 1062 1386 1080
rect 1368 1080 1386 1098
rect 1368 1098 1386 1116
rect 1368 1116 1386 1134
rect 1368 1134 1386 1152
rect 1368 1152 1386 1170
rect 1368 1170 1386 1188
rect 1368 1188 1386 1206
rect 1368 1206 1386 1224
rect 1368 1224 1386 1242
rect 1368 1242 1386 1260
rect 1368 1260 1386 1278
rect 1368 1278 1386 1296
rect 1368 1296 1386 1314
rect 1368 1314 1386 1332
rect 1368 1332 1386 1350
rect 1368 1350 1386 1368
rect 1368 1368 1386 1386
rect 1368 1386 1386 1404
rect 1368 1404 1386 1422
rect 1368 1422 1386 1440
rect 1368 1440 1386 1458
rect 1368 1458 1386 1476
rect 1368 1476 1386 1494
rect 1368 1494 1386 1512
rect 1368 1512 1386 1530
rect 1368 1530 1386 1548
rect 1368 1548 1386 1566
rect 1368 1566 1386 1584
rect 1368 1584 1386 1602
rect 1368 1602 1386 1620
rect 1368 1620 1386 1638
rect 1368 1638 1386 1656
rect 1368 5616 1386 5634
rect 1368 5634 1386 5652
rect 1368 5652 1386 5670
rect 1368 5670 1386 5688
rect 1368 5688 1386 5706
rect 1368 5706 1386 5724
rect 1368 5724 1386 5742
rect 1368 5742 1386 5760
rect 1368 5760 1386 5778
rect 1368 5778 1386 5796
rect 1368 5796 1386 5814
rect 1368 5814 1386 5832
rect 1368 5832 1386 5850
rect 1368 5850 1386 5868
rect 1368 5868 1386 5886
rect 1368 5886 1386 5904
rect 1368 5904 1386 5922
rect 1368 5922 1386 5940
rect 1368 5940 1386 5958
rect 1368 5958 1386 5976
rect 1368 5976 1386 5994
rect 1368 5994 1386 6012
rect 1368 6012 1386 6030
rect 1368 6030 1386 6048
rect 1368 6048 1386 6066
rect 1368 6066 1386 6084
rect 1368 6084 1386 6102
rect 1368 6102 1386 6120
rect 1368 6120 1386 6138
rect 1368 6138 1386 6156
rect 1368 6156 1386 6174
rect 1368 6174 1386 6192
rect 1368 6192 1386 6210
rect 1368 6210 1386 6228
rect 1368 6228 1386 6246
rect 1368 6246 1386 6264
rect 1368 6264 1386 6282
rect 1368 6282 1386 6300
rect 1368 6300 1386 6318
rect 1368 6318 1386 6336
rect 1368 6336 1386 6354
rect 1368 6354 1386 6372
rect 1368 6372 1386 6390
rect 1368 6390 1386 6408
rect 1368 6408 1386 6426
rect 1368 6426 1386 6444
rect 1368 6444 1386 6462
rect 1368 6462 1386 6480
rect 1386 774 1404 792
rect 1386 792 1404 810
rect 1386 810 1404 828
rect 1386 828 1404 846
rect 1386 846 1404 864
rect 1386 864 1404 882
rect 1386 882 1404 900
rect 1386 900 1404 918
rect 1386 918 1404 936
rect 1386 936 1404 954
rect 1386 954 1404 972
rect 1386 972 1404 990
rect 1386 990 1404 1008
rect 1386 1008 1404 1026
rect 1386 1026 1404 1044
rect 1386 1044 1404 1062
rect 1386 1062 1404 1080
rect 1386 1080 1404 1098
rect 1386 1098 1404 1116
rect 1386 1116 1404 1134
rect 1386 1134 1404 1152
rect 1386 1152 1404 1170
rect 1386 1170 1404 1188
rect 1386 1188 1404 1206
rect 1386 1206 1404 1224
rect 1386 1224 1404 1242
rect 1386 1242 1404 1260
rect 1386 1260 1404 1278
rect 1386 1278 1404 1296
rect 1386 1296 1404 1314
rect 1386 1314 1404 1332
rect 1386 1332 1404 1350
rect 1386 1350 1404 1368
rect 1386 1368 1404 1386
rect 1386 1386 1404 1404
rect 1386 1404 1404 1422
rect 1386 1422 1404 1440
rect 1386 1440 1404 1458
rect 1386 1458 1404 1476
rect 1386 1476 1404 1494
rect 1386 1494 1404 1512
rect 1386 1512 1404 1530
rect 1386 1530 1404 1548
rect 1386 1548 1404 1566
rect 1386 1566 1404 1584
rect 1386 1584 1404 1602
rect 1386 1602 1404 1620
rect 1386 5634 1404 5652
rect 1386 5652 1404 5670
rect 1386 5670 1404 5688
rect 1386 5688 1404 5706
rect 1386 5706 1404 5724
rect 1386 5724 1404 5742
rect 1386 5742 1404 5760
rect 1386 5760 1404 5778
rect 1386 5778 1404 5796
rect 1386 5796 1404 5814
rect 1386 5814 1404 5832
rect 1386 5832 1404 5850
rect 1386 5850 1404 5868
rect 1386 5868 1404 5886
rect 1386 5886 1404 5904
rect 1386 5904 1404 5922
rect 1386 5922 1404 5940
rect 1386 5940 1404 5958
rect 1386 5958 1404 5976
rect 1386 5976 1404 5994
rect 1386 5994 1404 6012
rect 1386 6012 1404 6030
rect 1386 6030 1404 6048
rect 1386 6048 1404 6066
rect 1386 6066 1404 6084
rect 1386 6084 1404 6102
rect 1386 6102 1404 6120
rect 1386 6120 1404 6138
rect 1386 6138 1404 6156
rect 1386 6156 1404 6174
rect 1386 6174 1404 6192
rect 1386 6192 1404 6210
rect 1386 6210 1404 6228
rect 1386 6228 1404 6246
rect 1386 6246 1404 6264
rect 1386 6264 1404 6282
rect 1386 6282 1404 6300
rect 1386 6300 1404 6318
rect 1386 6318 1404 6336
rect 1386 6336 1404 6354
rect 1386 6354 1404 6372
rect 1386 6372 1404 6390
rect 1386 6390 1404 6408
rect 1386 6408 1404 6426
rect 1386 6426 1404 6444
rect 1386 6444 1404 6462
rect 1386 6462 1404 6480
rect 1386 6480 1404 6498
rect 1404 756 1422 774
rect 1404 774 1422 792
rect 1404 792 1422 810
rect 1404 810 1422 828
rect 1404 828 1422 846
rect 1404 846 1422 864
rect 1404 864 1422 882
rect 1404 882 1422 900
rect 1404 900 1422 918
rect 1404 918 1422 936
rect 1404 936 1422 954
rect 1404 954 1422 972
rect 1404 972 1422 990
rect 1404 990 1422 1008
rect 1404 1008 1422 1026
rect 1404 1026 1422 1044
rect 1404 1044 1422 1062
rect 1404 1062 1422 1080
rect 1404 1080 1422 1098
rect 1404 1098 1422 1116
rect 1404 1116 1422 1134
rect 1404 1134 1422 1152
rect 1404 1152 1422 1170
rect 1404 1170 1422 1188
rect 1404 1188 1422 1206
rect 1404 1206 1422 1224
rect 1404 1224 1422 1242
rect 1404 1242 1422 1260
rect 1404 1260 1422 1278
rect 1404 1278 1422 1296
rect 1404 1296 1422 1314
rect 1404 1314 1422 1332
rect 1404 1332 1422 1350
rect 1404 1350 1422 1368
rect 1404 1368 1422 1386
rect 1404 1386 1422 1404
rect 1404 1404 1422 1422
rect 1404 1422 1422 1440
rect 1404 1440 1422 1458
rect 1404 1458 1422 1476
rect 1404 1476 1422 1494
rect 1404 1494 1422 1512
rect 1404 1512 1422 1530
rect 1404 1530 1422 1548
rect 1404 1548 1422 1566
rect 1404 1566 1422 1584
rect 1404 1584 1422 1602
rect 1404 5670 1422 5688
rect 1404 5688 1422 5706
rect 1404 5706 1422 5724
rect 1404 5724 1422 5742
rect 1404 5742 1422 5760
rect 1404 5760 1422 5778
rect 1404 5778 1422 5796
rect 1404 5796 1422 5814
rect 1404 5814 1422 5832
rect 1404 5832 1422 5850
rect 1404 5850 1422 5868
rect 1404 5868 1422 5886
rect 1404 5886 1422 5904
rect 1404 5904 1422 5922
rect 1404 5922 1422 5940
rect 1404 5940 1422 5958
rect 1404 5958 1422 5976
rect 1404 5976 1422 5994
rect 1404 5994 1422 6012
rect 1404 6012 1422 6030
rect 1404 6030 1422 6048
rect 1404 6048 1422 6066
rect 1404 6066 1422 6084
rect 1404 6084 1422 6102
rect 1404 6102 1422 6120
rect 1404 6120 1422 6138
rect 1404 6138 1422 6156
rect 1404 6156 1422 6174
rect 1404 6174 1422 6192
rect 1404 6192 1422 6210
rect 1404 6210 1422 6228
rect 1404 6228 1422 6246
rect 1404 6246 1422 6264
rect 1404 6264 1422 6282
rect 1404 6282 1422 6300
rect 1404 6300 1422 6318
rect 1404 6318 1422 6336
rect 1404 6336 1422 6354
rect 1404 6354 1422 6372
rect 1404 6372 1422 6390
rect 1404 6390 1422 6408
rect 1404 6408 1422 6426
rect 1404 6426 1422 6444
rect 1404 6444 1422 6462
rect 1404 6462 1422 6480
rect 1404 6480 1422 6498
rect 1404 6498 1422 6516
rect 1422 738 1440 756
rect 1422 756 1440 774
rect 1422 774 1440 792
rect 1422 792 1440 810
rect 1422 810 1440 828
rect 1422 828 1440 846
rect 1422 846 1440 864
rect 1422 864 1440 882
rect 1422 882 1440 900
rect 1422 900 1440 918
rect 1422 918 1440 936
rect 1422 936 1440 954
rect 1422 954 1440 972
rect 1422 972 1440 990
rect 1422 990 1440 1008
rect 1422 1008 1440 1026
rect 1422 1026 1440 1044
rect 1422 1044 1440 1062
rect 1422 1062 1440 1080
rect 1422 1080 1440 1098
rect 1422 1098 1440 1116
rect 1422 1116 1440 1134
rect 1422 1134 1440 1152
rect 1422 1152 1440 1170
rect 1422 1170 1440 1188
rect 1422 1188 1440 1206
rect 1422 1206 1440 1224
rect 1422 1224 1440 1242
rect 1422 1242 1440 1260
rect 1422 1260 1440 1278
rect 1422 1278 1440 1296
rect 1422 1296 1440 1314
rect 1422 1314 1440 1332
rect 1422 1332 1440 1350
rect 1422 1350 1440 1368
rect 1422 1368 1440 1386
rect 1422 1386 1440 1404
rect 1422 1404 1440 1422
rect 1422 1422 1440 1440
rect 1422 1440 1440 1458
rect 1422 1458 1440 1476
rect 1422 1476 1440 1494
rect 1422 1494 1440 1512
rect 1422 1512 1440 1530
rect 1422 1530 1440 1548
rect 1422 1548 1440 1566
rect 1422 1566 1440 1584
rect 1422 5688 1440 5706
rect 1422 5706 1440 5724
rect 1422 5724 1440 5742
rect 1422 5742 1440 5760
rect 1422 5760 1440 5778
rect 1422 5778 1440 5796
rect 1422 5796 1440 5814
rect 1422 5814 1440 5832
rect 1422 5832 1440 5850
rect 1422 5850 1440 5868
rect 1422 5868 1440 5886
rect 1422 5886 1440 5904
rect 1422 5904 1440 5922
rect 1422 5922 1440 5940
rect 1422 5940 1440 5958
rect 1422 5958 1440 5976
rect 1422 5976 1440 5994
rect 1422 5994 1440 6012
rect 1422 6012 1440 6030
rect 1422 6030 1440 6048
rect 1422 6048 1440 6066
rect 1422 6066 1440 6084
rect 1422 6084 1440 6102
rect 1422 6102 1440 6120
rect 1422 6120 1440 6138
rect 1422 6138 1440 6156
rect 1422 6156 1440 6174
rect 1422 6174 1440 6192
rect 1422 6192 1440 6210
rect 1422 6210 1440 6228
rect 1422 6228 1440 6246
rect 1422 6246 1440 6264
rect 1422 6264 1440 6282
rect 1422 6282 1440 6300
rect 1422 6300 1440 6318
rect 1422 6318 1440 6336
rect 1422 6336 1440 6354
rect 1422 6354 1440 6372
rect 1422 6372 1440 6390
rect 1422 6390 1440 6408
rect 1422 6408 1440 6426
rect 1422 6426 1440 6444
rect 1422 6444 1440 6462
rect 1422 6462 1440 6480
rect 1422 6480 1440 6498
rect 1422 6498 1440 6516
rect 1440 738 1458 756
rect 1440 756 1458 774
rect 1440 774 1458 792
rect 1440 792 1458 810
rect 1440 810 1458 828
rect 1440 828 1458 846
rect 1440 846 1458 864
rect 1440 864 1458 882
rect 1440 882 1458 900
rect 1440 900 1458 918
rect 1440 918 1458 936
rect 1440 936 1458 954
rect 1440 954 1458 972
rect 1440 972 1458 990
rect 1440 990 1458 1008
rect 1440 1008 1458 1026
rect 1440 1026 1458 1044
rect 1440 1044 1458 1062
rect 1440 1062 1458 1080
rect 1440 1080 1458 1098
rect 1440 1098 1458 1116
rect 1440 1116 1458 1134
rect 1440 1134 1458 1152
rect 1440 1152 1458 1170
rect 1440 1170 1458 1188
rect 1440 1188 1458 1206
rect 1440 1206 1458 1224
rect 1440 1224 1458 1242
rect 1440 1242 1458 1260
rect 1440 1260 1458 1278
rect 1440 1278 1458 1296
rect 1440 1296 1458 1314
rect 1440 1314 1458 1332
rect 1440 1332 1458 1350
rect 1440 1350 1458 1368
rect 1440 1368 1458 1386
rect 1440 1386 1458 1404
rect 1440 1404 1458 1422
rect 1440 1422 1458 1440
rect 1440 1440 1458 1458
rect 1440 1458 1458 1476
rect 1440 1476 1458 1494
rect 1440 1494 1458 1512
rect 1440 1512 1458 1530
rect 1440 1530 1458 1548
rect 1440 1548 1458 1566
rect 1440 5706 1458 5724
rect 1440 5724 1458 5742
rect 1440 5742 1458 5760
rect 1440 5760 1458 5778
rect 1440 5778 1458 5796
rect 1440 5796 1458 5814
rect 1440 5814 1458 5832
rect 1440 5832 1458 5850
rect 1440 5850 1458 5868
rect 1440 5868 1458 5886
rect 1440 5886 1458 5904
rect 1440 5904 1458 5922
rect 1440 5922 1458 5940
rect 1440 5940 1458 5958
rect 1440 5958 1458 5976
rect 1440 5976 1458 5994
rect 1440 5994 1458 6012
rect 1440 6012 1458 6030
rect 1440 6030 1458 6048
rect 1440 6048 1458 6066
rect 1440 6066 1458 6084
rect 1440 6084 1458 6102
rect 1440 6102 1458 6120
rect 1440 6120 1458 6138
rect 1440 6138 1458 6156
rect 1440 6156 1458 6174
rect 1440 6174 1458 6192
rect 1440 6192 1458 6210
rect 1440 6210 1458 6228
rect 1440 6228 1458 6246
rect 1440 6246 1458 6264
rect 1440 6264 1458 6282
rect 1440 6282 1458 6300
rect 1440 6300 1458 6318
rect 1440 6318 1458 6336
rect 1440 6336 1458 6354
rect 1440 6354 1458 6372
rect 1440 6372 1458 6390
rect 1440 6390 1458 6408
rect 1440 6408 1458 6426
rect 1440 6426 1458 6444
rect 1440 6444 1458 6462
rect 1440 6462 1458 6480
rect 1440 6480 1458 6498
rect 1440 6498 1458 6516
rect 1440 6516 1458 6534
rect 1458 720 1476 738
rect 1458 738 1476 756
rect 1458 756 1476 774
rect 1458 774 1476 792
rect 1458 792 1476 810
rect 1458 810 1476 828
rect 1458 828 1476 846
rect 1458 846 1476 864
rect 1458 864 1476 882
rect 1458 882 1476 900
rect 1458 900 1476 918
rect 1458 918 1476 936
rect 1458 936 1476 954
rect 1458 954 1476 972
rect 1458 972 1476 990
rect 1458 990 1476 1008
rect 1458 1008 1476 1026
rect 1458 1026 1476 1044
rect 1458 1044 1476 1062
rect 1458 1062 1476 1080
rect 1458 1080 1476 1098
rect 1458 1098 1476 1116
rect 1458 1116 1476 1134
rect 1458 1134 1476 1152
rect 1458 1152 1476 1170
rect 1458 1170 1476 1188
rect 1458 1188 1476 1206
rect 1458 1206 1476 1224
rect 1458 1224 1476 1242
rect 1458 1242 1476 1260
rect 1458 1260 1476 1278
rect 1458 1278 1476 1296
rect 1458 1296 1476 1314
rect 1458 1314 1476 1332
rect 1458 1332 1476 1350
rect 1458 1350 1476 1368
rect 1458 1368 1476 1386
rect 1458 1386 1476 1404
rect 1458 1404 1476 1422
rect 1458 1422 1476 1440
rect 1458 1440 1476 1458
rect 1458 1458 1476 1476
rect 1458 1476 1476 1494
rect 1458 1494 1476 1512
rect 1458 1512 1476 1530
rect 1458 1530 1476 1548
rect 1458 5724 1476 5742
rect 1458 5742 1476 5760
rect 1458 5760 1476 5778
rect 1458 5778 1476 5796
rect 1458 5796 1476 5814
rect 1458 5814 1476 5832
rect 1458 5832 1476 5850
rect 1458 5850 1476 5868
rect 1458 5868 1476 5886
rect 1458 5886 1476 5904
rect 1458 5904 1476 5922
rect 1458 5922 1476 5940
rect 1458 5940 1476 5958
rect 1458 5958 1476 5976
rect 1458 5976 1476 5994
rect 1458 5994 1476 6012
rect 1458 6012 1476 6030
rect 1458 6030 1476 6048
rect 1458 6048 1476 6066
rect 1458 6066 1476 6084
rect 1458 6084 1476 6102
rect 1458 6102 1476 6120
rect 1458 6120 1476 6138
rect 1458 6138 1476 6156
rect 1458 6156 1476 6174
rect 1458 6174 1476 6192
rect 1458 6192 1476 6210
rect 1458 6210 1476 6228
rect 1458 6228 1476 6246
rect 1458 6246 1476 6264
rect 1458 6264 1476 6282
rect 1458 6282 1476 6300
rect 1458 6300 1476 6318
rect 1458 6318 1476 6336
rect 1458 6336 1476 6354
rect 1458 6354 1476 6372
rect 1458 6372 1476 6390
rect 1458 6390 1476 6408
rect 1458 6408 1476 6426
rect 1458 6426 1476 6444
rect 1458 6444 1476 6462
rect 1458 6462 1476 6480
rect 1458 6480 1476 6498
rect 1458 6498 1476 6516
rect 1458 6516 1476 6534
rect 1458 6534 1476 6552
rect 1476 702 1494 720
rect 1476 720 1494 738
rect 1476 738 1494 756
rect 1476 756 1494 774
rect 1476 774 1494 792
rect 1476 792 1494 810
rect 1476 810 1494 828
rect 1476 828 1494 846
rect 1476 846 1494 864
rect 1476 864 1494 882
rect 1476 882 1494 900
rect 1476 900 1494 918
rect 1476 918 1494 936
rect 1476 936 1494 954
rect 1476 954 1494 972
rect 1476 972 1494 990
rect 1476 990 1494 1008
rect 1476 1008 1494 1026
rect 1476 1026 1494 1044
rect 1476 1044 1494 1062
rect 1476 1062 1494 1080
rect 1476 1080 1494 1098
rect 1476 1098 1494 1116
rect 1476 1116 1494 1134
rect 1476 1134 1494 1152
rect 1476 1152 1494 1170
rect 1476 1170 1494 1188
rect 1476 1188 1494 1206
rect 1476 1206 1494 1224
rect 1476 1224 1494 1242
rect 1476 1242 1494 1260
rect 1476 1260 1494 1278
rect 1476 1278 1494 1296
rect 1476 1296 1494 1314
rect 1476 1314 1494 1332
rect 1476 1332 1494 1350
rect 1476 1350 1494 1368
rect 1476 1368 1494 1386
rect 1476 1386 1494 1404
rect 1476 1404 1494 1422
rect 1476 1422 1494 1440
rect 1476 1440 1494 1458
rect 1476 1458 1494 1476
rect 1476 1476 1494 1494
rect 1476 1494 1494 1512
rect 1476 1512 1494 1530
rect 1476 5742 1494 5760
rect 1476 5760 1494 5778
rect 1476 5778 1494 5796
rect 1476 5796 1494 5814
rect 1476 5814 1494 5832
rect 1476 5832 1494 5850
rect 1476 5850 1494 5868
rect 1476 5868 1494 5886
rect 1476 5886 1494 5904
rect 1476 5904 1494 5922
rect 1476 5922 1494 5940
rect 1476 5940 1494 5958
rect 1476 5958 1494 5976
rect 1476 5976 1494 5994
rect 1476 5994 1494 6012
rect 1476 6012 1494 6030
rect 1476 6030 1494 6048
rect 1476 6048 1494 6066
rect 1476 6066 1494 6084
rect 1476 6084 1494 6102
rect 1476 6102 1494 6120
rect 1476 6120 1494 6138
rect 1476 6138 1494 6156
rect 1476 6156 1494 6174
rect 1476 6174 1494 6192
rect 1476 6192 1494 6210
rect 1476 6210 1494 6228
rect 1476 6228 1494 6246
rect 1476 6246 1494 6264
rect 1476 6264 1494 6282
rect 1476 6282 1494 6300
rect 1476 6300 1494 6318
rect 1476 6318 1494 6336
rect 1476 6336 1494 6354
rect 1476 6354 1494 6372
rect 1476 6372 1494 6390
rect 1476 6390 1494 6408
rect 1476 6408 1494 6426
rect 1476 6426 1494 6444
rect 1476 6444 1494 6462
rect 1476 6462 1494 6480
rect 1476 6480 1494 6498
rect 1476 6498 1494 6516
rect 1476 6516 1494 6534
rect 1476 6534 1494 6552
rect 1476 6552 1494 6570
rect 1494 684 1512 702
rect 1494 702 1512 720
rect 1494 720 1512 738
rect 1494 738 1512 756
rect 1494 756 1512 774
rect 1494 774 1512 792
rect 1494 792 1512 810
rect 1494 810 1512 828
rect 1494 828 1512 846
rect 1494 846 1512 864
rect 1494 864 1512 882
rect 1494 882 1512 900
rect 1494 900 1512 918
rect 1494 918 1512 936
rect 1494 936 1512 954
rect 1494 954 1512 972
rect 1494 972 1512 990
rect 1494 990 1512 1008
rect 1494 1008 1512 1026
rect 1494 1026 1512 1044
rect 1494 1044 1512 1062
rect 1494 1062 1512 1080
rect 1494 1080 1512 1098
rect 1494 1098 1512 1116
rect 1494 1116 1512 1134
rect 1494 1134 1512 1152
rect 1494 1152 1512 1170
rect 1494 1170 1512 1188
rect 1494 1188 1512 1206
rect 1494 1206 1512 1224
rect 1494 1224 1512 1242
rect 1494 1242 1512 1260
rect 1494 1260 1512 1278
rect 1494 1278 1512 1296
rect 1494 1296 1512 1314
rect 1494 1314 1512 1332
rect 1494 1332 1512 1350
rect 1494 1350 1512 1368
rect 1494 1368 1512 1386
rect 1494 1386 1512 1404
rect 1494 1404 1512 1422
rect 1494 1422 1512 1440
rect 1494 1440 1512 1458
rect 1494 1458 1512 1476
rect 1494 1476 1512 1494
rect 1494 1494 1512 1512
rect 1494 5760 1512 5778
rect 1494 5778 1512 5796
rect 1494 5796 1512 5814
rect 1494 5814 1512 5832
rect 1494 5832 1512 5850
rect 1494 5850 1512 5868
rect 1494 5868 1512 5886
rect 1494 5886 1512 5904
rect 1494 5904 1512 5922
rect 1494 5922 1512 5940
rect 1494 5940 1512 5958
rect 1494 5958 1512 5976
rect 1494 5976 1512 5994
rect 1494 5994 1512 6012
rect 1494 6012 1512 6030
rect 1494 6030 1512 6048
rect 1494 6048 1512 6066
rect 1494 6066 1512 6084
rect 1494 6084 1512 6102
rect 1494 6102 1512 6120
rect 1494 6120 1512 6138
rect 1494 6138 1512 6156
rect 1494 6156 1512 6174
rect 1494 6174 1512 6192
rect 1494 6192 1512 6210
rect 1494 6210 1512 6228
rect 1494 6228 1512 6246
rect 1494 6246 1512 6264
rect 1494 6264 1512 6282
rect 1494 6282 1512 6300
rect 1494 6300 1512 6318
rect 1494 6318 1512 6336
rect 1494 6336 1512 6354
rect 1494 6354 1512 6372
rect 1494 6372 1512 6390
rect 1494 6390 1512 6408
rect 1494 6408 1512 6426
rect 1494 6426 1512 6444
rect 1494 6444 1512 6462
rect 1494 6462 1512 6480
rect 1494 6480 1512 6498
rect 1494 6498 1512 6516
rect 1494 6516 1512 6534
rect 1494 6534 1512 6552
rect 1494 6552 1512 6570
rect 1512 684 1530 702
rect 1512 702 1530 720
rect 1512 720 1530 738
rect 1512 738 1530 756
rect 1512 756 1530 774
rect 1512 774 1530 792
rect 1512 792 1530 810
rect 1512 810 1530 828
rect 1512 828 1530 846
rect 1512 846 1530 864
rect 1512 864 1530 882
rect 1512 882 1530 900
rect 1512 900 1530 918
rect 1512 918 1530 936
rect 1512 936 1530 954
rect 1512 954 1530 972
rect 1512 972 1530 990
rect 1512 990 1530 1008
rect 1512 1008 1530 1026
rect 1512 1026 1530 1044
rect 1512 1044 1530 1062
rect 1512 1062 1530 1080
rect 1512 1080 1530 1098
rect 1512 1098 1530 1116
rect 1512 1116 1530 1134
rect 1512 1134 1530 1152
rect 1512 1152 1530 1170
rect 1512 1170 1530 1188
rect 1512 1188 1530 1206
rect 1512 1206 1530 1224
rect 1512 1224 1530 1242
rect 1512 1242 1530 1260
rect 1512 1260 1530 1278
rect 1512 1278 1530 1296
rect 1512 1296 1530 1314
rect 1512 1314 1530 1332
rect 1512 1332 1530 1350
rect 1512 1350 1530 1368
rect 1512 1368 1530 1386
rect 1512 1386 1530 1404
rect 1512 1404 1530 1422
rect 1512 1422 1530 1440
rect 1512 1440 1530 1458
rect 1512 1458 1530 1476
rect 1512 1476 1530 1494
rect 1512 5778 1530 5796
rect 1512 5796 1530 5814
rect 1512 5814 1530 5832
rect 1512 5832 1530 5850
rect 1512 5850 1530 5868
rect 1512 5868 1530 5886
rect 1512 5886 1530 5904
rect 1512 5904 1530 5922
rect 1512 5922 1530 5940
rect 1512 5940 1530 5958
rect 1512 5958 1530 5976
rect 1512 5976 1530 5994
rect 1512 5994 1530 6012
rect 1512 6012 1530 6030
rect 1512 6030 1530 6048
rect 1512 6048 1530 6066
rect 1512 6066 1530 6084
rect 1512 6084 1530 6102
rect 1512 6102 1530 6120
rect 1512 6120 1530 6138
rect 1512 6138 1530 6156
rect 1512 6156 1530 6174
rect 1512 6174 1530 6192
rect 1512 6192 1530 6210
rect 1512 6210 1530 6228
rect 1512 6228 1530 6246
rect 1512 6246 1530 6264
rect 1512 6264 1530 6282
rect 1512 6282 1530 6300
rect 1512 6300 1530 6318
rect 1512 6318 1530 6336
rect 1512 6336 1530 6354
rect 1512 6354 1530 6372
rect 1512 6372 1530 6390
rect 1512 6390 1530 6408
rect 1512 6408 1530 6426
rect 1512 6426 1530 6444
rect 1512 6444 1530 6462
rect 1512 6462 1530 6480
rect 1512 6480 1530 6498
rect 1512 6498 1530 6516
rect 1512 6516 1530 6534
rect 1512 6534 1530 6552
rect 1512 6552 1530 6570
rect 1512 6570 1530 6588
rect 1530 666 1548 684
rect 1530 684 1548 702
rect 1530 702 1548 720
rect 1530 720 1548 738
rect 1530 738 1548 756
rect 1530 756 1548 774
rect 1530 774 1548 792
rect 1530 792 1548 810
rect 1530 810 1548 828
rect 1530 828 1548 846
rect 1530 846 1548 864
rect 1530 864 1548 882
rect 1530 882 1548 900
rect 1530 900 1548 918
rect 1530 918 1548 936
rect 1530 936 1548 954
rect 1530 954 1548 972
rect 1530 972 1548 990
rect 1530 990 1548 1008
rect 1530 1008 1548 1026
rect 1530 1026 1548 1044
rect 1530 1044 1548 1062
rect 1530 1062 1548 1080
rect 1530 1080 1548 1098
rect 1530 1098 1548 1116
rect 1530 1116 1548 1134
rect 1530 1134 1548 1152
rect 1530 1152 1548 1170
rect 1530 1170 1548 1188
rect 1530 1188 1548 1206
rect 1530 1206 1548 1224
rect 1530 1224 1548 1242
rect 1530 1242 1548 1260
rect 1530 1260 1548 1278
rect 1530 1278 1548 1296
rect 1530 1296 1548 1314
rect 1530 1314 1548 1332
rect 1530 1332 1548 1350
rect 1530 1350 1548 1368
rect 1530 1368 1548 1386
rect 1530 1386 1548 1404
rect 1530 1404 1548 1422
rect 1530 1422 1548 1440
rect 1530 1440 1548 1458
rect 1530 1458 1548 1476
rect 1530 5796 1548 5814
rect 1530 5814 1548 5832
rect 1530 5832 1548 5850
rect 1530 5850 1548 5868
rect 1530 5868 1548 5886
rect 1530 5886 1548 5904
rect 1530 5904 1548 5922
rect 1530 5922 1548 5940
rect 1530 5940 1548 5958
rect 1530 5958 1548 5976
rect 1530 5976 1548 5994
rect 1530 5994 1548 6012
rect 1530 6012 1548 6030
rect 1530 6030 1548 6048
rect 1530 6048 1548 6066
rect 1530 6066 1548 6084
rect 1530 6084 1548 6102
rect 1530 6102 1548 6120
rect 1530 6120 1548 6138
rect 1530 6138 1548 6156
rect 1530 6156 1548 6174
rect 1530 6174 1548 6192
rect 1530 6192 1548 6210
rect 1530 6210 1548 6228
rect 1530 6228 1548 6246
rect 1530 6246 1548 6264
rect 1530 6264 1548 6282
rect 1530 6282 1548 6300
rect 1530 6300 1548 6318
rect 1530 6318 1548 6336
rect 1530 6336 1548 6354
rect 1530 6354 1548 6372
rect 1530 6372 1548 6390
rect 1530 6390 1548 6408
rect 1530 6408 1548 6426
rect 1530 6426 1548 6444
rect 1530 6444 1548 6462
rect 1530 6462 1548 6480
rect 1530 6480 1548 6498
rect 1530 6498 1548 6516
rect 1530 6516 1548 6534
rect 1530 6534 1548 6552
rect 1530 6552 1548 6570
rect 1530 6570 1548 6588
rect 1530 6588 1548 6606
rect 1548 648 1566 666
rect 1548 666 1566 684
rect 1548 684 1566 702
rect 1548 702 1566 720
rect 1548 720 1566 738
rect 1548 738 1566 756
rect 1548 756 1566 774
rect 1548 774 1566 792
rect 1548 792 1566 810
rect 1548 810 1566 828
rect 1548 828 1566 846
rect 1548 846 1566 864
rect 1548 864 1566 882
rect 1548 882 1566 900
rect 1548 900 1566 918
rect 1548 918 1566 936
rect 1548 936 1566 954
rect 1548 954 1566 972
rect 1548 972 1566 990
rect 1548 990 1566 1008
rect 1548 1008 1566 1026
rect 1548 1026 1566 1044
rect 1548 1044 1566 1062
rect 1548 1062 1566 1080
rect 1548 1080 1566 1098
rect 1548 1098 1566 1116
rect 1548 1116 1566 1134
rect 1548 1134 1566 1152
rect 1548 1152 1566 1170
rect 1548 1170 1566 1188
rect 1548 1188 1566 1206
rect 1548 1206 1566 1224
rect 1548 1224 1566 1242
rect 1548 1242 1566 1260
rect 1548 1260 1566 1278
rect 1548 1278 1566 1296
rect 1548 1296 1566 1314
rect 1548 1314 1566 1332
rect 1548 1332 1566 1350
rect 1548 1350 1566 1368
rect 1548 1368 1566 1386
rect 1548 1386 1566 1404
rect 1548 1404 1566 1422
rect 1548 1422 1566 1440
rect 1548 1440 1566 1458
rect 1548 5814 1566 5832
rect 1548 5832 1566 5850
rect 1548 5850 1566 5868
rect 1548 5868 1566 5886
rect 1548 5886 1566 5904
rect 1548 5904 1566 5922
rect 1548 5922 1566 5940
rect 1548 5940 1566 5958
rect 1548 5958 1566 5976
rect 1548 5976 1566 5994
rect 1548 5994 1566 6012
rect 1548 6012 1566 6030
rect 1548 6030 1566 6048
rect 1548 6048 1566 6066
rect 1548 6066 1566 6084
rect 1548 6084 1566 6102
rect 1548 6102 1566 6120
rect 1548 6120 1566 6138
rect 1548 6138 1566 6156
rect 1548 6156 1566 6174
rect 1548 6174 1566 6192
rect 1548 6192 1566 6210
rect 1548 6210 1566 6228
rect 1548 6228 1566 6246
rect 1548 6246 1566 6264
rect 1548 6264 1566 6282
rect 1548 6282 1566 6300
rect 1548 6300 1566 6318
rect 1548 6318 1566 6336
rect 1548 6336 1566 6354
rect 1548 6354 1566 6372
rect 1548 6372 1566 6390
rect 1548 6390 1566 6408
rect 1548 6408 1566 6426
rect 1548 6426 1566 6444
rect 1548 6444 1566 6462
rect 1548 6462 1566 6480
rect 1548 6480 1566 6498
rect 1548 6498 1566 6516
rect 1548 6516 1566 6534
rect 1548 6534 1566 6552
rect 1548 6552 1566 6570
rect 1548 6570 1566 6588
rect 1548 6588 1566 6606
rect 1548 6606 1566 6624
rect 1566 648 1584 666
rect 1566 666 1584 684
rect 1566 684 1584 702
rect 1566 702 1584 720
rect 1566 720 1584 738
rect 1566 738 1584 756
rect 1566 756 1584 774
rect 1566 774 1584 792
rect 1566 792 1584 810
rect 1566 810 1584 828
rect 1566 828 1584 846
rect 1566 846 1584 864
rect 1566 864 1584 882
rect 1566 882 1584 900
rect 1566 900 1584 918
rect 1566 918 1584 936
rect 1566 936 1584 954
rect 1566 954 1584 972
rect 1566 972 1584 990
rect 1566 990 1584 1008
rect 1566 1008 1584 1026
rect 1566 1026 1584 1044
rect 1566 1044 1584 1062
rect 1566 1062 1584 1080
rect 1566 1080 1584 1098
rect 1566 1098 1584 1116
rect 1566 1116 1584 1134
rect 1566 1134 1584 1152
rect 1566 1152 1584 1170
rect 1566 1170 1584 1188
rect 1566 1188 1584 1206
rect 1566 1206 1584 1224
rect 1566 1224 1584 1242
rect 1566 1242 1584 1260
rect 1566 1260 1584 1278
rect 1566 1278 1584 1296
rect 1566 1296 1584 1314
rect 1566 1314 1584 1332
rect 1566 1332 1584 1350
rect 1566 1350 1584 1368
rect 1566 1368 1584 1386
rect 1566 1386 1584 1404
rect 1566 1404 1584 1422
rect 1566 1422 1584 1440
rect 1566 5832 1584 5850
rect 1566 5850 1584 5868
rect 1566 5868 1584 5886
rect 1566 5886 1584 5904
rect 1566 5904 1584 5922
rect 1566 5922 1584 5940
rect 1566 5940 1584 5958
rect 1566 5958 1584 5976
rect 1566 5976 1584 5994
rect 1566 5994 1584 6012
rect 1566 6012 1584 6030
rect 1566 6030 1584 6048
rect 1566 6048 1584 6066
rect 1566 6066 1584 6084
rect 1566 6084 1584 6102
rect 1566 6102 1584 6120
rect 1566 6120 1584 6138
rect 1566 6138 1584 6156
rect 1566 6156 1584 6174
rect 1566 6174 1584 6192
rect 1566 6192 1584 6210
rect 1566 6210 1584 6228
rect 1566 6228 1584 6246
rect 1566 6246 1584 6264
rect 1566 6264 1584 6282
rect 1566 6282 1584 6300
rect 1566 6300 1584 6318
rect 1566 6318 1584 6336
rect 1566 6336 1584 6354
rect 1566 6354 1584 6372
rect 1566 6372 1584 6390
rect 1566 6390 1584 6408
rect 1566 6408 1584 6426
rect 1566 6426 1584 6444
rect 1566 6444 1584 6462
rect 1566 6462 1584 6480
rect 1566 6480 1584 6498
rect 1566 6498 1584 6516
rect 1566 6516 1584 6534
rect 1566 6534 1584 6552
rect 1566 6552 1584 6570
rect 1566 6570 1584 6588
rect 1566 6588 1584 6606
rect 1566 6606 1584 6624
rect 1584 630 1602 648
rect 1584 648 1602 666
rect 1584 666 1602 684
rect 1584 684 1602 702
rect 1584 702 1602 720
rect 1584 720 1602 738
rect 1584 738 1602 756
rect 1584 756 1602 774
rect 1584 774 1602 792
rect 1584 792 1602 810
rect 1584 810 1602 828
rect 1584 828 1602 846
rect 1584 846 1602 864
rect 1584 864 1602 882
rect 1584 882 1602 900
rect 1584 900 1602 918
rect 1584 918 1602 936
rect 1584 936 1602 954
rect 1584 954 1602 972
rect 1584 972 1602 990
rect 1584 990 1602 1008
rect 1584 1008 1602 1026
rect 1584 1026 1602 1044
rect 1584 1044 1602 1062
rect 1584 1062 1602 1080
rect 1584 1080 1602 1098
rect 1584 1098 1602 1116
rect 1584 1116 1602 1134
rect 1584 1134 1602 1152
rect 1584 1152 1602 1170
rect 1584 1170 1602 1188
rect 1584 1188 1602 1206
rect 1584 1206 1602 1224
rect 1584 1224 1602 1242
rect 1584 1242 1602 1260
rect 1584 1260 1602 1278
rect 1584 1278 1602 1296
rect 1584 1296 1602 1314
rect 1584 1314 1602 1332
rect 1584 1332 1602 1350
rect 1584 1350 1602 1368
rect 1584 1368 1602 1386
rect 1584 1386 1602 1404
rect 1584 1404 1602 1422
rect 1584 5850 1602 5868
rect 1584 5868 1602 5886
rect 1584 5886 1602 5904
rect 1584 5904 1602 5922
rect 1584 5922 1602 5940
rect 1584 5940 1602 5958
rect 1584 5958 1602 5976
rect 1584 5976 1602 5994
rect 1584 5994 1602 6012
rect 1584 6012 1602 6030
rect 1584 6030 1602 6048
rect 1584 6048 1602 6066
rect 1584 6066 1602 6084
rect 1584 6084 1602 6102
rect 1584 6102 1602 6120
rect 1584 6120 1602 6138
rect 1584 6138 1602 6156
rect 1584 6156 1602 6174
rect 1584 6174 1602 6192
rect 1584 6192 1602 6210
rect 1584 6210 1602 6228
rect 1584 6228 1602 6246
rect 1584 6246 1602 6264
rect 1584 6264 1602 6282
rect 1584 6282 1602 6300
rect 1584 6300 1602 6318
rect 1584 6318 1602 6336
rect 1584 6336 1602 6354
rect 1584 6354 1602 6372
rect 1584 6372 1602 6390
rect 1584 6390 1602 6408
rect 1584 6408 1602 6426
rect 1584 6426 1602 6444
rect 1584 6444 1602 6462
rect 1584 6462 1602 6480
rect 1584 6480 1602 6498
rect 1584 6498 1602 6516
rect 1584 6516 1602 6534
rect 1584 6534 1602 6552
rect 1584 6552 1602 6570
rect 1584 6570 1602 6588
rect 1584 6588 1602 6606
rect 1584 6606 1602 6624
rect 1584 6624 1602 6642
rect 1602 612 1620 630
rect 1602 630 1620 648
rect 1602 648 1620 666
rect 1602 666 1620 684
rect 1602 684 1620 702
rect 1602 702 1620 720
rect 1602 720 1620 738
rect 1602 738 1620 756
rect 1602 756 1620 774
rect 1602 774 1620 792
rect 1602 792 1620 810
rect 1602 810 1620 828
rect 1602 828 1620 846
rect 1602 846 1620 864
rect 1602 864 1620 882
rect 1602 882 1620 900
rect 1602 900 1620 918
rect 1602 918 1620 936
rect 1602 936 1620 954
rect 1602 954 1620 972
rect 1602 972 1620 990
rect 1602 990 1620 1008
rect 1602 1008 1620 1026
rect 1602 1026 1620 1044
rect 1602 1044 1620 1062
rect 1602 1062 1620 1080
rect 1602 1080 1620 1098
rect 1602 1098 1620 1116
rect 1602 1116 1620 1134
rect 1602 1134 1620 1152
rect 1602 1152 1620 1170
rect 1602 1170 1620 1188
rect 1602 1188 1620 1206
rect 1602 1206 1620 1224
rect 1602 1224 1620 1242
rect 1602 1242 1620 1260
rect 1602 1260 1620 1278
rect 1602 1278 1620 1296
rect 1602 1296 1620 1314
rect 1602 1314 1620 1332
rect 1602 1332 1620 1350
rect 1602 1350 1620 1368
rect 1602 1368 1620 1386
rect 1602 1386 1620 1404
rect 1602 5868 1620 5886
rect 1602 5886 1620 5904
rect 1602 5904 1620 5922
rect 1602 5922 1620 5940
rect 1602 5940 1620 5958
rect 1602 5958 1620 5976
rect 1602 5976 1620 5994
rect 1602 5994 1620 6012
rect 1602 6012 1620 6030
rect 1602 6030 1620 6048
rect 1602 6048 1620 6066
rect 1602 6066 1620 6084
rect 1602 6084 1620 6102
rect 1602 6102 1620 6120
rect 1602 6120 1620 6138
rect 1602 6138 1620 6156
rect 1602 6156 1620 6174
rect 1602 6174 1620 6192
rect 1602 6192 1620 6210
rect 1602 6210 1620 6228
rect 1602 6228 1620 6246
rect 1602 6246 1620 6264
rect 1602 6264 1620 6282
rect 1602 6282 1620 6300
rect 1602 6300 1620 6318
rect 1602 6318 1620 6336
rect 1602 6336 1620 6354
rect 1602 6354 1620 6372
rect 1602 6372 1620 6390
rect 1602 6390 1620 6408
rect 1602 6408 1620 6426
rect 1602 6426 1620 6444
rect 1602 6444 1620 6462
rect 1602 6462 1620 6480
rect 1602 6480 1620 6498
rect 1602 6498 1620 6516
rect 1602 6516 1620 6534
rect 1602 6534 1620 6552
rect 1602 6552 1620 6570
rect 1602 6570 1620 6588
rect 1602 6588 1620 6606
rect 1602 6606 1620 6624
rect 1602 6624 1620 6642
rect 1602 6642 1620 6660
rect 1620 594 1638 612
rect 1620 612 1638 630
rect 1620 630 1638 648
rect 1620 648 1638 666
rect 1620 666 1638 684
rect 1620 684 1638 702
rect 1620 702 1638 720
rect 1620 720 1638 738
rect 1620 738 1638 756
rect 1620 756 1638 774
rect 1620 774 1638 792
rect 1620 792 1638 810
rect 1620 810 1638 828
rect 1620 828 1638 846
rect 1620 846 1638 864
rect 1620 864 1638 882
rect 1620 882 1638 900
rect 1620 900 1638 918
rect 1620 918 1638 936
rect 1620 936 1638 954
rect 1620 954 1638 972
rect 1620 972 1638 990
rect 1620 990 1638 1008
rect 1620 1008 1638 1026
rect 1620 1026 1638 1044
rect 1620 1044 1638 1062
rect 1620 1062 1638 1080
rect 1620 1080 1638 1098
rect 1620 1098 1638 1116
rect 1620 1116 1638 1134
rect 1620 1134 1638 1152
rect 1620 1152 1638 1170
rect 1620 1170 1638 1188
rect 1620 1188 1638 1206
rect 1620 1206 1638 1224
rect 1620 1224 1638 1242
rect 1620 1242 1638 1260
rect 1620 1260 1638 1278
rect 1620 1278 1638 1296
rect 1620 1296 1638 1314
rect 1620 1314 1638 1332
rect 1620 1332 1638 1350
rect 1620 1350 1638 1368
rect 1620 1368 1638 1386
rect 1620 5868 1638 5886
rect 1620 5886 1638 5904
rect 1620 5904 1638 5922
rect 1620 5922 1638 5940
rect 1620 5940 1638 5958
rect 1620 5958 1638 5976
rect 1620 5976 1638 5994
rect 1620 5994 1638 6012
rect 1620 6012 1638 6030
rect 1620 6030 1638 6048
rect 1620 6048 1638 6066
rect 1620 6066 1638 6084
rect 1620 6084 1638 6102
rect 1620 6102 1638 6120
rect 1620 6120 1638 6138
rect 1620 6138 1638 6156
rect 1620 6156 1638 6174
rect 1620 6174 1638 6192
rect 1620 6192 1638 6210
rect 1620 6210 1638 6228
rect 1620 6228 1638 6246
rect 1620 6246 1638 6264
rect 1620 6264 1638 6282
rect 1620 6282 1638 6300
rect 1620 6300 1638 6318
rect 1620 6318 1638 6336
rect 1620 6336 1638 6354
rect 1620 6354 1638 6372
rect 1620 6372 1638 6390
rect 1620 6390 1638 6408
rect 1620 6408 1638 6426
rect 1620 6426 1638 6444
rect 1620 6444 1638 6462
rect 1620 6462 1638 6480
rect 1620 6480 1638 6498
rect 1620 6498 1638 6516
rect 1620 6516 1638 6534
rect 1620 6534 1638 6552
rect 1620 6552 1638 6570
rect 1620 6570 1638 6588
rect 1620 6588 1638 6606
rect 1620 6606 1638 6624
rect 1620 6624 1638 6642
rect 1620 6642 1638 6660
rect 1638 594 1656 612
rect 1638 612 1656 630
rect 1638 630 1656 648
rect 1638 648 1656 666
rect 1638 666 1656 684
rect 1638 684 1656 702
rect 1638 702 1656 720
rect 1638 720 1656 738
rect 1638 738 1656 756
rect 1638 756 1656 774
rect 1638 774 1656 792
rect 1638 792 1656 810
rect 1638 810 1656 828
rect 1638 828 1656 846
rect 1638 846 1656 864
rect 1638 864 1656 882
rect 1638 882 1656 900
rect 1638 900 1656 918
rect 1638 918 1656 936
rect 1638 936 1656 954
rect 1638 954 1656 972
rect 1638 972 1656 990
rect 1638 990 1656 1008
rect 1638 1008 1656 1026
rect 1638 1026 1656 1044
rect 1638 1044 1656 1062
rect 1638 1062 1656 1080
rect 1638 1080 1656 1098
rect 1638 1098 1656 1116
rect 1638 1116 1656 1134
rect 1638 1134 1656 1152
rect 1638 1152 1656 1170
rect 1638 1170 1656 1188
rect 1638 1188 1656 1206
rect 1638 1206 1656 1224
rect 1638 1224 1656 1242
rect 1638 1242 1656 1260
rect 1638 1260 1656 1278
rect 1638 1278 1656 1296
rect 1638 1296 1656 1314
rect 1638 1314 1656 1332
rect 1638 1332 1656 1350
rect 1638 1350 1656 1368
rect 1638 1368 1656 1386
rect 1638 5886 1656 5904
rect 1638 5904 1656 5922
rect 1638 5922 1656 5940
rect 1638 5940 1656 5958
rect 1638 5958 1656 5976
rect 1638 5976 1656 5994
rect 1638 5994 1656 6012
rect 1638 6012 1656 6030
rect 1638 6030 1656 6048
rect 1638 6048 1656 6066
rect 1638 6066 1656 6084
rect 1638 6084 1656 6102
rect 1638 6102 1656 6120
rect 1638 6120 1656 6138
rect 1638 6138 1656 6156
rect 1638 6156 1656 6174
rect 1638 6174 1656 6192
rect 1638 6192 1656 6210
rect 1638 6210 1656 6228
rect 1638 6228 1656 6246
rect 1638 6246 1656 6264
rect 1638 6264 1656 6282
rect 1638 6282 1656 6300
rect 1638 6300 1656 6318
rect 1638 6318 1656 6336
rect 1638 6336 1656 6354
rect 1638 6354 1656 6372
rect 1638 6372 1656 6390
rect 1638 6390 1656 6408
rect 1638 6408 1656 6426
rect 1638 6426 1656 6444
rect 1638 6444 1656 6462
rect 1638 6462 1656 6480
rect 1638 6480 1656 6498
rect 1638 6498 1656 6516
rect 1638 6516 1656 6534
rect 1638 6534 1656 6552
rect 1638 6552 1656 6570
rect 1638 6570 1656 6588
rect 1638 6588 1656 6606
rect 1638 6606 1656 6624
rect 1638 6624 1656 6642
rect 1638 6642 1656 6660
rect 1638 6660 1656 6678
rect 1656 576 1674 594
rect 1656 594 1674 612
rect 1656 612 1674 630
rect 1656 630 1674 648
rect 1656 648 1674 666
rect 1656 666 1674 684
rect 1656 684 1674 702
rect 1656 702 1674 720
rect 1656 720 1674 738
rect 1656 738 1674 756
rect 1656 756 1674 774
rect 1656 774 1674 792
rect 1656 792 1674 810
rect 1656 810 1674 828
rect 1656 828 1674 846
rect 1656 846 1674 864
rect 1656 864 1674 882
rect 1656 882 1674 900
rect 1656 900 1674 918
rect 1656 918 1674 936
rect 1656 936 1674 954
rect 1656 954 1674 972
rect 1656 972 1674 990
rect 1656 990 1674 1008
rect 1656 1008 1674 1026
rect 1656 1026 1674 1044
rect 1656 1044 1674 1062
rect 1656 1062 1674 1080
rect 1656 1080 1674 1098
rect 1656 1098 1674 1116
rect 1656 1116 1674 1134
rect 1656 1134 1674 1152
rect 1656 1152 1674 1170
rect 1656 1170 1674 1188
rect 1656 1188 1674 1206
rect 1656 1206 1674 1224
rect 1656 1224 1674 1242
rect 1656 1242 1674 1260
rect 1656 1260 1674 1278
rect 1656 1278 1674 1296
rect 1656 1296 1674 1314
rect 1656 1314 1674 1332
rect 1656 1332 1674 1350
rect 1656 1350 1674 1368
rect 1656 5904 1674 5922
rect 1656 5922 1674 5940
rect 1656 5940 1674 5958
rect 1656 5958 1674 5976
rect 1656 5976 1674 5994
rect 1656 5994 1674 6012
rect 1656 6012 1674 6030
rect 1656 6030 1674 6048
rect 1656 6048 1674 6066
rect 1656 6066 1674 6084
rect 1656 6084 1674 6102
rect 1656 6102 1674 6120
rect 1656 6120 1674 6138
rect 1656 6138 1674 6156
rect 1656 6156 1674 6174
rect 1656 6174 1674 6192
rect 1656 6192 1674 6210
rect 1656 6210 1674 6228
rect 1656 6228 1674 6246
rect 1656 6246 1674 6264
rect 1656 6264 1674 6282
rect 1656 6282 1674 6300
rect 1656 6300 1674 6318
rect 1656 6318 1674 6336
rect 1656 6336 1674 6354
rect 1656 6354 1674 6372
rect 1656 6372 1674 6390
rect 1656 6390 1674 6408
rect 1656 6408 1674 6426
rect 1656 6426 1674 6444
rect 1656 6444 1674 6462
rect 1656 6462 1674 6480
rect 1656 6480 1674 6498
rect 1656 6498 1674 6516
rect 1656 6516 1674 6534
rect 1656 6534 1674 6552
rect 1656 6552 1674 6570
rect 1656 6570 1674 6588
rect 1656 6588 1674 6606
rect 1656 6606 1674 6624
rect 1656 6624 1674 6642
rect 1656 6642 1674 6660
rect 1656 6660 1674 6678
rect 1656 6678 1674 6696
rect 1674 576 1692 594
rect 1674 594 1692 612
rect 1674 612 1692 630
rect 1674 630 1692 648
rect 1674 648 1692 666
rect 1674 666 1692 684
rect 1674 684 1692 702
rect 1674 702 1692 720
rect 1674 720 1692 738
rect 1674 738 1692 756
rect 1674 756 1692 774
rect 1674 774 1692 792
rect 1674 792 1692 810
rect 1674 810 1692 828
rect 1674 828 1692 846
rect 1674 846 1692 864
rect 1674 864 1692 882
rect 1674 882 1692 900
rect 1674 900 1692 918
rect 1674 918 1692 936
rect 1674 936 1692 954
rect 1674 954 1692 972
rect 1674 972 1692 990
rect 1674 990 1692 1008
rect 1674 1008 1692 1026
rect 1674 1026 1692 1044
rect 1674 1044 1692 1062
rect 1674 1062 1692 1080
rect 1674 1080 1692 1098
rect 1674 1098 1692 1116
rect 1674 1116 1692 1134
rect 1674 1134 1692 1152
rect 1674 1152 1692 1170
rect 1674 1170 1692 1188
rect 1674 1188 1692 1206
rect 1674 1206 1692 1224
rect 1674 1224 1692 1242
rect 1674 1242 1692 1260
rect 1674 1260 1692 1278
rect 1674 1278 1692 1296
rect 1674 1296 1692 1314
rect 1674 1314 1692 1332
rect 1674 1332 1692 1350
rect 1674 5922 1692 5940
rect 1674 5940 1692 5958
rect 1674 5958 1692 5976
rect 1674 5976 1692 5994
rect 1674 5994 1692 6012
rect 1674 6012 1692 6030
rect 1674 6030 1692 6048
rect 1674 6048 1692 6066
rect 1674 6066 1692 6084
rect 1674 6084 1692 6102
rect 1674 6102 1692 6120
rect 1674 6120 1692 6138
rect 1674 6138 1692 6156
rect 1674 6156 1692 6174
rect 1674 6174 1692 6192
rect 1674 6192 1692 6210
rect 1674 6210 1692 6228
rect 1674 6228 1692 6246
rect 1674 6246 1692 6264
rect 1674 6264 1692 6282
rect 1674 6282 1692 6300
rect 1674 6300 1692 6318
rect 1674 6318 1692 6336
rect 1674 6336 1692 6354
rect 1674 6354 1692 6372
rect 1674 6372 1692 6390
rect 1674 6390 1692 6408
rect 1674 6408 1692 6426
rect 1674 6426 1692 6444
rect 1674 6444 1692 6462
rect 1674 6462 1692 6480
rect 1674 6480 1692 6498
rect 1674 6498 1692 6516
rect 1674 6516 1692 6534
rect 1674 6534 1692 6552
rect 1674 6552 1692 6570
rect 1674 6570 1692 6588
rect 1674 6588 1692 6606
rect 1674 6606 1692 6624
rect 1674 6624 1692 6642
rect 1674 6642 1692 6660
rect 1674 6660 1692 6678
rect 1674 6678 1692 6696
rect 1692 558 1710 576
rect 1692 576 1710 594
rect 1692 594 1710 612
rect 1692 612 1710 630
rect 1692 630 1710 648
rect 1692 648 1710 666
rect 1692 666 1710 684
rect 1692 684 1710 702
rect 1692 702 1710 720
rect 1692 720 1710 738
rect 1692 738 1710 756
rect 1692 756 1710 774
rect 1692 774 1710 792
rect 1692 792 1710 810
rect 1692 810 1710 828
rect 1692 828 1710 846
rect 1692 846 1710 864
rect 1692 864 1710 882
rect 1692 882 1710 900
rect 1692 900 1710 918
rect 1692 918 1710 936
rect 1692 936 1710 954
rect 1692 954 1710 972
rect 1692 972 1710 990
rect 1692 990 1710 1008
rect 1692 1008 1710 1026
rect 1692 1026 1710 1044
rect 1692 1044 1710 1062
rect 1692 1062 1710 1080
rect 1692 1080 1710 1098
rect 1692 1098 1710 1116
rect 1692 1116 1710 1134
rect 1692 1134 1710 1152
rect 1692 1152 1710 1170
rect 1692 1170 1710 1188
rect 1692 1188 1710 1206
rect 1692 1206 1710 1224
rect 1692 1224 1710 1242
rect 1692 1242 1710 1260
rect 1692 1260 1710 1278
rect 1692 1278 1710 1296
rect 1692 1296 1710 1314
rect 1692 1314 1710 1332
rect 1692 5940 1710 5958
rect 1692 5958 1710 5976
rect 1692 5976 1710 5994
rect 1692 5994 1710 6012
rect 1692 6012 1710 6030
rect 1692 6030 1710 6048
rect 1692 6048 1710 6066
rect 1692 6066 1710 6084
rect 1692 6084 1710 6102
rect 1692 6102 1710 6120
rect 1692 6120 1710 6138
rect 1692 6138 1710 6156
rect 1692 6156 1710 6174
rect 1692 6174 1710 6192
rect 1692 6192 1710 6210
rect 1692 6210 1710 6228
rect 1692 6228 1710 6246
rect 1692 6246 1710 6264
rect 1692 6264 1710 6282
rect 1692 6282 1710 6300
rect 1692 6300 1710 6318
rect 1692 6318 1710 6336
rect 1692 6336 1710 6354
rect 1692 6354 1710 6372
rect 1692 6372 1710 6390
rect 1692 6390 1710 6408
rect 1692 6408 1710 6426
rect 1692 6426 1710 6444
rect 1692 6444 1710 6462
rect 1692 6462 1710 6480
rect 1692 6480 1710 6498
rect 1692 6498 1710 6516
rect 1692 6516 1710 6534
rect 1692 6534 1710 6552
rect 1692 6552 1710 6570
rect 1692 6570 1710 6588
rect 1692 6588 1710 6606
rect 1692 6606 1710 6624
rect 1692 6624 1710 6642
rect 1692 6642 1710 6660
rect 1692 6660 1710 6678
rect 1692 6678 1710 6696
rect 1692 6696 1710 6714
rect 1710 540 1728 558
rect 1710 558 1728 576
rect 1710 576 1728 594
rect 1710 594 1728 612
rect 1710 612 1728 630
rect 1710 630 1728 648
rect 1710 648 1728 666
rect 1710 666 1728 684
rect 1710 684 1728 702
rect 1710 702 1728 720
rect 1710 720 1728 738
rect 1710 738 1728 756
rect 1710 756 1728 774
rect 1710 774 1728 792
rect 1710 792 1728 810
rect 1710 810 1728 828
rect 1710 828 1728 846
rect 1710 846 1728 864
rect 1710 864 1728 882
rect 1710 882 1728 900
rect 1710 900 1728 918
rect 1710 918 1728 936
rect 1710 936 1728 954
rect 1710 954 1728 972
rect 1710 972 1728 990
rect 1710 990 1728 1008
rect 1710 1008 1728 1026
rect 1710 1026 1728 1044
rect 1710 1044 1728 1062
rect 1710 1062 1728 1080
rect 1710 1080 1728 1098
rect 1710 1098 1728 1116
rect 1710 1116 1728 1134
rect 1710 1134 1728 1152
rect 1710 1152 1728 1170
rect 1710 1170 1728 1188
rect 1710 1188 1728 1206
rect 1710 1206 1728 1224
rect 1710 1224 1728 1242
rect 1710 1242 1728 1260
rect 1710 1260 1728 1278
rect 1710 1278 1728 1296
rect 1710 1296 1728 1314
rect 1710 5958 1728 5976
rect 1710 5976 1728 5994
rect 1710 5994 1728 6012
rect 1710 6012 1728 6030
rect 1710 6030 1728 6048
rect 1710 6048 1728 6066
rect 1710 6066 1728 6084
rect 1710 6084 1728 6102
rect 1710 6102 1728 6120
rect 1710 6120 1728 6138
rect 1710 6138 1728 6156
rect 1710 6156 1728 6174
rect 1710 6174 1728 6192
rect 1710 6192 1728 6210
rect 1710 6210 1728 6228
rect 1710 6228 1728 6246
rect 1710 6246 1728 6264
rect 1710 6264 1728 6282
rect 1710 6282 1728 6300
rect 1710 6300 1728 6318
rect 1710 6318 1728 6336
rect 1710 6336 1728 6354
rect 1710 6354 1728 6372
rect 1710 6372 1728 6390
rect 1710 6390 1728 6408
rect 1710 6408 1728 6426
rect 1710 6426 1728 6444
rect 1710 6444 1728 6462
rect 1710 6462 1728 6480
rect 1710 6480 1728 6498
rect 1710 6498 1728 6516
rect 1710 6516 1728 6534
rect 1710 6534 1728 6552
rect 1710 6552 1728 6570
rect 1710 6570 1728 6588
rect 1710 6588 1728 6606
rect 1710 6606 1728 6624
rect 1710 6624 1728 6642
rect 1710 6642 1728 6660
rect 1710 6660 1728 6678
rect 1710 6678 1728 6696
rect 1710 6696 1728 6714
rect 1728 540 1746 558
rect 1728 558 1746 576
rect 1728 576 1746 594
rect 1728 594 1746 612
rect 1728 612 1746 630
rect 1728 630 1746 648
rect 1728 648 1746 666
rect 1728 666 1746 684
rect 1728 684 1746 702
rect 1728 702 1746 720
rect 1728 720 1746 738
rect 1728 738 1746 756
rect 1728 756 1746 774
rect 1728 774 1746 792
rect 1728 792 1746 810
rect 1728 810 1746 828
rect 1728 828 1746 846
rect 1728 846 1746 864
rect 1728 864 1746 882
rect 1728 882 1746 900
rect 1728 900 1746 918
rect 1728 918 1746 936
rect 1728 936 1746 954
rect 1728 954 1746 972
rect 1728 972 1746 990
rect 1728 990 1746 1008
rect 1728 1008 1746 1026
rect 1728 1026 1746 1044
rect 1728 1044 1746 1062
rect 1728 1062 1746 1080
rect 1728 1080 1746 1098
rect 1728 1098 1746 1116
rect 1728 1116 1746 1134
rect 1728 1134 1746 1152
rect 1728 1152 1746 1170
rect 1728 1170 1746 1188
rect 1728 1188 1746 1206
rect 1728 1206 1746 1224
rect 1728 1224 1746 1242
rect 1728 1242 1746 1260
rect 1728 1260 1746 1278
rect 1728 1278 1746 1296
rect 1728 5976 1746 5994
rect 1728 5994 1746 6012
rect 1728 6012 1746 6030
rect 1728 6030 1746 6048
rect 1728 6048 1746 6066
rect 1728 6066 1746 6084
rect 1728 6084 1746 6102
rect 1728 6102 1746 6120
rect 1728 6120 1746 6138
rect 1728 6138 1746 6156
rect 1728 6156 1746 6174
rect 1728 6174 1746 6192
rect 1728 6192 1746 6210
rect 1728 6210 1746 6228
rect 1728 6228 1746 6246
rect 1728 6246 1746 6264
rect 1728 6264 1746 6282
rect 1728 6282 1746 6300
rect 1728 6300 1746 6318
rect 1728 6318 1746 6336
rect 1728 6336 1746 6354
rect 1728 6354 1746 6372
rect 1728 6372 1746 6390
rect 1728 6390 1746 6408
rect 1728 6408 1746 6426
rect 1728 6426 1746 6444
rect 1728 6444 1746 6462
rect 1728 6462 1746 6480
rect 1728 6480 1746 6498
rect 1728 6498 1746 6516
rect 1728 6516 1746 6534
rect 1728 6534 1746 6552
rect 1728 6552 1746 6570
rect 1728 6570 1746 6588
rect 1728 6588 1746 6606
rect 1728 6606 1746 6624
rect 1728 6624 1746 6642
rect 1728 6642 1746 6660
rect 1728 6660 1746 6678
rect 1728 6678 1746 6696
rect 1728 6696 1746 6714
rect 1728 6714 1746 6732
rect 1746 522 1764 540
rect 1746 540 1764 558
rect 1746 558 1764 576
rect 1746 576 1764 594
rect 1746 594 1764 612
rect 1746 612 1764 630
rect 1746 630 1764 648
rect 1746 648 1764 666
rect 1746 666 1764 684
rect 1746 684 1764 702
rect 1746 702 1764 720
rect 1746 720 1764 738
rect 1746 738 1764 756
rect 1746 756 1764 774
rect 1746 774 1764 792
rect 1746 792 1764 810
rect 1746 810 1764 828
rect 1746 828 1764 846
rect 1746 846 1764 864
rect 1746 864 1764 882
rect 1746 882 1764 900
rect 1746 900 1764 918
rect 1746 918 1764 936
rect 1746 936 1764 954
rect 1746 954 1764 972
rect 1746 972 1764 990
rect 1746 990 1764 1008
rect 1746 1008 1764 1026
rect 1746 1026 1764 1044
rect 1746 1044 1764 1062
rect 1746 1062 1764 1080
rect 1746 1080 1764 1098
rect 1746 1098 1764 1116
rect 1746 1116 1764 1134
rect 1746 1134 1764 1152
rect 1746 1152 1764 1170
rect 1746 1170 1764 1188
rect 1746 1188 1764 1206
rect 1746 1206 1764 1224
rect 1746 1224 1764 1242
rect 1746 1242 1764 1260
rect 1746 1260 1764 1278
rect 1746 5976 1764 5994
rect 1746 5994 1764 6012
rect 1746 6012 1764 6030
rect 1746 6030 1764 6048
rect 1746 6048 1764 6066
rect 1746 6066 1764 6084
rect 1746 6084 1764 6102
rect 1746 6102 1764 6120
rect 1746 6120 1764 6138
rect 1746 6138 1764 6156
rect 1746 6156 1764 6174
rect 1746 6174 1764 6192
rect 1746 6192 1764 6210
rect 1746 6210 1764 6228
rect 1746 6228 1764 6246
rect 1746 6246 1764 6264
rect 1746 6264 1764 6282
rect 1746 6282 1764 6300
rect 1746 6300 1764 6318
rect 1746 6318 1764 6336
rect 1746 6336 1764 6354
rect 1746 6354 1764 6372
rect 1746 6372 1764 6390
rect 1746 6390 1764 6408
rect 1746 6408 1764 6426
rect 1746 6426 1764 6444
rect 1746 6444 1764 6462
rect 1746 6462 1764 6480
rect 1746 6480 1764 6498
rect 1746 6498 1764 6516
rect 1746 6516 1764 6534
rect 1746 6534 1764 6552
rect 1746 6552 1764 6570
rect 1746 6570 1764 6588
rect 1746 6588 1764 6606
rect 1746 6606 1764 6624
rect 1746 6624 1764 6642
rect 1746 6642 1764 6660
rect 1746 6660 1764 6678
rect 1746 6678 1764 6696
rect 1746 6696 1764 6714
rect 1746 6714 1764 6732
rect 1746 6732 1764 6750
rect 1764 504 1782 522
rect 1764 522 1782 540
rect 1764 540 1782 558
rect 1764 558 1782 576
rect 1764 576 1782 594
rect 1764 594 1782 612
rect 1764 612 1782 630
rect 1764 630 1782 648
rect 1764 648 1782 666
rect 1764 666 1782 684
rect 1764 684 1782 702
rect 1764 702 1782 720
rect 1764 720 1782 738
rect 1764 738 1782 756
rect 1764 756 1782 774
rect 1764 774 1782 792
rect 1764 792 1782 810
rect 1764 810 1782 828
rect 1764 828 1782 846
rect 1764 846 1782 864
rect 1764 864 1782 882
rect 1764 882 1782 900
rect 1764 900 1782 918
rect 1764 918 1782 936
rect 1764 936 1782 954
rect 1764 954 1782 972
rect 1764 972 1782 990
rect 1764 990 1782 1008
rect 1764 1008 1782 1026
rect 1764 1026 1782 1044
rect 1764 1044 1782 1062
rect 1764 1062 1782 1080
rect 1764 1080 1782 1098
rect 1764 1098 1782 1116
rect 1764 1116 1782 1134
rect 1764 1134 1782 1152
rect 1764 1152 1782 1170
rect 1764 1170 1782 1188
rect 1764 1188 1782 1206
rect 1764 1206 1782 1224
rect 1764 1224 1782 1242
rect 1764 1242 1782 1260
rect 1764 1260 1782 1278
rect 1764 5994 1782 6012
rect 1764 6012 1782 6030
rect 1764 6030 1782 6048
rect 1764 6048 1782 6066
rect 1764 6066 1782 6084
rect 1764 6084 1782 6102
rect 1764 6102 1782 6120
rect 1764 6120 1782 6138
rect 1764 6138 1782 6156
rect 1764 6156 1782 6174
rect 1764 6174 1782 6192
rect 1764 6192 1782 6210
rect 1764 6210 1782 6228
rect 1764 6228 1782 6246
rect 1764 6246 1782 6264
rect 1764 6264 1782 6282
rect 1764 6282 1782 6300
rect 1764 6300 1782 6318
rect 1764 6318 1782 6336
rect 1764 6336 1782 6354
rect 1764 6354 1782 6372
rect 1764 6372 1782 6390
rect 1764 6390 1782 6408
rect 1764 6408 1782 6426
rect 1764 6426 1782 6444
rect 1764 6444 1782 6462
rect 1764 6462 1782 6480
rect 1764 6480 1782 6498
rect 1764 6498 1782 6516
rect 1764 6516 1782 6534
rect 1764 6534 1782 6552
rect 1764 6552 1782 6570
rect 1764 6570 1782 6588
rect 1764 6588 1782 6606
rect 1764 6606 1782 6624
rect 1764 6624 1782 6642
rect 1764 6642 1782 6660
rect 1764 6660 1782 6678
rect 1764 6678 1782 6696
rect 1764 6696 1782 6714
rect 1764 6714 1782 6732
rect 1764 6732 1782 6750
rect 1782 504 1800 522
rect 1782 522 1800 540
rect 1782 540 1800 558
rect 1782 558 1800 576
rect 1782 576 1800 594
rect 1782 594 1800 612
rect 1782 612 1800 630
rect 1782 630 1800 648
rect 1782 648 1800 666
rect 1782 666 1800 684
rect 1782 684 1800 702
rect 1782 702 1800 720
rect 1782 720 1800 738
rect 1782 738 1800 756
rect 1782 756 1800 774
rect 1782 774 1800 792
rect 1782 792 1800 810
rect 1782 810 1800 828
rect 1782 828 1800 846
rect 1782 846 1800 864
rect 1782 864 1800 882
rect 1782 882 1800 900
rect 1782 900 1800 918
rect 1782 918 1800 936
rect 1782 936 1800 954
rect 1782 954 1800 972
rect 1782 972 1800 990
rect 1782 990 1800 1008
rect 1782 1008 1800 1026
rect 1782 1026 1800 1044
rect 1782 1044 1800 1062
rect 1782 1062 1800 1080
rect 1782 1080 1800 1098
rect 1782 1098 1800 1116
rect 1782 1116 1800 1134
rect 1782 1134 1800 1152
rect 1782 1152 1800 1170
rect 1782 1170 1800 1188
rect 1782 1188 1800 1206
rect 1782 1206 1800 1224
rect 1782 1224 1800 1242
rect 1782 1242 1800 1260
rect 1782 6012 1800 6030
rect 1782 6030 1800 6048
rect 1782 6048 1800 6066
rect 1782 6066 1800 6084
rect 1782 6084 1800 6102
rect 1782 6102 1800 6120
rect 1782 6120 1800 6138
rect 1782 6138 1800 6156
rect 1782 6156 1800 6174
rect 1782 6174 1800 6192
rect 1782 6192 1800 6210
rect 1782 6210 1800 6228
rect 1782 6228 1800 6246
rect 1782 6246 1800 6264
rect 1782 6264 1800 6282
rect 1782 6282 1800 6300
rect 1782 6300 1800 6318
rect 1782 6318 1800 6336
rect 1782 6336 1800 6354
rect 1782 6354 1800 6372
rect 1782 6372 1800 6390
rect 1782 6390 1800 6408
rect 1782 6408 1800 6426
rect 1782 6426 1800 6444
rect 1782 6444 1800 6462
rect 1782 6462 1800 6480
rect 1782 6480 1800 6498
rect 1782 6498 1800 6516
rect 1782 6516 1800 6534
rect 1782 6534 1800 6552
rect 1782 6552 1800 6570
rect 1782 6570 1800 6588
rect 1782 6588 1800 6606
rect 1782 6606 1800 6624
rect 1782 6624 1800 6642
rect 1782 6642 1800 6660
rect 1782 6660 1800 6678
rect 1782 6678 1800 6696
rect 1782 6696 1800 6714
rect 1782 6714 1800 6732
rect 1782 6732 1800 6750
rect 1782 6750 1800 6768
rect 1800 486 1818 504
rect 1800 504 1818 522
rect 1800 522 1818 540
rect 1800 540 1818 558
rect 1800 558 1818 576
rect 1800 576 1818 594
rect 1800 594 1818 612
rect 1800 612 1818 630
rect 1800 630 1818 648
rect 1800 648 1818 666
rect 1800 666 1818 684
rect 1800 684 1818 702
rect 1800 702 1818 720
rect 1800 720 1818 738
rect 1800 738 1818 756
rect 1800 756 1818 774
rect 1800 774 1818 792
rect 1800 792 1818 810
rect 1800 810 1818 828
rect 1800 828 1818 846
rect 1800 846 1818 864
rect 1800 864 1818 882
rect 1800 882 1818 900
rect 1800 900 1818 918
rect 1800 918 1818 936
rect 1800 936 1818 954
rect 1800 954 1818 972
rect 1800 972 1818 990
rect 1800 990 1818 1008
rect 1800 1008 1818 1026
rect 1800 1026 1818 1044
rect 1800 1044 1818 1062
rect 1800 1062 1818 1080
rect 1800 1080 1818 1098
rect 1800 1098 1818 1116
rect 1800 1116 1818 1134
rect 1800 1134 1818 1152
rect 1800 1152 1818 1170
rect 1800 1170 1818 1188
rect 1800 1188 1818 1206
rect 1800 1206 1818 1224
rect 1800 1224 1818 1242
rect 1800 6030 1818 6048
rect 1800 6048 1818 6066
rect 1800 6066 1818 6084
rect 1800 6084 1818 6102
rect 1800 6102 1818 6120
rect 1800 6120 1818 6138
rect 1800 6138 1818 6156
rect 1800 6156 1818 6174
rect 1800 6174 1818 6192
rect 1800 6192 1818 6210
rect 1800 6210 1818 6228
rect 1800 6228 1818 6246
rect 1800 6246 1818 6264
rect 1800 6264 1818 6282
rect 1800 6282 1818 6300
rect 1800 6300 1818 6318
rect 1800 6318 1818 6336
rect 1800 6336 1818 6354
rect 1800 6354 1818 6372
rect 1800 6372 1818 6390
rect 1800 6390 1818 6408
rect 1800 6408 1818 6426
rect 1800 6426 1818 6444
rect 1800 6444 1818 6462
rect 1800 6462 1818 6480
rect 1800 6480 1818 6498
rect 1800 6498 1818 6516
rect 1800 6516 1818 6534
rect 1800 6534 1818 6552
rect 1800 6552 1818 6570
rect 1800 6570 1818 6588
rect 1800 6588 1818 6606
rect 1800 6606 1818 6624
rect 1800 6624 1818 6642
rect 1800 6642 1818 6660
rect 1800 6660 1818 6678
rect 1800 6678 1818 6696
rect 1800 6696 1818 6714
rect 1800 6714 1818 6732
rect 1800 6732 1818 6750
rect 1800 6750 1818 6768
rect 1800 6768 1818 6786
rect 1818 486 1836 504
rect 1818 504 1836 522
rect 1818 522 1836 540
rect 1818 540 1836 558
rect 1818 558 1836 576
rect 1818 576 1836 594
rect 1818 594 1836 612
rect 1818 612 1836 630
rect 1818 630 1836 648
rect 1818 648 1836 666
rect 1818 666 1836 684
rect 1818 684 1836 702
rect 1818 702 1836 720
rect 1818 720 1836 738
rect 1818 738 1836 756
rect 1818 756 1836 774
rect 1818 774 1836 792
rect 1818 792 1836 810
rect 1818 810 1836 828
rect 1818 828 1836 846
rect 1818 846 1836 864
rect 1818 864 1836 882
rect 1818 882 1836 900
rect 1818 900 1836 918
rect 1818 918 1836 936
rect 1818 936 1836 954
rect 1818 954 1836 972
rect 1818 972 1836 990
rect 1818 990 1836 1008
rect 1818 1008 1836 1026
rect 1818 1026 1836 1044
rect 1818 1044 1836 1062
rect 1818 1062 1836 1080
rect 1818 1080 1836 1098
rect 1818 1098 1836 1116
rect 1818 1116 1836 1134
rect 1818 1134 1836 1152
rect 1818 1152 1836 1170
rect 1818 1170 1836 1188
rect 1818 1188 1836 1206
rect 1818 1206 1836 1224
rect 1818 6048 1836 6066
rect 1818 6066 1836 6084
rect 1818 6084 1836 6102
rect 1818 6102 1836 6120
rect 1818 6120 1836 6138
rect 1818 6138 1836 6156
rect 1818 6156 1836 6174
rect 1818 6174 1836 6192
rect 1818 6192 1836 6210
rect 1818 6210 1836 6228
rect 1818 6228 1836 6246
rect 1818 6246 1836 6264
rect 1818 6264 1836 6282
rect 1818 6282 1836 6300
rect 1818 6300 1836 6318
rect 1818 6318 1836 6336
rect 1818 6336 1836 6354
rect 1818 6354 1836 6372
rect 1818 6372 1836 6390
rect 1818 6390 1836 6408
rect 1818 6408 1836 6426
rect 1818 6426 1836 6444
rect 1818 6444 1836 6462
rect 1818 6462 1836 6480
rect 1818 6480 1836 6498
rect 1818 6498 1836 6516
rect 1818 6516 1836 6534
rect 1818 6534 1836 6552
rect 1818 6552 1836 6570
rect 1818 6570 1836 6588
rect 1818 6588 1836 6606
rect 1818 6606 1836 6624
rect 1818 6624 1836 6642
rect 1818 6642 1836 6660
rect 1818 6660 1836 6678
rect 1818 6678 1836 6696
rect 1818 6696 1836 6714
rect 1818 6714 1836 6732
rect 1818 6732 1836 6750
rect 1818 6750 1836 6768
rect 1818 6768 1836 6786
rect 1836 468 1854 486
rect 1836 486 1854 504
rect 1836 504 1854 522
rect 1836 522 1854 540
rect 1836 540 1854 558
rect 1836 558 1854 576
rect 1836 576 1854 594
rect 1836 594 1854 612
rect 1836 612 1854 630
rect 1836 630 1854 648
rect 1836 648 1854 666
rect 1836 666 1854 684
rect 1836 684 1854 702
rect 1836 702 1854 720
rect 1836 720 1854 738
rect 1836 738 1854 756
rect 1836 756 1854 774
rect 1836 774 1854 792
rect 1836 792 1854 810
rect 1836 810 1854 828
rect 1836 828 1854 846
rect 1836 846 1854 864
rect 1836 864 1854 882
rect 1836 882 1854 900
rect 1836 900 1854 918
rect 1836 918 1854 936
rect 1836 936 1854 954
rect 1836 954 1854 972
rect 1836 972 1854 990
rect 1836 990 1854 1008
rect 1836 1008 1854 1026
rect 1836 1026 1854 1044
rect 1836 1044 1854 1062
rect 1836 1062 1854 1080
rect 1836 1080 1854 1098
rect 1836 1098 1854 1116
rect 1836 1116 1854 1134
rect 1836 1134 1854 1152
rect 1836 1152 1854 1170
rect 1836 1170 1854 1188
rect 1836 1188 1854 1206
rect 1836 6048 1854 6066
rect 1836 6066 1854 6084
rect 1836 6084 1854 6102
rect 1836 6102 1854 6120
rect 1836 6120 1854 6138
rect 1836 6138 1854 6156
rect 1836 6156 1854 6174
rect 1836 6174 1854 6192
rect 1836 6192 1854 6210
rect 1836 6210 1854 6228
rect 1836 6228 1854 6246
rect 1836 6246 1854 6264
rect 1836 6264 1854 6282
rect 1836 6282 1854 6300
rect 1836 6300 1854 6318
rect 1836 6318 1854 6336
rect 1836 6336 1854 6354
rect 1836 6354 1854 6372
rect 1836 6372 1854 6390
rect 1836 6390 1854 6408
rect 1836 6408 1854 6426
rect 1836 6426 1854 6444
rect 1836 6444 1854 6462
rect 1836 6462 1854 6480
rect 1836 6480 1854 6498
rect 1836 6498 1854 6516
rect 1836 6516 1854 6534
rect 1836 6534 1854 6552
rect 1836 6552 1854 6570
rect 1836 6570 1854 6588
rect 1836 6588 1854 6606
rect 1836 6606 1854 6624
rect 1836 6624 1854 6642
rect 1836 6642 1854 6660
rect 1836 6660 1854 6678
rect 1836 6678 1854 6696
rect 1836 6696 1854 6714
rect 1836 6714 1854 6732
rect 1836 6732 1854 6750
rect 1836 6750 1854 6768
rect 1836 6768 1854 6786
rect 1836 6786 1854 6804
rect 1854 450 1872 468
rect 1854 468 1872 486
rect 1854 486 1872 504
rect 1854 504 1872 522
rect 1854 522 1872 540
rect 1854 540 1872 558
rect 1854 558 1872 576
rect 1854 576 1872 594
rect 1854 594 1872 612
rect 1854 612 1872 630
rect 1854 630 1872 648
rect 1854 648 1872 666
rect 1854 666 1872 684
rect 1854 684 1872 702
rect 1854 702 1872 720
rect 1854 720 1872 738
rect 1854 738 1872 756
rect 1854 756 1872 774
rect 1854 774 1872 792
rect 1854 792 1872 810
rect 1854 810 1872 828
rect 1854 828 1872 846
rect 1854 846 1872 864
rect 1854 864 1872 882
rect 1854 882 1872 900
rect 1854 900 1872 918
rect 1854 918 1872 936
rect 1854 936 1872 954
rect 1854 954 1872 972
rect 1854 972 1872 990
rect 1854 990 1872 1008
rect 1854 1008 1872 1026
rect 1854 1026 1872 1044
rect 1854 1044 1872 1062
rect 1854 1062 1872 1080
rect 1854 1080 1872 1098
rect 1854 1098 1872 1116
rect 1854 1116 1872 1134
rect 1854 1134 1872 1152
rect 1854 1152 1872 1170
rect 1854 1170 1872 1188
rect 1854 1188 1872 1206
rect 1854 6066 1872 6084
rect 1854 6084 1872 6102
rect 1854 6102 1872 6120
rect 1854 6120 1872 6138
rect 1854 6138 1872 6156
rect 1854 6156 1872 6174
rect 1854 6174 1872 6192
rect 1854 6192 1872 6210
rect 1854 6210 1872 6228
rect 1854 6228 1872 6246
rect 1854 6246 1872 6264
rect 1854 6264 1872 6282
rect 1854 6282 1872 6300
rect 1854 6300 1872 6318
rect 1854 6318 1872 6336
rect 1854 6336 1872 6354
rect 1854 6354 1872 6372
rect 1854 6372 1872 6390
rect 1854 6390 1872 6408
rect 1854 6408 1872 6426
rect 1854 6426 1872 6444
rect 1854 6444 1872 6462
rect 1854 6462 1872 6480
rect 1854 6480 1872 6498
rect 1854 6498 1872 6516
rect 1854 6516 1872 6534
rect 1854 6534 1872 6552
rect 1854 6552 1872 6570
rect 1854 6570 1872 6588
rect 1854 6588 1872 6606
rect 1854 6606 1872 6624
rect 1854 6624 1872 6642
rect 1854 6642 1872 6660
rect 1854 6660 1872 6678
rect 1854 6678 1872 6696
rect 1854 6696 1872 6714
rect 1854 6714 1872 6732
rect 1854 6732 1872 6750
rect 1854 6750 1872 6768
rect 1854 6768 1872 6786
rect 1854 6786 1872 6804
rect 1872 450 1890 468
rect 1872 468 1890 486
rect 1872 486 1890 504
rect 1872 504 1890 522
rect 1872 522 1890 540
rect 1872 540 1890 558
rect 1872 558 1890 576
rect 1872 576 1890 594
rect 1872 594 1890 612
rect 1872 612 1890 630
rect 1872 630 1890 648
rect 1872 648 1890 666
rect 1872 666 1890 684
rect 1872 684 1890 702
rect 1872 702 1890 720
rect 1872 720 1890 738
rect 1872 738 1890 756
rect 1872 756 1890 774
rect 1872 774 1890 792
rect 1872 792 1890 810
rect 1872 810 1890 828
rect 1872 828 1890 846
rect 1872 846 1890 864
rect 1872 864 1890 882
rect 1872 882 1890 900
rect 1872 900 1890 918
rect 1872 918 1890 936
rect 1872 936 1890 954
rect 1872 954 1890 972
rect 1872 972 1890 990
rect 1872 990 1890 1008
rect 1872 1008 1890 1026
rect 1872 1026 1890 1044
rect 1872 1044 1890 1062
rect 1872 1062 1890 1080
rect 1872 1080 1890 1098
rect 1872 1098 1890 1116
rect 1872 1116 1890 1134
rect 1872 1134 1890 1152
rect 1872 1152 1890 1170
rect 1872 1170 1890 1188
rect 1872 6084 1890 6102
rect 1872 6102 1890 6120
rect 1872 6120 1890 6138
rect 1872 6138 1890 6156
rect 1872 6156 1890 6174
rect 1872 6174 1890 6192
rect 1872 6192 1890 6210
rect 1872 6210 1890 6228
rect 1872 6228 1890 6246
rect 1872 6246 1890 6264
rect 1872 6264 1890 6282
rect 1872 6282 1890 6300
rect 1872 6300 1890 6318
rect 1872 6318 1890 6336
rect 1872 6336 1890 6354
rect 1872 6354 1890 6372
rect 1872 6372 1890 6390
rect 1872 6390 1890 6408
rect 1872 6408 1890 6426
rect 1872 6426 1890 6444
rect 1872 6444 1890 6462
rect 1872 6462 1890 6480
rect 1872 6480 1890 6498
rect 1872 6498 1890 6516
rect 1872 6516 1890 6534
rect 1872 6534 1890 6552
rect 1872 6552 1890 6570
rect 1872 6570 1890 6588
rect 1872 6588 1890 6606
rect 1872 6606 1890 6624
rect 1872 6624 1890 6642
rect 1872 6642 1890 6660
rect 1872 6660 1890 6678
rect 1872 6678 1890 6696
rect 1872 6696 1890 6714
rect 1872 6714 1890 6732
rect 1872 6732 1890 6750
rect 1872 6750 1890 6768
rect 1872 6768 1890 6786
rect 1872 6786 1890 6804
rect 1872 6804 1890 6822
rect 1890 432 1908 450
rect 1890 450 1908 468
rect 1890 468 1908 486
rect 1890 486 1908 504
rect 1890 504 1908 522
rect 1890 522 1908 540
rect 1890 540 1908 558
rect 1890 558 1908 576
rect 1890 576 1908 594
rect 1890 594 1908 612
rect 1890 612 1908 630
rect 1890 630 1908 648
rect 1890 648 1908 666
rect 1890 666 1908 684
rect 1890 684 1908 702
rect 1890 702 1908 720
rect 1890 720 1908 738
rect 1890 738 1908 756
rect 1890 756 1908 774
rect 1890 774 1908 792
rect 1890 792 1908 810
rect 1890 810 1908 828
rect 1890 828 1908 846
rect 1890 846 1908 864
rect 1890 864 1908 882
rect 1890 882 1908 900
rect 1890 900 1908 918
rect 1890 918 1908 936
rect 1890 936 1908 954
rect 1890 954 1908 972
rect 1890 972 1908 990
rect 1890 990 1908 1008
rect 1890 1008 1908 1026
rect 1890 1026 1908 1044
rect 1890 1044 1908 1062
rect 1890 1062 1908 1080
rect 1890 1080 1908 1098
rect 1890 1098 1908 1116
rect 1890 1116 1908 1134
rect 1890 1134 1908 1152
rect 1890 1152 1908 1170
rect 1890 6084 1908 6102
rect 1890 6102 1908 6120
rect 1890 6120 1908 6138
rect 1890 6138 1908 6156
rect 1890 6156 1908 6174
rect 1890 6174 1908 6192
rect 1890 6192 1908 6210
rect 1890 6210 1908 6228
rect 1890 6228 1908 6246
rect 1890 6246 1908 6264
rect 1890 6264 1908 6282
rect 1890 6282 1908 6300
rect 1890 6300 1908 6318
rect 1890 6318 1908 6336
rect 1890 6336 1908 6354
rect 1890 6354 1908 6372
rect 1890 6372 1908 6390
rect 1890 6390 1908 6408
rect 1890 6408 1908 6426
rect 1890 6426 1908 6444
rect 1890 6444 1908 6462
rect 1890 6462 1908 6480
rect 1890 6480 1908 6498
rect 1890 6498 1908 6516
rect 1890 6516 1908 6534
rect 1890 6534 1908 6552
rect 1890 6552 1908 6570
rect 1890 6570 1908 6588
rect 1890 6588 1908 6606
rect 1890 6606 1908 6624
rect 1890 6624 1908 6642
rect 1890 6642 1908 6660
rect 1890 6660 1908 6678
rect 1890 6678 1908 6696
rect 1890 6696 1908 6714
rect 1890 6714 1908 6732
rect 1890 6732 1908 6750
rect 1890 6750 1908 6768
rect 1890 6768 1908 6786
rect 1890 6786 1908 6804
rect 1890 6804 1908 6822
rect 1908 432 1926 450
rect 1908 450 1926 468
rect 1908 468 1926 486
rect 1908 486 1926 504
rect 1908 504 1926 522
rect 1908 522 1926 540
rect 1908 540 1926 558
rect 1908 558 1926 576
rect 1908 576 1926 594
rect 1908 594 1926 612
rect 1908 612 1926 630
rect 1908 630 1926 648
rect 1908 648 1926 666
rect 1908 666 1926 684
rect 1908 684 1926 702
rect 1908 702 1926 720
rect 1908 720 1926 738
rect 1908 738 1926 756
rect 1908 756 1926 774
rect 1908 774 1926 792
rect 1908 792 1926 810
rect 1908 810 1926 828
rect 1908 828 1926 846
rect 1908 846 1926 864
rect 1908 864 1926 882
rect 1908 882 1926 900
rect 1908 900 1926 918
rect 1908 918 1926 936
rect 1908 936 1926 954
rect 1908 954 1926 972
rect 1908 972 1926 990
rect 1908 990 1926 1008
rect 1908 1008 1926 1026
rect 1908 1026 1926 1044
rect 1908 1044 1926 1062
rect 1908 1062 1926 1080
rect 1908 1080 1926 1098
rect 1908 1098 1926 1116
rect 1908 1116 1926 1134
rect 1908 1134 1926 1152
rect 1908 6102 1926 6120
rect 1908 6120 1926 6138
rect 1908 6138 1926 6156
rect 1908 6156 1926 6174
rect 1908 6174 1926 6192
rect 1908 6192 1926 6210
rect 1908 6210 1926 6228
rect 1908 6228 1926 6246
rect 1908 6246 1926 6264
rect 1908 6264 1926 6282
rect 1908 6282 1926 6300
rect 1908 6300 1926 6318
rect 1908 6318 1926 6336
rect 1908 6336 1926 6354
rect 1908 6354 1926 6372
rect 1908 6372 1926 6390
rect 1908 6390 1926 6408
rect 1908 6408 1926 6426
rect 1908 6426 1926 6444
rect 1908 6444 1926 6462
rect 1908 6462 1926 6480
rect 1908 6480 1926 6498
rect 1908 6498 1926 6516
rect 1908 6516 1926 6534
rect 1908 6534 1926 6552
rect 1908 6552 1926 6570
rect 1908 6570 1926 6588
rect 1908 6588 1926 6606
rect 1908 6606 1926 6624
rect 1908 6624 1926 6642
rect 1908 6642 1926 6660
rect 1908 6660 1926 6678
rect 1908 6678 1926 6696
rect 1908 6696 1926 6714
rect 1908 6714 1926 6732
rect 1908 6732 1926 6750
rect 1908 6750 1926 6768
rect 1908 6768 1926 6786
rect 1908 6786 1926 6804
rect 1908 6804 1926 6822
rect 1908 6822 1926 6840
rect 1926 414 1944 432
rect 1926 432 1944 450
rect 1926 450 1944 468
rect 1926 468 1944 486
rect 1926 486 1944 504
rect 1926 504 1944 522
rect 1926 522 1944 540
rect 1926 540 1944 558
rect 1926 558 1944 576
rect 1926 576 1944 594
rect 1926 594 1944 612
rect 1926 612 1944 630
rect 1926 630 1944 648
rect 1926 648 1944 666
rect 1926 666 1944 684
rect 1926 684 1944 702
rect 1926 702 1944 720
rect 1926 720 1944 738
rect 1926 738 1944 756
rect 1926 756 1944 774
rect 1926 774 1944 792
rect 1926 792 1944 810
rect 1926 810 1944 828
rect 1926 828 1944 846
rect 1926 846 1944 864
rect 1926 864 1944 882
rect 1926 882 1944 900
rect 1926 900 1944 918
rect 1926 918 1944 936
rect 1926 936 1944 954
rect 1926 954 1944 972
rect 1926 972 1944 990
rect 1926 990 1944 1008
rect 1926 1008 1944 1026
rect 1926 1026 1944 1044
rect 1926 1044 1944 1062
rect 1926 1062 1944 1080
rect 1926 1080 1944 1098
rect 1926 1098 1944 1116
rect 1926 1116 1944 1134
rect 1926 1134 1944 1152
rect 1926 6120 1944 6138
rect 1926 6138 1944 6156
rect 1926 6156 1944 6174
rect 1926 6174 1944 6192
rect 1926 6192 1944 6210
rect 1926 6210 1944 6228
rect 1926 6228 1944 6246
rect 1926 6246 1944 6264
rect 1926 6264 1944 6282
rect 1926 6282 1944 6300
rect 1926 6300 1944 6318
rect 1926 6318 1944 6336
rect 1926 6336 1944 6354
rect 1926 6354 1944 6372
rect 1926 6372 1944 6390
rect 1926 6390 1944 6408
rect 1926 6408 1944 6426
rect 1926 6426 1944 6444
rect 1926 6444 1944 6462
rect 1926 6462 1944 6480
rect 1926 6480 1944 6498
rect 1926 6498 1944 6516
rect 1926 6516 1944 6534
rect 1926 6534 1944 6552
rect 1926 6552 1944 6570
rect 1926 6570 1944 6588
rect 1926 6588 1944 6606
rect 1926 6606 1944 6624
rect 1926 6624 1944 6642
rect 1926 6642 1944 6660
rect 1926 6660 1944 6678
rect 1926 6678 1944 6696
rect 1926 6696 1944 6714
rect 1926 6714 1944 6732
rect 1926 6732 1944 6750
rect 1926 6750 1944 6768
rect 1926 6768 1944 6786
rect 1926 6786 1944 6804
rect 1926 6804 1944 6822
rect 1926 6822 1944 6840
rect 1944 414 1962 432
rect 1944 432 1962 450
rect 1944 450 1962 468
rect 1944 468 1962 486
rect 1944 486 1962 504
rect 1944 504 1962 522
rect 1944 522 1962 540
rect 1944 540 1962 558
rect 1944 558 1962 576
rect 1944 576 1962 594
rect 1944 594 1962 612
rect 1944 612 1962 630
rect 1944 630 1962 648
rect 1944 648 1962 666
rect 1944 666 1962 684
rect 1944 684 1962 702
rect 1944 702 1962 720
rect 1944 720 1962 738
rect 1944 738 1962 756
rect 1944 756 1962 774
rect 1944 774 1962 792
rect 1944 792 1962 810
rect 1944 810 1962 828
rect 1944 828 1962 846
rect 1944 846 1962 864
rect 1944 864 1962 882
rect 1944 882 1962 900
rect 1944 900 1962 918
rect 1944 918 1962 936
rect 1944 936 1962 954
rect 1944 954 1962 972
rect 1944 972 1962 990
rect 1944 990 1962 1008
rect 1944 1008 1962 1026
rect 1944 1026 1962 1044
rect 1944 1044 1962 1062
rect 1944 1062 1962 1080
rect 1944 1080 1962 1098
rect 1944 1098 1962 1116
rect 1944 1116 1962 1134
rect 1944 6138 1962 6156
rect 1944 6156 1962 6174
rect 1944 6174 1962 6192
rect 1944 6192 1962 6210
rect 1944 6210 1962 6228
rect 1944 6228 1962 6246
rect 1944 6246 1962 6264
rect 1944 6264 1962 6282
rect 1944 6282 1962 6300
rect 1944 6300 1962 6318
rect 1944 6318 1962 6336
rect 1944 6336 1962 6354
rect 1944 6354 1962 6372
rect 1944 6372 1962 6390
rect 1944 6390 1962 6408
rect 1944 6408 1962 6426
rect 1944 6426 1962 6444
rect 1944 6444 1962 6462
rect 1944 6462 1962 6480
rect 1944 6480 1962 6498
rect 1944 6498 1962 6516
rect 1944 6516 1962 6534
rect 1944 6534 1962 6552
rect 1944 6552 1962 6570
rect 1944 6570 1962 6588
rect 1944 6588 1962 6606
rect 1944 6606 1962 6624
rect 1944 6624 1962 6642
rect 1944 6642 1962 6660
rect 1944 6660 1962 6678
rect 1944 6678 1962 6696
rect 1944 6696 1962 6714
rect 1944 6714 1962 6732
rect 1944 6732 1962 6750
rect 1944 6750 1962 6768
rect 1944 6768 1962 6786
rect 1944 6786 1962 6804
rect 1944 6804 1962 6822
rect 1944 6822 1962 6840
rect 1944 6840 1962 6858
rect 1962 396 1980 414
rect 1962 414 1980 432
rect 1962 432 1980 450
rect 1962 450 1980 468
rect 1962 468 1980 486
rect 1962 486 1980 504
rect 1962 504 1980 522
rect 1962 522 1980 540
rect 1962 540 1980 558
rect 1962 558 1980 576
rect 1962 576 1980 594
rect 1962 594 1980 612
rect 1962 612 1980 630
rect 1962 630 1980 648
rect 1962 648 1980 666
rect 1962 666 1980 684
rect 1962 684 1980 702
rect 1962 702 1980 720
rect 1962 720 1980 738
rect 1962 738 1980 756
rect 1962 756 1980 774
rect 1962 774 1980 792
rect 1962 792 1980 810
rect 1962 810 1980 828
rect 1962 828 1980 846
rect 1962 846 1980 864
rect 1962 864 1980 882
rect 1962 882 1980 900
rect 1962 900 1980 918
rect 1962 918 1980 936
rect 1962 936 1980 954
rect 1962 954 1980 972
rect 1962 972 1980 990
rect 1962 990 1980 1008
rect 1962 1008 1980 1026
rect 1962 1026 1980 1044
rect 1962 1044 1980 1062
rect 1962 1062 1980 1080
rect 1962 1080 1980 1098
rect 1962 1098 1980 1116
rect 1962 6138 1980 6156
rect 1962 6156 1980 6174
rect 1962 6174 1980 6192
rect 1962 6192 1980 6210
rect 1962 6210 1980 6228
rect 1962 6228 1980 6246
rect 1962 6246 1980 6264
rect 1962 6264 1980 6282
rect 1962 6282 1980 6300
rect 1962 6300 1980 6318
rect 1962 6318 1980 6336
rect 1962 6336 1980 6354
rect 1962 6354 1980 6372
rect 1962 6372 1980 6390
rect 1962 6390 1980 6408
rect 1962 6408 1980 6426
rect 1962 6426 1980 6444
rect 1962 6444 1980 6462
rect 1962 6462 1980 6480
rect 1962 6480 1980 6498
rect 1962 6498 1980 6516
rect 1962 6516 1980 6534
rect 1962 6534 1980 6552
rect 1962 6552 1980 6570
rect 1962 6570 1980 6588
rect 1962 6588 1980 6606
rect 1962 6606 1980 6624
rect 1962 6624 1980 6642
rect 1962 6642 1980 6660
rect 1962 6660 1980 6678
rect 1962 6678 1980 6696
rect 1962 6696 1980 6714
rect 1962 6714 1980 6732
rect 1962 6732 1980 6750
rect 1962 6750 1980 6768
rect 1962 6768 1980 6786
rect 1962 6786 1980 6804
rect 1962 6804 1980 6822
rect 1962 6822 1980 6840
rect 1962 6840 1980 6858
rect 1980 396 1998 414
rect 1980 414 1998 432
rect 1980 432 1998 450
rect 1980 450 1998 468
rect 1980 468 1998 486
rect 1980 486 1998 504
rect 1980 504 1998 522
rect 1980 522 1998 540
rect 1980 540 1998 558
rect 1980 558 1998 576
rect 1980 576 1998 594
rect 1980 594 1998 612
rect 1980 612 1998 630
rect 1980 630 1998 648
rect 1980 648 1998 666
rect 1980 666 1998 684
rect 1980 684 1998 702
rect 1980 702 1998 720
rect 1980 720 1998 738
rect 1980 738 1998 756
rect 1980 756 1998 774
rect 1980 774 1998 792
rect 1980 792 1998 810
rect 1980 810 1998 828
rect 1980 828 1998 846
rect 1980 846 1998 864
rect 1980 864 1998 882
rect 1980 882 1998 900
rect 1980 900 1998 918
rect 1980 918 1998 936
rect 1980 936 1998 954
rect 1980 954 1998 972
rect 1980 972 1998 990
rect 1980 990 1998 1008
rect 1980 1008 1998 1026
rect 1980 1026 1998 1044
rect 1980 1044 1998 1062
rect 1980 1062 1998 1080
rect 1980 1080 1998 1098
rect 1980 1098 1998 1116
rect 1980 6156 1998 6174
rect 1980 6174 1998 6192
rect 1980 6192 1998 6210
rect 1980 6210 1998 6228
rect 1980 6228 1998 6246
rect 1980 6246 1998 6264
rect 1980 6264 1998 6282
rect 1980 6282 1998 6300
rect 1980 6300 1998 6318
rect 1980 6318 1998 6336
rect 1980 6336 1998 6354
rect 1980 6354 1998 6372
rect 1980 6372 1998 6390
rect 1980 6390 1998 6408
rect 1980 6408 1998 6426
rect 1980 6426 1998 6444
rect 1980 6444 1998 6462
rect 1980 6462 1998 6480
rect 1980 6480 1998 6498
rect 1980 6498 1998 6516
rect 1980 6516 1998 6534
rect 1980 6534 1998 6552
rect 1980 6552 1998 6570
rect 1980 6570 1998 6588
rect 1980 6588 1998 6606
rect 1980 6606 1998 6624
rect 1980 6624 1998 6642
rect 1980 6642 1998 6660
rect 1980 6660 1998 6678
rect 1980 6678 1998 6696
rect 1980 6696 1998 6714
rect 1980 6714 1998 6732
rect 1980 6732 1998 6750
rect 1980 6750 1998 6768
rect 1980 6768 1998 6786
rect 1980 6786 1998 6804
rect 1980 6804 1998 6822
rect 1980 6822 1998 6840
rect 1980 6840 1998 6858
rect 1980 6858 1998 6876
rect 1998 378 2016 396
rect 1998 396 2016 414
rect 1998 414 2016 432
rect 1998 432 2016 450
rect 1998 450 2016 468
rect 1998 468 2016 486
rect 1998 486 2016 504
rect 1998 504 2016 522
rect 1998 522 2016 540
rect 1998 540 2016 558
rect 1998 558 2016 576
rect 1998 576 2016 594
rect 1998 594 2016 612
rect 1998 612 2016 630
rect 1998 630 2016 648
rect 1998 648 2016 666
rect 1998 666 2016 684
rect 1998 684 2016 702
rect 1998 702 2016 720
rect 1998 720 2016 738
rect 1998 738 2016 756
rect 1998 756 2016 774
rect 1998 774 2016 792
rect 1998 792 2016 810
rect 1998 810 2016 828
rect 1998 828 2016 846
rect 1998 846 2016 864
rect 1998 864 2016 882
rect 1998 882 2016 900
rect 1998 900 2016 918
rect 1998 918 2016 936
rect 1998 936 2016 954
rect 1998 954 2016 972
rect 1998 972 2016 990
rect 1998 990 2016 1008
rect 1998 1008 2016 1026
rect 1998 1026 2016 1044
rect 1998 1044 2016 1062
rect 1998 1062 2016 1080
rect 1998 1080 2016 1098
rect 1998 6156 2016 6174
rect 1998 6174 2016 6192
rect 1998 6192 2016 6210
rect 1998 6210 2016 6228
rect 1998 6228 2016 6246
rect 1998 6246 2016 6264
rect 1998 6264 2016 6282
rect 1998 6282 2016 6300
rect 1998 6300 2016 6318
rect 1998 6318 2016 6336
rect 1998 6336 2016 6354
rect 1998 6354 2016 6372
rect 1998 6372 2016 6390
rect 1998 6390 2016 6408
rect 1998 6408 2016 6426
rect 1998 6426 2016 6444
rect 1998 6444 2016 6462
rect 1998 6462 2016 6480
rect 1998 6480 2016 6498
rect 1998 6498 2016 6516
rect 1998 6516 2016 6534
rect 1998 6534 2016 6552
rect 1998 6552 2016 6570
rect 1998 6570 2016 6588
rect 1998 6588 2016 6606
rect 1998 6606 2016 6624
rect 1998 6624 2016 6642
rect 1998 6642 2016 6660
rect 1998 6660 2016 6678
rect 1998 6678 2016 6696
rect 1998 6696 2016 6714
rect 1998 6714 2016 6732
rect 1998 6732 2016 6750
rect 1998 6750 2016 6768
rect 1998 6768 2016 6786
rect 1998 6786 2016 6804
rect 1998 6804 2016 6822
rect 1998 6822 2016 6840
rect 1998 6840 2016 6858
rect 1998 6858 2016 6876
rect 2016 360 2034 378
rect 2016 378 2034 396
rect 2016 396 2034 414
rect 2016 414 2034 432
rect 2016 432 2034 450
rect 2016 450 2034 468
rect 2016 468 2034 486
rect 2016 486 2034 504
rect 2016 504 2034 522
rect 2016 522 2034 540
rect 2016 540 2034 558
rect 2016 558 2034 576
rect 2016 576 2034 594
rect 2016 594 2034 612
rect 2016 612 2034 630
rect 2016 630 2034 648
rect 2016 648 2034 666
rect 2016 666 2034 684
rect 2016 684 2034 702
rect 2016 702 2034 720
rect 2016 720 2034 738
rect 2016 738 2034 756
rect 2016 756 2034 774
rect 2016 774 2034 792
rect 2016 792 2034 810
rect 2016 810 2034 828
rect 2016 828 2034 846
rect 2016 846 2034 864
rect 2016 864 2034 882
rect 2016 882 2034 900
rect 2016 900 2034 918
rect 2016 918 2034 936
rect 2016 936 2034 954
rect 2016 954 2034 972
rect 2016 972 2034 990
rect 2016 990 2034 1008
rect 2016 1008 2034 1026
rect 2016 1026 2034 1044
rect 2016 1044 2034 1062
rect 2016 1062 2034 1080
rect 2016 6174 2034 6192
rect 2016 6192 2034 6210
rect 2016 6210 2034 6228
rect 2016 6228 2034 6246
rect 2016 6246 2034 6264
rect 2016 6264 2034 6282
rect 2016 6282 2034 6300
rect 2016 6300 2034 6318
rect 2016 6318 2034 6336
rect 2016 6336 2034 6354
rect 2016 6354 2034 6372
rect 2016 6372 2034 6390
rect 2016 6390 2034 6408
rect 2016 6408 2034 6426
rect 2016 6426 2034 6444
rect 2016 6444 2034 6462
rect 2016 6462 2034 6480
rect 2016 6480 2034 6498
rect 2016 6498 2034 6516
rect 2016 6516 2034 6534
rect 2016 6534 2034 6552
rect 2016 6552 2034 6570
rect 2016 6570 2034 6588
rect 2016 6588 2034 6606
rect 2016 6606 2034 6624
rect 2016 6624 2034 6642
rect 2016 6642 2034 6660
rect 2016 6660 2034 6678
rect 2016 6678 2034 6696
rect 2016 6696 2034 6714
rect 2016 6714 2034 6732
rect 2016 6732 2034 6750
rect 2016 6750 2034 6768
rect 2016 6768 2034 6786
rect 2016 6786 2034 6804
rect 2016 6804 2034 6822
rect 2016 6822 2034 6840
rect 2016 6840 2034 6858
rect 2016 6858 2034 6876
rect 2016 6876 2034 6894
rect 2034 360 2052 378
rect 2034 378 2052 396
rect 2034 396 2052 414
rect 2034 414 2052 432
rect 2034 432 2052 450
rect 2034 450 2052 468
rect 2034 468 2052 486
rect 2034 486 2052 504
rect 2034 504 2052 522
rect 2034 522 2052 540
rect 2034 540 2052 558
rect 2034 558 2052 576
rect 2034 576 2052 594
rect 2034 594 2052 612
rect 2034 612 2052 630
rect 2034 630 2052 648
rect 2034 648 2052 666
rect 2034 666 2052 684
rect 2034 684 2052 702
rect 2034 702 2052 720
rect 2034 720 2052 738
rect 2034 738 2052 756
rect 2034 756 2052 774
rect 2034 774 2052 792
rect 2034 792 2052 810
rect 2034 810 2052 828
rect 2034 828 2052 846
rect 2034 846 2052 864
rect 2034 864 2052 882
rect 2034 882 2052 900
rect 2034 900 2052 918
rect 2034 918 2052 936
rect 2034 936 2052 954
rect 2034 954 2052 972
rect 2034 972 2052 990
rect 2034 990 2052 1008
rect 2034 1008 2052 1026
rect 2034 1026 2052 1044
rect 2034 1044 2052 1062
rect 2034 1062 2052 1080
rect 2034 6192 2052 6210
rect 2034 6210 2052 6228
rect 2034 6228 2052 6246
rect 2034 6246 2052 6264
rect 2034 6264 2052 6282
rect 2034 6282 2052 6300
rect 2034 6300 2052 6318
rect 2034 6318 2052 6336
rect 2034 6336 2052 6354
rect 2034 6354 2052 6372
rect 2034 6372 2052 6390
rect 2034 6390 2052 6408
rect 2034 6408 2052 6426
rect 2034 6426 2052 6444
rect 2034 6444 2052 6462
rect 2034 6462 2052 6480
rect 2034 6480 2052 6498
rect 2034 6498 2052 6516
rect 2034 6516 2052 6534
rect 2034 6534 2052 6552
rect 2034 6552 2052 6570
rect 2034 6570 2052 6588
rect 2034 6588 2052 6606
rect 2034 6606 2052 6624
rect 2034 6624 2052 6642
rect 2034 6642 2052 6660
rect 2034 6660 2052 6678
rect 2034 6678 2052 6696
rect 2034 6696 2052 6714
rect 2034 6714 2052 6732
rect 2034 6732 2052 6750
rect 2034 6750 2052 6768
rect 2034 6768 2052 6786
rect 2034 6786 2052 6804
rect 2034 6804 2052 6822
rect 2034 6822 2052 6840
rect 2034 6840 2052 6858
rect 2034 6858 2052 6876
rect 2034 6876 2052 6894
rect 2052 342 2070 360
rect 2052 360 2070 378
rect 2052 378 2070 396
rect 2052 396 2070 414
rect 2052 414 2070 432
rect 2052 432 2070 450
rect 2052 450 2070 468
rect 2052 468 2070 486
rect 2052 486 2070 504
rect 2052 504 2070 522
rect 2052 522 2070 540
rect 2052 540 2070 558
rect 2052 558 2070 576
rect 2052 576 2070 594
rect 2052 594 2070 612
rect 2052 612 2070 630
rect 2052 630 2070 648
rect 2052 648 2070 666
rect 2052 666 2070 684
rect 2052 684 2070 702
rect 2052 702 2070 720
rect 2052 720 2070 738
rect 2052 738 2070 756
rect 2052 756 2070 774
rect 2052 774 2070 792
rect 2052 792 2070 810
rect 2052 810 2070 828
rect 2052 828 2070 846
rect 2052 846 2070 864
rect 2052 864 2070 882
rect 2052 882 2070 900
rect 2052 900 2070 918
rect 2052 918 2070 936
rect 2052 936 2070 954
rect 2052 954 2070 972
rect 2052 972 2070 990
rect 2052 990 2070 1008
rect 2052 1008 2070 1026
rect 2052 1026 2070 1044
rect 2052 1044 2070 1062
rect 2052 6192 2070 6210
rect 2052 6210 2070 6228
rect 2052 6228 2070 6246
rect 2052 6246 2070 6264
rect 2052 6264 2070 6282
rect 2052 6282 2070 6300
rect 2052 6300 2070 6318
rect 2052 6318 2070 6336
rect 2052 6336 2070 6354
rect 2052 6354 2070 6372
rect 2052 6372 2070 6390
rect 2052 6390 2070 6408
rect 2052 6408 2070 6426
rect 2052 6426 2070 6444
rect 2052 6444 2070 6462
rect 2052 6462 2070 6480
rect 2052 6480 2070 6498
rect 2052 6498 2070 6516
rect 2052 6516 2070 6534
rect 2052 6534 2070 6552
rect 2052 6552 2070 6570
rect 2052 6570 2070 6588
rect 2052 6588 2070 6606
rect 2052 6606 2070 6624
rect 2052 6624 2070 6642
rect 2052 6642 2070 6660
rect 2052 6660 2070 6678
rect 2052 6678 2070 6696
rect 2052 6696 2070 6714
rect 2052 6714 2070 6732
rect 2052 6732 2070 6750
rect 2052 6750 2070 6768
rect 2052 6768 2070 6786
rect 2052 6786 2070 6804
rect 2052 6804 2070 6822
rect 2052 6822 2070 6840
rect 2052 6840 2070 6858
rect 2052 6858 2070 6876
rect 2052 6876 2070 6894
rect 2052 6894 2070 6912
rect 2070 342 2088 360
rect 2070 360 2088 378
rect 2070 378 2088 396
rect 2070 396 2088 414
rect 2070 414 2088 432
rect 2070 432 2088 450
rect 2070 450 2088 468
rect 2070 468 2088 486
rect 2070 486 2088 504
rect 2070 504 2088 522
rect 2070 522 2088 540
rect 2070 540 2088 558
rect 2070 558 2088 576
rect 2070 576 2088 594
rect 2070 594 2088 612
rect 2070 612 2088 630
rect 2070 630 2088 648
rect 2070 648 2088 666
rect 2070 666 2088 684
rect 2070 684 2088 702
rect 2070 702 2088 720
rect 2070 720 2088 738
rect 2070 738 2088 756
rect 2070 756 2088 774
rect 2070 774 2088 792
rect 2070 792 2088 810
rect 2070 810 2088 828
rect 2070 828 2088 846
rect 2070 846 2088 864
rect 2070 864 2088 882
rect 2070 882 2088 900
rect 2070 900 2088 918
rect 2070 918 2088 936
rect 2070 936 2088 954
rect 2070 954 2088 972
rect 2070 972 2088 990
rect 2070 990 2088 1008
rect 2070 1008 2088 1026
rect 2070 1026 2088 1044
rect 2070 6210 2088 6228
rect 2070 6228 2088 6246
rect 2070 6246 2088 6264
rect 2070 6264 2088 6282
rect 2070 6282 2088 6300
rect 2070 6300 2088 6318
rect 2070 6318 2088 6336
rect 2070 6336 2088 6354
rect 2070 6354 2088 6372
rect 2070 6372 2088 6390
rect 2070 6390 2088 6408
rect 2070 6408 2088 6426
rect 2070 6426 2088 6444
rect 2070 6444 2088 6462
rect 2070 6462 2088 6480
rect 2070 6480 2088 6498
rect 2070 6498 2088 6516
rect 2070 6516 2088 6534
rect 2070 6534 2088 6552
rect 2070 6552 2088 6570
rect 2070 6570 2088 6588
rect 2070 6588 2088 6606
rect 2070 6606 2088 6624
rect 2070 6624 2088 6642
rect 2070 6642 2088 6660
rect 2070 6660 2088 6678
rect 2070 6678 2088 6696
rect 2070 6696 2088 6714
rect 2070 6714 2088 6732
rect 2070 6732 2088 6750
rect 2070 6750 2088 6768
rect 2070 6768 2088 6786
rect 2070 6786 2088 6804
rect 2070 6804 2088 6822
rect 2070 6822 2088 6840
rect 2070 6840 2088 6858
rect 2070 6858 2088 6876
rect 2070 6876 2088 6894
rect 2070 6894 2088 6912
rect 2088 324 2106 342
rect 2088 342 2106 360
rect 2088 360 2106 378
rect 2088 378 2106 396
rect 2088 396 2106 414
rect 2088 414 2106 432
rect 2088 432 2106 450
rect 2088 450 2106 468
rect 2088 468 2106 486
rect 2088 486 2106 504
rect 2088 504 2106 522
rect 2088 522 2106 540
rect 2088 540 2106 558
rect 2088 558 2106 576
rect 2088 576 2106 594
rect 2088 594 2106 612
rect 2088 612 2106 630
rect 2088 630 2106 648
rect 2088 648 2106 666
rect 2088 666 2106 684
rect 2088 684 2106 702
rect 2088 702 2106 720
rect 2088 720 2106 738
rect 2088 738 2106 756
rect 2088 756 2106 774
rect 2088 774 2106 792
rect 2088 792 2106 810
rect 2088 810 2106 828
rect 2088 828 2106 846
rect 2088 846 2106 864
rect 2088 864 2106 882
rect 2088 882 2106 900
rect 2088 900 2106 918
rect 2088 918 2106 936
rect 2088 936 2106 954
rect 2088 954 2106 972
rect 2088 972 2106 990
rect 2088 990 2106 1008
rect 2088 1008 2106 1026
rect 2088 1026 2106 1044
rect 2088 6228 2106 6246
rect 2088 6246 2106 6264
rect 2088 6264 2106 6282
rect 2088 6282 2106 6300
rect 2088 6300 2106 6318
rect 2088 6318 2106 6336
rect 2088 6336 2106 6354
rect 2088 6354 2106 6372
rect 2088 6372 2106 6390
rect 2088 6390 2106 6408
rect 2088 6408 2106 6426
rect 2088 6426 2106 6444
rect 2088 6444 2106 6462
rect 2088 6462 2106 6480
rect 2088 6480 2106 6498
rect 2088 6498 2106 6516
rect 2088 6516 2106 6534
rect 2088 6534 2106 6552
rect 2088 6552 2106 6570
rect 2088 6570 2106 6588
rect 2088 6588 2106 6606
rect 2088 6606 2106 6624
rect 2088 6624 2106 6642
rect 2088 6642 2106 6660
rect 2088 6660 2106 6678
rect 2088 6678 2106 6696
rect 2088 6696 2106 6714
rect 2088 6714 2106 6732
rect 2088 6732 2106 6750
rect 2088 6750 2106 6768
rect 2088 6768 2106 6786
rect 2088 6786 2106 6804
rect 2088 6804 2106 6822
rect 2088 6822 2106 6840
rect 2088 6840 2106 6858
rect 2088 6858 2106 6876
rect 2088 6876 2106 6894
rect 2088 6894 2106 6912
rect 2088 6912 2106 6930
rect 2106 324 2124 342
rect 2106 342 2124 360
rect 2106 360 2124 378
rect 2106 378 2124 396
rect 2106 396 2124 414
rect 2106 414 2124 432
rect 2106 432 2124 450
rect 2106 450 2124 468
rect 2106 468 2124 486
rect 2106 486 2124 504
rect 2106 504 2124 522
rect 2106 522 2124 540
rect 2106 540 2124 558
rect 2106 558 2124 576
rect 2106 576 2124 594
rect 2106 594 2124 612
rect 2106 612 2124 630
rect 2106 630 2124 648
rect 2106 648 2124 666
rect 2106 666 2124 684
rect 2106 684 2124 702
rect 2106 702 2124 720
rect 2106 720 2124 738
rect 2106 738 2124 756
rect 2106 756 2124 774
rect 2106 774 2124 792
rect 2106 792 2124 810
rect 2106 810 2124 828
rect 2106 828 2124 846
rect 2106 846 2124 864
rect 2106 864 2124 882
rect 2106 882 2124 900
rect 2106 900 2124 918
rect 2106 918 2124 936
rect 2106 936 2124 954
rect 2106 954 2124 972
rect 2106 972 2124 990
rect 2106 990 2124 1008
rect 2106 1008 2124 1026
rect 2106 6228 2124 6246
rect 2106 6246 2124 6264
rect 2106 6264 2124 6282
rect 2106 6282 2124 6300
rect 2106 6300 2124 6318
rect 2106 6318 2124 6336
rect 2106 6336 2124 6354
rect 2106 6354 2124 6372
rect 2106 6372 2124 6390
rect 2106 6390 2124 6408
rect 2106 6408 2124 6426
rect 2106 6426 2124 6444
rect 2106 6444 2124 6462
rect 2106 6462 2124 6480
rect 2106 6480 2124 6498
rect 2106 6498 2124 6516
rect 2106 6516 2124 6534
rect 2106 6534 2124 6552
rect 2106 6552 2124 6570
rect 2106 6570 2124 6588
rect 2106 6588 2124 6606
rect 2106 6606 2124 6624
rect 2106 6624 2124 6642
rect 2106 6642 2124 6660
rect 2106 6660 2124 6678
rect 2106 6678 2124 6696
rect 2106 6696 2124 6714
rect 2106 6714 2124 6732
rect 2106 6732 2124 6750
rect 2106 6750 2124 6768
rect 2106 6768 2124 6786
rect 2106 6786 2124 6804
rect 2106 6804 2124 6822
rect 2106 6822 2124 6840
rect 2106 6840 2124 6858
rect 2106 6858 2124 6876
rect 2106 6876 2124 6894
rect 2106 6894 2124 6912
rect 2106 6912 2124 6930
rect 2124 306 2142 324
rect 2124 324 2142 342
rect 2124 342 2142 360
rect 2124 360 2142 378
rect 2124 378 2142 396
rect 2124 396 2142 414
rect 2124 414 2142 432
rect 2124 432 2142 450
rect 2124 450 2142 468
rect 2124 468 2142 486
rect 2124 486 2142 504
rect 2124 504 2142 522
rect 2124 522 2142 540
rect 2124 540 2142 558
rect 2124 558 2142 576
rect 2124 576 2142 594
rect 2124 594 2142 612
rect 2124 612 2142 630
rect 2124 630 2142 648
rect 2124 648 2142 666
rect 2124 666 2142 684
rect 2124 684 2142 702
rect 2124 702 2142 720
rect 2124 720 2142 738
rect 2124 738 2142 756
rect 2124 756 2142 774
rect 2124 774 2142 792
rect 2124 792 2142 810
rect 2124 810 2142 828
rect 2124 828 2142 846
rect 2124 846 2142 864
rect 2124 864 2142 882
rect 2124 882 2142 900
rect 2124 900 2142 918
rect 2124 918 2142 936
rect 2124 936 2142 954
rect 2124 954 2142 972
rect 2124 972 2142 990
rect 2124 990 2142 1008
rect 2124 1008 2142 1026
rect 2124 6246 2142 6264
rect 2124 6264 2142 6282
rect 2124 6282 2142 6300
rect 2124 6300 2142 6318
rect 2124 6318 2142 6336
rect 2124 6336 2142 6354
rect 2124 6354 2142 6372
rect 2124 6372 2142 6390
rect 2124 6390 2142 6408
rect 2124 6408 2142 6426
rect 2124 6426 2142 6444
rect 2124 6444 2142 6462
rect 2124 6462 2142 6480
rect 2124 6480 2142 6498
rect 2124 6498 2142 6516
rect 2124 6516 2142 6534
rect 2124 6534 2142 6552
rect 2124 6552 2142 6570
rect 2124 6570 2142 6588
rect 2124 6588 2142 6606
rect 2124 6606 2142 6624
rect 2124 6624 2142 6642
rect 2124 6642 2142 6660
rect 2124 6660 2142 6678
rect 2124 6678 2142 6696
rect 2124 6696 2142 6714
rect 2124 6714 2142 6732
rect 2124 6732 2142 6750
rect 2124 6750 2142 6768
rect 2124 6768 2142 6786
rect 2124 6786 2142 6804
rect 2124 6804 2142 6822
rect 2124 6822 2142 6840
rect 2124 6840 2142 6858
rect 2124 6858 2142 6876
rect 2124 6876 2142 6894
rect 2124 6894 2142 6912
rect 2124 6912 2142 6930
rect 2124 6930 2142 6948
rect 2142 378 2160 396
rect 2142 396 2160 414
rect 2142 414 2160 432
rect 2142 432 2160 450
rect 2142 450 2160 468
rect 2142 468 2160 486
rect 2142 486 2160 504
rect 2142 504 2160 522
rect 2142 522 2160 540
rect 2142 540 2160 558
rect 2142 558 2160 576
rect 2142 576 2160 594
rect 2142 594 2160 612
rect 2142 612 2160 630
rect 2142 630 2160 648
rect 2142 648 2160 666
rect 2142 666 2160 684
rect 2142 684 2160 702
rect 2142 702 2160 720
rect 2142 720 2160 738
rect 2142 738 2160 756
rect 2142 756 2160 774
rect 2142 774 2160 792
rect 2142 792 2160 810
rect 2142 810 2160 828
rect 2142 828 2160 846
rect 2142 846 2160 864
rect 2142 864 2160 882
rect 2142 882 2160 900
rect 2142 900 2160 918
rect 2142 918 2160 936
rect 2142 936 2160 954
rect 2142 954 2160 972
rect 2142 972 2160 990
rect 2142 990 2160 1008
rect 2142 6246 2160 6264
rect 2142 6264 2160 6282
rect 2142 6282 2160 6300
rect 2142 6300 2160 6318
rect 2142 6318 2160 6336
rect 2142 6336 2160 6354
rect 2142 6354 2160 6372
rect 2142 6372 2160 6390
rect 2142 6390 2160 6408
rect 2142 6408 2160 6426
rect 2142 6426 2160 6444
rect 2142 6444 2160 6462
rect 2142 6462 2160 6480
rect 2142 6480 2160 6498
rect 2142 6498 2160 6516
rect 2142 6516 2160 6534
rect 2142 6534 2160 6552
rect 2142 6552 2160 6570
rect 2142 6570 2160 6588
rect 2142 6588 2160 6606
rect 2142 6606 2160 6624
rect 2142 6624 2160 6642
rect 2142 6642 2160 6660
rect 2142 6660 2160 6678
rect 2142 6678 2160 6696
rect 2142 6696 2160 6714
rect 2142 6714 2160 6732
rect 2142 6732 2160 6750
rect 2142 6750 2160 6768
rect 2142 6768 2160 6786
rect 2142 6786 2160 6804
rect 2142 6804 2160 6822
rect 2142 6822 2160 6840
rect 2142 6840 2160 6858
rect 2142 6858 2160 6876
rect 2142 6876 2160 6894
rect 2142 6894 2160 6912
rect 2142 6912 2160 6930
rect 2142 6930 2160 6948
rect 2160 522 2178 540
rect 2160 540 2178 558
rect 2160 558 2178 576
rect 2160 576 2178 594
rect 2160 594 2178 612
rect 2160 612 2178 630
rect 2160 630 2178 648
rect 2160 648 2178 666
rect 2160 666 2178 684
rect 2160 684 2178 702
rect 2160 702 2178 720
rect 2160 720 2178 738
rect 2160 738 2178 756
rect 2160 756 2178 774
rect 2160 774 2178 792
rect 2160 792 2178 810
rect 2160 810 2178 828
rect 2160 828 2178 846
rect 2160 846 2178 864
rect 2160 864 2178 882
rect 2160 882 2178 900
rect 2160 900 2178 918
rect 2160 918 2178 936
rect 2160 936 2178 954
rect 2160 954 2178 972
rect 2160 972 2178 990
rect 2160 990 2178 1008
rect 2160 6264 2178 6282
rect 2160 6282 2178 6300
rect 2160 6300 2178 6318
rect 2160 6318 2178 6336
rect 2160 6336 2178 6354
rect 2160 6354 2178 6372
rect 2160 6372 2178 6390
rect 2160 6390 2178 6408
rect 2160 6408 2178 6426
rect 2160 6426 2178 6444
rect 2160 6444 2178 6462
rect 2160 6462 2178 6480
rect 2160 6480 2178 6498
rect 2160 6498 2178 6516
rect 2160 6516 2178 6534
rect 2160 6534 2178 6552
rect 2160 6552 2178 6570
rect 2160 6570 2178 6588
rect 2160 6588 2178 6606
rect 2160 6606 2178 6624
rect 2160 6624 2178 6642
rect 2160 6642 2178 6660
rect 2160 6660 2178 6678
rect 2160 6678 2178 6696
rect 2160 6696 2178 6714
rect 2160 6714 2178 6732
rect 2160 6732 2178 6750
rect 2160 6750 2178 6768
rect 2160 6768 2178 6786
rect 2160 6786 2178 6804
rect 2160 6804 2178 6822
rect 2160 6822 2178 6840
rect 2160 6840 2178 6858
rect 2160 6858 2178 6876
rect 2160 6876 2178 6894
rect 2160 6894 2178 6912
rect 2160 6912 2178 6930
rect 2160 6930 2178 6948
rect 2160 6948 2178 6966
rect 2178 666 2196 684
rect 2178 684 2196 702
rect 2178 702 2196 720
rect 2178 720 2196 738
rect 2178 738 2196 756
rect 2178 756 2196 774
rect 2178 774 2196 792
rect 2178 792 2196 810
rect 2178 810 2196 828
rect 2178 828 2196 846
rect 2178 846 2196 864
rect 2178 864 2196 882
rect 2178 882 2196 900
rect 2178 900 2196 918
rect 2178 918 2196 936
rect 2178 936 2196 954
rect 2178 954 2196 972
rect 2178 972 2196 990
rect 2178 6264 2196 6282
rect 2178 6282 2196 6300
rect 2178 6300 2196 6318
rect 2178 6318 2196 6336
rect 2178 6336 2196 6354
rect 2178 6354 2196 6372
rect 2178 6372 2196 6390
rect 2178 6390 2196 6408
rect 2178 6408 2196 6426
rect 2178 6426 2196 6444
rect 2178 6444 2196 6462
rect 2178 6462 2196 6480
rect 2178 6480 2196 6498
rect 2178 6498 2196 6516
rect 2178 6516 2196 6534
rect 2178 6534 2196 6552
rect 2178 6552 2196 6570
rect 2178 6570 2196 6588
rect 2178 6588 2196 6606
rect 2178 6606 2196 6624
rect 2178 6624 2196 6642
rect 2178 6642 2196 6660
rect 2178 6660 2196 6678
rect 2178 6678 2196 6696
rect 2178 6696 2196 6714
rect 2178 6714 2196 6732
rect 2178 6732 2196 6750
rect 2178 6750 2196 6768
rect 2178 6768 2196 6786
rect 2178 6786 2196 6804
rect 2178 6804 2196 6822
rect 2178 6822 2196 6840
rect 2178 6840 2196 6858
rect 2178 6858 2196 6876
rect 2178 6876 2196 6894
rect 2178 6894 2196 6912
rect 2178 6912 2196 6930
rect 2178 6930 2196 6948
rect 2178 6948 2196 6966
rect 2196 828 2214 846
rect 2196 846 2214 864
rect 2196 864 2214 882
rect 2196 882 2214 900
rect 2196 900 2214 918
rect 2196 918 2214 936
rect 2196 936 2214 954
rect 2196 954 2214 972
rect 2196 972 2214 990
rect 2196 6282 2214 6300
rect 2196 6300 2214 6318
rect 2196 6318 2214 6336
rect 2196 6336 2214 6354
rect 2196 6354 2214 6372
rect 2196 6372 2214 6390
rect 2196 6390 2214 6408
rect 2196 6408 2214 6426
rect 2196 6426 2214 6444
rect 2196 6444 2214 6462
rect 2196 6462 2214 6480
rect 2196 6480 2214 6498
rect 2196 6498 2214 6516
rect 2196 6516 2214 6534
rect 2196 6534 2214 6552
rect 2196 6552 2214 6570
rect 2196 6570 2214 6588
rect 2196 6588 2214 6606
rect 2196 6606 2214 6624
rect 2196 6624 2214 6642
rect 2196 6642 2214 6660
rect 2196 6660 2214 6678
rect 2196 6678 2214 6696
rect 2196 6696 2214 6714
rect 2196 6714 2214 6732
rect 2196 6732 2214 6750
rect 2196 6750 2214 6768
rect 2196 6768 2214 6786
rect 2196 6786 2214 6804
rect 2196 6804 2214 6822
rect 2196 6822 2214 6840
rect 2196 6840 2214 6858
rect 2196 6858 2214 6876
rect 2196 6876 2214 6894
rect 2196 6894 2214 6912
rect 2196 6912 2214 6930
rect 2196 6930 2214 6948
rect 2196 6948 2214 6966
rect 2196 6966 2214 6984
rect 2214 6300 2232 6318
rect 2214 6318 2232 6336
rect 2214 6336 2232 6354
rect 2214 6354 2232 6372
rect 2214 6372 2232 6390
rect 2214 6390 2232 6408
rect 2214 6408 2232 6426
rect 2214 6426 2232 6444
rect 2214 6444 2232 6462
rect 2214 6462 2232 6480
rect 2214 6480 2232 6498
rect 2214 6498 2232 6516
rect 2214 6516 2232 6534
rect 2214 6534 2232 6552
rect 2214 6552 2232 6570
rect 2214 6570 2232 6588
rect 2214 6588 2232 6606
rect 2214 6606 2232 6624
rect 2214 6624 2232 6642
rect 2214 6642 2232 6660
rect 2214 6660 2232 6678
rect 2214 6678 2232 6696
rect 2214 6696 2232 6714
rect 2214 6714 2232 6732
rect 2214 6732 2232 6750
rect 2214 6750 2232 6768
rect 2214 6768 2232 6786
rect 2214 6786 2232 6804
rect 2214 6804 2232 6822
rect 2214 6822 2232 6840
rect 2214 6840 2232 6858
rect 2214 6858 2232 6876
rect 2214 6876 2232 6894
rect 2214 6894 2232 6912
rect 2214 6912 2232 6930
rect 2214 6930 2232 6948
rect 2214 6948 2232 6966
rect 2214 6966 2232 6984
rect 2232 6300 2250 6318
rect 2232 6318 2250 6336
rect 2232 6336 2250 6354
rect 2232 6354 2250 6372
rect 2232 6372 2250 6390
rect 2232 6390 2250 6408
rect 2232 6408 2250 6426
rect 2232 6426 2250 6444
rect 2232 6444 2250 6462
rect 2232 6462 2250 6480
rect 2232 6480 2250 6498
rect 2232 6498 2250 6516
rect 2232 6516 2250 6534
rect 2232 6534 2250 6552
rect 2232 6552 2250 6570
rect 2232 6570 2250 6588
rect 2232 6588 2250 6606
rect 2232 6606 2250 6624
rect 2232 6624 2250 6642
rect 2232 6642 2250 6660
rect 2232 6660 2250 6678
rect 2232 6678 2250 6696
rect 2232 6696 2250 6714
rect 2232 6714 2250 6732
rect 2232 6732 2250 6750
rect 2232 6750 2250 6768
rect 2232 6768 2250 6786
rect 2232 6786 2250 6804
rect 2232 6804 2250 6822
rect 2232 6822 2250 6840
rect 2232 6840 2250 6858
rect 2232 6858 2250 6876
rect 2232 6876 2250 6894
rect 2232 6894 2250 6912
rect 2232 6912 2250 6930
rect 2232 6930 2250 6948
rect 2232 6948 2250 6966
rect 2232 6966 2250 6984
rect 2250 6318 2268 6336
rect 2250 6336 2268 6354
rect 2250 6354 2268 6372
rect 2250 6372 2268 6390
rect 2250 6390 2268 6408
rect 2250 6408 2268 6426
rect 2250 6426 2268 6444
rect 2250 6444 2268 6462
rect 2250 6462 2268 6480
rect 2250 6480 2268 6498
rect 2250 6498 2268 6516
rect 2250 6516 2268 6534
rect 2250 6534 2268 6552
rect 2250 6552 2268 6570
rect 2250 6570 2268 6588
rect 2250 6588 2268 6606
rect 2250 6606 2268 6624
rect 2250 6624 2268 6642
rect 2250 6642 2268 6660
rect 2250 6660 2268 6678
rect 2250 6678 2268 6696
rect 2250 6696 2268 6714
rect 2250 6714 2268 6732
rect 2250 6732 2268 6750
rect 2250 6750 2268 6768
rect 2250 6768 2268 6786
rect 2250 6786 2268 6804
rect 2250 6804 2268 6822
rect 2250 6822 2268 6840
rect 2250 6840 2268 6858
rect 2250 6858 2268 6876
rect 2250 6876 2268 6894
rect 2250 6894 2268 6912
rect 2250 6912 2268 6930
rect 2250 6930 2268 6948
rect 2250 6948 2268 6966
rect 2250 6966 2268 6984
rect 2250 6984 2268 7002
rect 2268 6318 2286 6336
rect 2268 6336 2286 6354
rect 2268 6354 2286 6372
rect 2268 6372 2286 6390
rect 2268 6390 2286 6408
rect 2268 6408 2286 6426
rect 2268 6426 2286 6444
rect 2268 6444 2286 6462
rect 2268 6462 2286 6480
rect 2268 6480 2286 6498
rect 2268 6498 2286 6516
rect 2268 6516 2286 6534
rect 2268 6534 2286 6552
rect 2268 6552 2286 6570
rect 2268 6570 2286 6588
rect 2268 6588 2286 6606
rect 2268 6606 2286 6624
rect 2268 6624 2286 6642
rect 2268 6642 2286 6660
rect 2268 6660 2286 6678
rect 2268 6678 2286 6696
rect 2268 6696 2286 6714
rect 2268 6714 2286 6732
rect 2268 6732 2286 6750
rect 2268 6750 2286 6768
rect 2268 6768 2286 6786
rect 2268 6786 2286 6804
rect 2268 6804 2286 6822
rect 2268 6822 2286 6840
rect 2268 6840 2286 6858
rect 2268 6858 2286 6876
rect 2268 6876 2286 6894
rect 2268 6894 2286 6912
rect 2268 6912 2286 6930
rect 2268 6930 2286 6948
rect 2268 6948 2286 6966
rect 2268 6966 2286 6984
rect 2268 6984 2286 7002
rect 2286 6336 2304 6354
rect 2286 6354 2304 6372
rect 2286 6372 2304 6390
rect 2286 6390 2304 6408
rect 2286 6408 2304 6426
rect 2286 6426 2304 6444
rect 2286 6444 2304 6462
rect 2286 6462 2304 6480
rect 2286 6480 2304 6498
rect 2286 6498 2304 6516
rect 2286 6516 2304 6534
rect 2286 6534 2304 6552
rect 2286 6552 2304 6570
rect 2286 6570 2304 6588
rect 2286 6588 2304 6606
rect 2286 6606 2304 6624
rect 2286 6624 2304 6642
rect 2286 6642 2304 6660
rect 2286 6660 2304 6678
rect 2286 6678 2304 6696
rect 2286 6696 2304 6714
rect 2286 6714 2304 6732
rect 2286 6732 2304 6750
rect 2286 6750 2304 6768
rect 2286 6768 2304 6786
rect 2286 6786 2304 6804
rect 2286 6804 2304 6822
rect 2286 6822 2304 6840
rect 2286 6840 2304 6858
rect 2286 6858 2304 6876
rect 2286 6876 2304 6894
rect 2286 6894 2304 6912
rect 2286 6912 2304 6930
rect 2286 6930 2304 6948
rect 2286 6948 2304 6966
rect 2286 6966 2304 6984
rect 2286 6984 2304 7002
rect 2286 7002 2304 7020
rect 2304 360 2322 378
rect 2304 378 2322 396
rect 2304 396 2322 414
rect 2304 414 2322 432
rect 2304 6336 2322 6354
rect 2304 6354 2322 6372
rect 2304 6372 2322 6390
rect 2304 6390 2322 6408
rect 2304 6408 2322 6426
rect 2304 6426 2322 6444
rect 2304 6444 2322 6462
rect 2304 6462 2322 6480
rect 2304 6480 2322 6498
rect 2304 6498 2322 6516
rect 2304 6516 2322 6534
rect 2304 6534 2322 6552
rect 2304 6552 2322 6570
rect 2304 6570 2322 6588
rect 2304 6588 2322 6606
rect 2304 6606 2322 6624
rect 2304 6624 2322 6642
rect 2304 6642 2322 6660
rect 2304 6660 2322 6678
rect 2304 6678 2322 6696
rect 2304 6696 2322 6714
rect 2304 6714 2322 6732
rect 2304 6732 2322 6750
rect 2304 6750 2322 6768
rect 2304 6768 2322 6786
rect 2304 6786 2322 6804
rect 2304 6804 2322 6822
rect 2304 6822 2322 6840
rect 2304 6840 2322 6858
rect 2304 6858 2322 6876
rect 2304 6876 2322 6894
rect 2304 6894 2322 6912
rect 2304 6912 2322 6930
rect 2304 6930 2322 6948
rect 2304 6948 2322 6966
rect 2304 6966 2322 6984
rect 2304 6984 2322 7002
rect 2304 7002 2322 7020
rect 2322 396 2340 414
rect 2322 414 2340 432
rect 2322 432 2340 450
rect 2322 450 2340 468
rect 2322 468 2340 486
rect 2322 486 2340 504
rect 2322 504 2340 522
rect 2322 6354 2340 6372
rect 2322 6372 2340 6390
rect 2322 6390 2340 6408
rect 2322 6408 2340 6426
rect 2322 6426 2340 6444
rect 2322 6444 2340 6462
rect 2322 6462 2340 6480
rect 2322 6480 2340 6498
rect 2322 6498 2340 6516
rect 2322 6516 2340 6534
rect 2322 6534 2340 6552
rect 2322 6552 2340 6570
rect 2322 6570 2340 6588
rect 2322 6588 2340 6606
rect 2322 6606 2340 6624
rect 2322 6624 2340 6642
rect 2322 6642 2340 6660
rect 2322 6660 2340 6678
rect 2322 6678 2340 6696
rect 2322 6696 2340 6714
rect 2322 6714 2340 6732
rect 2322 6732 2340 6750
rect 2322 6750 2340 6768
rect 2322 6768 2340 6786
rect 2322 6786 2340 6804
rect 2322 6804 2340 6822
rect 2322 6822 2340 6840
rect 2322 6840 2340 6858
rect 2322 6858 2340 6876
rect 2322 6876 2340 6894
rect 2322 6894 2340 6912
rect 2322 6912 2340 6930
rect 2322 6930 2340 6948
rect 2322 6948 2340 6966
rect 2322 6966 2340 6984
rect 2322 6984 2340 7002
rect 2322 7002 2340 7020
rect 2340 432 2358 450
rect 2340 450 2358 468
rect 2340 468 2358 486
rect 2340 486 2358 504
rect 2340 504 2358 522
rect 2340 522 2358 540
rect 2340 540 2358 558
rect 2340 558 2358 576
rect 2340 576 2358 594
rect 2340 594 2358 612
rect 2340 612 2358 630
rect 2340 6354 2358 6372
rect 2340 6372 2358 6390
rect 2340 6390 2358 6408
rect 2340 6408 2358 6426
rect 2340 6426 2358 6444
rect 2340 6444 2358 6462
rect 2340 6462 2358 6480
rect 2340 6480 2358 6498
rect 2340 6498 2358 6516
rect 2340 6516 2358 6534
rect 2340 6534 2358 6552
rect 2340 6552 2358 6570
rect 2340 6570 2358 6588
rect 2340 6588 2358 6606
rect 2340 6606 2358 6624
rect 2340 6624 2358 6642
rect 2340 6642 2358 6660
rect 2340 6660 2358 6678
rect 2340 6678 2358 6696
rect 2340 6696 2358 6714
rect 2340 6714 2358 6732
rect 2340 6732 2358 6750
rect 2340 6750 2358 6768
rect 2340 6768 2358 6786
rect 2340 6786 2358 6804
rect 2340 6804 2358 6822
rect 2340 6822 2358 6840
rect 2340 6840 2358 6858
rect 2340 6858 2358 6876
rect 2340 6876 2358 6894
rect 2340 6894 2358 6912
rect 2340 6912 2358 6930
rect 2340 6930 2358 6948
rect 2340 6948 2358 6966
rect 2340 6966 2358 6984
rect 2340 6984 2358 7002
rect 2340 7002 2358 7020
rect 2340 7020 2358 7038
rect 2358 468 2376 486
rect 2358 486 2376 504
rect 2358 504 2376 522
rect 2358 522 2376 540
rect 2358 540 2376 558
rect 2358 558 2376 576
rect 2358 576 2376 594
rect 2358 594 2376 612
rect 2358 612 2376 630
rect 2358 630 2376 648
rect 2358 648 2376 666
rect 2358 666 2376 684
rect 2358 684 2376 702
rect 2358 702 2376 720
rect 2358 6372 2376 6390
rect 2358 6390 2376 6408
rect 2358 6408 2376 6426
rect 2358 6426 2376 6444
rect 2358 6444 2376 6462
rect 2358 6462 2376 6480
rect 2358 6480 2376 6498
rect 2358 6498 2376 6516
rect 2358 6516 2376 6534
rect 2358 6534 2376 6552
rect 2358 6552 2376 6570
rect 2358 6570 2376 6588
rect 2358 6588 2376 6606
rect 2358 6606 2376 6624
rect 2358 6624 2376 6642
rect 2358 6642 2376 6660
rect 2358 6660 2376 6678
rect 2358 6678 2376 6696
rect 2358 6696 2376 6714
rect 2358 6714 2376 6732
rect 2358 6732 2376 6750
rect 2358 6750 2376 6768
rect 2358 6768 2376 6786
rect 2358 6786 2376 6804
rect 2358 6804 2376 6822
rect 2358 6822 2376 6840
rect 2358 6840 2376 6858
rect 2358 6858 2376 6876
rect 2358 6876 2376 6894
rect 2358 6894 2376 6912
rect 2358 6912 2376 6930
rect 2358 6930 2376 6948
rect 2358 6948 2376 6966
rect 2358 6966 2376 6984
rect 2358 6984 2376 7002
rect 2358 7002 2376 7020
rect 2358 7020 2376 7038
rect 2376 504 2394 522
rect 2376 522 2394 540
rect 2376 540 2394 558
rect 2376 558 2394 576
rect 2376 576 2394 594
rect 2376 594 2394 612
rect 2376 612 2394 630
rect 2376 630 2394 648
rect 2376 648 2394 666
rect 2376 666 2394 684
rect 2376 684 2394 702
rect 2376 702 2394 720
rect 2376 720 2394 738
rect 2376 738 2394 756
rect 2376 756 2394 774
rect 2376 774 2394 792
rect 2376 792 2394 810
rect 2376 6372 2394 6390
rect 2376 6390 2394 6408
rect 2376 6408 2394 6426
rect 2376 6426 2394 6444
rect 2376 6444 2394 6462
rect 2376 6462 2394 6480
rect 2376 6480 2394 6498
rect 2376 6498 2394 6516
rect 2376 6516 2394 6534
rect 2376 6534 2394 6552
rect 2376 6552 2394 6570
rect 2376 6570 2394 6588
rect 2376 6588 2394 6606
rect 2376 6606 2394 6624
rect 2376 6624 2394 6642
rect 2376 6642 2394 6660
rect 2376 6660 2394 6678
rect 2376 6678 2394 6696
rect 2376 6696 2394 6714
rect 2376 6714 2394 6732
rect 2376 6732 2394 6750
rect 2376 6750 2394 6768
rect 2376 6768 2394 6786
rect 2376 6786 2394 6804
rect 2376 6804 2394 6822
rect 2376 6822 2394 6840
rect 2376 6840 2394 6858
rect 2376 6858 2394 6876
rect 2376 6876 2394 6894
rect 2376 6894 2394 6912
rect 2376 6912 2394 6930
rect 2376 6930 2394 6948
rect 2376 6948 2394 6966
rect 2376 6966 2394 6984
rect 2376 6984 2394 7002
rect 2376 7002 2394 7020
rect 2376 7020 2394 7038
rect 2376 7038 2394 7056
rect 2394 540 2412 558
rect 2394 558 2412 576
rect 2394 576 2412 594
rect 2394 594 2412 612
rect 2394 612 2412 630
rect 2394 630 2412 648
rect 2394 648 2412 666
rect 2394 666 2412 684
rect 2394 684 2412 702
rect 2394 702 2412 720
rect 2394 720 2412 738
rect 2394 738 2412 756
rect 2394 756 2412 774
rect 2394 774 2412 792
rect 2394 792 2412 810
rect 2394 810 2412 828
rect 2394 828 2412 846
rect 2394 846 2412 864
rect 2394 864 2412 882
rect 2394 882 2412 900
rect 2394 6372 2412 6390
rect 2394 6390 2412 6408
rect 2394 6408 2412 6426
rect 2394 6426 2412 6444
rect 2394 6444 2412 6462
rect 2394 6462 2412 6480
rect 2394 6480 2412 6498
rect 2394 6498 2412 6516
rect 2394 6516 2412 6534
rect 2394 6534 2412 6552
rect 2394 6552 2412 6570
rect 2394 6570 2412 6588
rect 2394 6588 2412 6606
rect 2394 6606 2412 6624
rect 2394 6624 2412 6642
rect 2394 6642 2412 6660
rect 2394 6660 2412 6678
rect 2394 6678 2412 6696
rect 2394 6696 2412 6714
rect 2394 6714 2412 6732
rect 2394 6732 2412 6750
rect 2394 6750 2412 6768
rect 2394 6768 2412 6786
rect 2394 6786 2412 6804
rect 2394 6804 2412 6822
rect 2394 6822 2412 6840
rect 2394 6840 2412 6858
rect 2394 6858 2412 6876
rect 2394 6876 2412 6894
rect 2394 6894 2412 6912
rect 2394 6912 2412 6930
rect 2394 6930 2412 6948
rect 2394 6948 2412 6966
rect 2394 6966 2412 6984
rect 2394 6984 2412 7002
rect 2394 7002 2412 7020
rect 2394 7020 2412 7038
rect 2394 7038 2412 7056
rect 2412 576 2430 594
rect 2412 594 2430 612
rect 2412 612 2430 630
rect 2412 630 2430 648
rect 2412 648 2430 666
rect 2412 666 2430 684
rect 2412 684 2430 702
rect 2412 702 2430 720
rect 2412 720 2430 738
rect 2412 738 2430 756
rect 2412 756 2430 774
rect 2412 774 2430 792
rect 2412 792 2430 810
rect 2412 810 2430 828
rect 2412 828 2430 846
rect 2412 846 2430 864
rect 2412 864 2430 882
rect 2412 882 2430 900
rect 2412 900 2430 918
rect 2412 918 2430 936
rect 2412 936 2430 954
rect 2412 954 2430 972
rect 2412 972 2430 990
rect 2412 6390 2430 6408
rect 2412 6408 2430 6426
rect 2412 6426 2430 6444
rect 2412 6444 2430 6462
rect 2412 6462 2430 6480
rect 2412 6480 2430 6498
rect 2412 6498 2430 6516
rect 2412 6516 2430 6534
rect 2412 6534 2430 6552
rect 2412 6552 2430 6570
rect 2412 6570 2430 6588
rect 2412 6588 2430 6606
rect 2412 6606 2430 6624
rect 2412 6624 2430 6642
rect 2412 6642 2430 6660
rect 2412 6660 2430 6678
rect 2412 6678 2430 6696
rect 2412 6696 2430 6714
rect 2412 6714 2430 6732
rect 2412 6732 2430 6750
rect 2412 6750 2430 6768
rect 2412 6768 2430 6786
rect 2412 6786 2430 6804
rect 2412 6804 2430 6822
rect 2412 6822 2430 6840
rect 2412 6840 2430 6858
rect 2412 6858 2430 6876
rect 2412 6876 2430 6894
rect 2412 6894 2430 6912
rect 2412 6912 2430 6930
rect 2412 6930 2430 6948
rect 2412 6948 2430 6966
rect 2412 6966 2430 6984
rect 2412 6984 2430 7002
rect 2412 7002 2430 7020
rect 2412 7020 2430 7038
rect 2412 7038 2430 7056
rect 2430 612 2448 630
rect 2430 630 2448 648
rect 2430 648 2448 666
rect 2430 666 2448 684
rect 2430 684 2448 702
rect 2430 702 2448 720
rect 2430 720 2448 738
rect 2430 738 2448 756
rect 2430 756 2448 774
rect 2430 774 2448 792
rect 2430 792 2448 810
rect 2430 810 2448 828
rect 2430 828 2448 846
rect 2430 846 2448 864
rect 2430 864 2448 882
rect 2430 882 2448 900
rect 2430 900 2448 918
rect 2430 918 2448 936
rect 2430 936 2448 954
rect 2430 954 2448 972
rect 2430 972 2448 990
rect 2430 990 2448 1008
rect 2430 1008 2448 1026
rect 2430 1026 2448 1044
rect 2430 1044 2448 1062
rect 2430 1062 2448 1080
rect 2430 1080 2448 1098
rect 2430 6390 2448 6408
rect 2430 6408 2448 6426
rect 2430 6426 2448 6444
rect 2430 6444 2448 6462
rect 2430 6462 2448 6480
rect 2430 6480 2448 6498
rect 2430 6498 2448 6516
rect 2430 6516 2448 6534
rect 2430 6534 2448 6552
rect 2430 6552 2448 6570
rect 2430 6570 2448 6588
rect 2430 6588 2448 6606
rect 2430 6606 2448 6624
rect 2430 6624 2448 6642
rect 2430 6642 2448 6660
rect 2430 6660 2448 6678
rect 2430 6678 2448 6696
rect 2430 6696 2448 6714
rect 2430 6714 2448 6732
rect 2430 6732 2448 6750
rect 2430 6750 2448 6768
rect 2430 6768 2448 6786
rect 2430 6786 2448 6804
rect 2430 6804 2448 6822
rect 2430 6822 2448 6840
rect 2430 6840 2448 6858
rect 2430 6858 2448 6876
rect 2430 6876 2448 6894
rect 2430 6894 2448 6912
rect 2430 6912 2448 6930
rect 2430 6930 2448 6948
rect 2430 6948 2448 6966
rect 2430 6966 2448 6984
rect 2430 6984 2448 7002
rect 2430 7002 2448 7020
rect 2430 7020 2448 7038
rect 2430 7038 2448 7056
rect 2430 7056 2448 7074
rect 2448 666 2466 684
rect 2448 684 2466 702
rect 2448 702 2466 720
rect 2448 720 2466 738
rect 2448 738 2466 756
rect 2448 756 2466 774
rect 2448 774 2466 792
rect 2448 792 2466 810
rect 2448 810 2466 828
rect 2448 828 2466 846
rect 2448 846 2466 864
rect 2448 864 2466 882
rect 2448 882 2466 900
rect 2448 900 2466 918
rect 2448 918 2466 936
rect 2448 936 2466 954
rect 2448 954 2466 972
rect 2448 972 2466 990
rect 2448 990 2466 1008
rect 2448 1008 2466 1026
rect 2448 1026 2466 1044
rect 2448 1044 2466 1062
rect 2448 1062 2466 1080
rect 2448 1080 2466 1098
rect 2448 1098 2466 1116
rect 2448 1116 2466 1134
rect 2448 1134 2466 1152
rect 2448 1152 2466 1170
rect 2448 1170 2466 1188
rect 2448 6408 2466 6426
rect 2448 6426 2466 6444
rect 2448 6444 2466 6462
rect 2448 6462 2466 6480
rect 2448 6480 2466 6498
rect 2448 6498 2466 6516
rect 2448 6516 2466 6534
rect 2448 6534 2466 6552
rect 2448 6552 2466 6570
rect 2448 6570 2466 6588
rect 2448 6588 2466 6606
rect 2448 6606 2466 6624
rect 2448 6624 2466 6642
rect 2448 6642 2466 6660
rect 2448 6660 2466 6678
rect 2448 6678 2466 6696
rect 2448 6696 2466 6714
rect 2448 6714 2466 6732
rect 2448 6732 2466 6750
rect 2448 6750 2466 6768
rect 2448 6768 2466 6786
rect 2448 6786 2466 6804
rect 2448 6804 2466 6822
rect 2448 6822 2466 6840
rect 2448 6840 2466 6858
rect 2448 6858 2466 6876
rect 2448 6876 2466 6894
rect 2448 6894 2466 6912
rect 2448 6912 2466 6930
rect 2448 6930 2466 6948
rect 2448 6948 2466 6966
rect 2448 6966 2466 6984
rect 2448 6984 2466 7002
rect 2448 7002 2466 7020
rect 2448 7020 2466 7038
rect 2448 7038 2466 7056
rect 2448 7056 2466 7074
rect 2466 702 2484 720
rect 2466 720 2484 738
rect 2466 738 2484 756
rect 2466 756 2484 774
rect 2466 774 2484 792
rect 2466 792 2484 810
rect 2466 810 2484 828
rect 2466 828 2484 846
rect 2466 846 2484 864
rect 2466 864 2484 882
rect 2466 882 2484 900
rect 2466 900 2484 918
rect 2466 918 2484 936
rect 2466 936 2484 954
rect 2466 954 2484 972
rect 2466 972 2484 990
rect 2466 990 2484 1008
rect 2466 1008 2484 1026
rect 2466 1026 2484 1044
rect 2466 1044 2484 1062
rect 2466 1062 2484 1080
rect 2466 1080 2484 1098
rect 2466 1098 2484 1116
rect 2466 1116 2484 1134
rect 2466 1134 2484 1152
rect 2466 1152 2484 1170
rect 2466 1170 2484 1188
rect 2466 1188 2484 1206
rect 2466 1206 2484 1224
rect 2466 1224 2484 1242
rect 2466 1242 2484 1260
rect 2466 6408 2484 6426
rect 2466 6426 2484 6444
rect 2466 6444 2484 6462
rect 2466 6462 2484 6480
rect 2466 6480 2484 6498
rect 2466 6498 2484 6516
rect 2466 6516 2484 6534
rect 2466 6534 2484 6552
rect 2466 6552 2484 6570
rect 2466 6570 2484 6588
rect 2466 6588 2484 6606
rect 2466 6606 2484 6624
rect 2466 6624 2484 6642
rect 2466 6642 2484 6660
rect 2466 6660 2484 6678
rect 2466 6678 2484 6696
rect 2466 6696 2484 6714
rect 2466 6714 2484 6732
rect 2466 6732 2484 6750
rect 2466 6750 2484 6768
rect 2466 6768 2484 6786
rect 2466 6786 2484 6804
rect 2466 6804 2484 6822
rect 2466 6822 2484 6840
rect 2466 6840 2484 6858
rect 2466 6858 2484 6876
rect 2466 6876 2484 6894
rect 2466 6894 2484 6912
rect 2466 6912 2484 6930
rect 2466 6930 2484 6948
rect 2466 6948 2484 6966
rect 2466 6966 2484 6984
rect 2466 6984 2484 7002
rect 2466 7002 2484 7020
rect 2466 7020 2484 7038
rect 2466 7038 2484 7056
rect 2466 7056 2484 7074
rect 2484 216 2502 234
rect 2484 234 2502 252
rect 2484 738 2502 756
rect 2484 756 2502 774
rect 2484 774 2502 792
rect 2484 792 2502 810
rect 2484 810 2502 828
rect 2484 828 2502 846
rect 2484 846 2502 864
rect 2484 864 2502 882
rect 2484 882 2502 900
rect 2484 900 2502 918
rect 2484 918 2502 936
rect 2484 936 2502 954
rect 2484 954 2502 972
rect 2484 972 2502 990
rect 2484 990 2502 1008
rect 2484 1008 2502 1026
rect 2484 1026 2502 1044
rect 2484 1044 2502 1062
rect 2484 1062 2502 1080
rect 2484 1080 2502 1098
rect 2484 1098 2502 1116
rect 2484 1116 2502 1134
rect 2484 1134 2502 1152
rect 2484 1152 2502 1170
rect 2484 1170 2502 1188
rect 2484 1188 2502 1206
rect 2484 1206 2502 1224
rect 2484 1224 2502 1242
rect 2484 1242 2502 1260
rect 2484 1260 2502 1278
rect 2484 1278 2502 1296
rect 2484 1296 2502 1314
rect 2484 1314 2502 1332
rect 2484 1332 2502 1350
rect 2484 6426 2502 6444
rect 2484 6444 2502 6462
rect 2484 6462 2502 6480
rect 2484 6480 2502 6498
rect 2484 6498 2502 6516
rect 2484 6516 2502 6534
rect 2484 6534 2502 6552
rect 2484 6552 2502 6570
rect 2484 6570 2502 6588
rect 2484 6588 2502 6606
rect 2484 6606 2502 6624
rect 2484 6624 2502 6642
rect 2484 6642 2502 6660
rect 2484 6660 2502 6678
rect 2484 6678 2502 6696
rect 2484 6696 2502 6714
rect 2484 6714 2502 6732
rect 2484 6732 2502 6750
rect 2484 6750 2502 6768
rect 2484 6768 2502 6786
rect 2484 6786 2502 6804
rect 2484 6804 2502 6822
rect 2484 6822 2502 6840
rect 2484 6840 2502 6858
rect 2484 6858 2502 6876
rect 2484 6876 2502 6894
rect 2484 6894 2502 6912
rect 2484 6912 2502 6930
rect 2484 6930 2502 6948
rect 2484 6948 2502 6966
rect 2484 6966 2502 6984
rect 2484 6984 2502 7002
rect 2484 7002 2502 7020
rect 2484 7020 2502 7038
rect 2484 7038 2502 7056
rect 2484 7056 2502 7074
rect 2484 7074 2502 7092
rect 2502 216 2520 234
rect 2502 234 2520 252
rect 2502 252 2520 270
rect 2502 270 2520 288
rect 2502 774 2520 792
rect 2502 792 2520 810
rect 2502 810 2520 828
rect 2502 828 2520 846
rect 2502 846 2520 864
rect 2502 864 2520 882
rect 2502 882 2520 900
rect 2502 900 2520 918
rect 2502 918 2520 936
rect 2502 936 2520 954
rect 2502 954 2520 972
rect 2502 972 2520 990
rect 2502 990 2520 1008
rect 2502 1008 2520 1026
rect 2502 1026 2520 1044
rect 2502 1044 2520 1062
rect 2502 1062 2520 1080
rect 2502 1080 2520 1098
rect 2502 1098 2520 1116
rect 2502 1116 2520 1134
rect 2502 1134 2520 1152
rect 2502 1152 2520 1170
rect 2502 1170 2520 1188
rect 2502 1188 2520 1206
rect 2502 1206 2520 1224
rect 2502 1224 2520 1242
rect 2502 1242 2520 1260
rect 2502 1260 2520 1278
rect 2502 1278 2520 1296
rect 2502 1296 2520 1314
rect 2502 1314 2520 1332
rect 2502 1332 2520 1350
rect 2502 1350 2520 1368
rect 2502 1368 2520 1386
rect 2502 1386 2520 1404
rect 2502 1404 2520 1422
rect 2502 1422 2520 1440
rect 2502 6426 2520 6444
rect 2502 6444 2520 6462
rect 2502 6462 2520 6480
rect 2502 6480 2520 6498
rect 2502 6498 2520 6516
rect 2502 6516 2520 6534
rect 2502 6534 2520 6552
rect 2502 6552 2520 6570
rect 2502 6570 2520 6588
rect 2502 6588 2520 6606
rect 2502 6606 2520 6624
rect 2502 6624 2520 6642
rect 2502 6642 2520 6660
rect 2502 6660 2520 6678
rect 2502 6678 2520 6696
rect 2502 6696 2520 6714
rect 2502 6714 2520 6732
rect 2502 6732 2520 6750
rect 2502 6750 2520 6768
rect 2502 6768 2520 6786
rect 2502 6786 2520 6804
rect 2502 6804 2520 6822
rect 2502 6822 2520 6840
rect 2502 6840 2520 6858
rect 2502 6858 2520 6876
rect 2502 6876 2520 6894
rect 2502 6894 2520 6912
rect 2502 6912 2520 6930
rect 2502 6930 2520 6948
rect 2502 6948 2520 6966
rect 2502 6966 2520 6984
rect 2502 6984 2520 7002
rect 2502 7002 2520 7020
rect 2502 7020 2520 7038
rect 2502 7038 2520 7056
rect 2502 7056 2520 7074
rect 2502 7074 2520 7092
rect 2520 234 2538 252
rect 2520 252 2538 270
rect 2520 270 2538 288
rect 2520 288 2538 306
rect 2520 306 2538 324
rect 2520 810 2538 828
rect 2520 828 2538 846
rect 2520 846 2538 864
rect 2520 864 2538 882
rect 2520 882 2538 900
rect 2520 900 2538 918
rect 2520 918 2538 936
rect 2520 936 2538 954
rect 2520 954 2538 972
rect 2520 972 2538 990
rect 2520 990 2538 1008
rect 2520 1008 2538 1026
rect 2520 1026 2538 1044
rect 2520 1044 2538 1062
rect 2520 1062 2538 1080
rect 2520 1080 2538 1098
rect 2520 1098 2538 1116
rect 2520 1116 2538 1134
rect 2520 1134 2538 1152
rect 2520 1152 2538 1170
rect 2520 1170 2538 1188
rect 2520 1188 2538 1206
rect 2520 1206 2538 1224
rect 2520 1224 2538 1242
rect 2520 1242 2538 1260
rect 2520 1260 2538 1278
rect 2520 1278 2538 1296
rect 2520 1296 2538 1314
rect 2520 1314 2538 1332
rect 2520 1332 2538 1350
rect 2520 1350 2538 1368
rect 2520 1368 2538 1386
rect 2520 1386 2538 1404
rect 2520 1404 2538 1422
rect 2520 1422 2538 1440
rect 2520 1440 2538 1458
rect 2520 1458 2538 1476
rect 2520 1476 2538 1494
rect 2520 1494 2538 1512
rect 2520 1512 2538 1530
rect 2520 6426 2538 6444
rect 2520 6444 2538 6462
rect 2520 6462 2538 6480
rect 2520 6480 2538 6498
rect 2520 6498 2538 6516
rect 2520 6516 2538 6534
rect 2520 6534 2538 6552
rect 2520 6552 2538 6570
rect 2520 6570 2538 6588
rect 2520 6588 2538 6606
rect 2520 6606 2538 6624
rect 2520 6624 2538 6642
rect 2520 6642 2538 6660
rect 2520 6660 2538 6678
rect 2520 6678 2538 6696
rect 2520 6696 2538 6714
rect 2520 6714 2538 6732
rect 2520 6732 2538 6750
rect 2520 6750 2538 6768
rect 2520 6768 2538 6786
rect 2520 6786 2538 6804
rect 2520 6804 2538 6822
rect 2520 6822 2538 6840
rect 2520 6840 2538 6858
rect 2520 6858 2538 6876
rect 2520 6876 2538 6894
rect 2520 6894 2538 6912
rect 2520 6912 2538 6930
rect 2520 6930 2538 6948
rect 2520 6948 2538 6966
rect 2520 6966 2538 6984
rect 2520 6984 2538 7002
rect 2520 7002 2538 7020
rect 2520 7020 2538 7038
rect 2520 7038 2538 7056
rect 2520 7056 2538 7074
rect 2520 7074 2538 7092
rect 2538 252 2556 270
rect 2538 270 2556 288
rect 2538 288 2556 306
rect 2538 306 2556 324
rect 2538 324 2556 342
rect 2538 342 2556 360
rect 2538 846 2556 864
rect 2538 864 2556 882
rect 2538 882 2556 900
rect 2538 900 2556 918
rect 2538 918 2556 936
rect 2538 936 2556 954
rect 2538 954 2556 972
rect 2538 972 2556 990
rect 2538 990 2556 1008
rect 2538 1008 2556 1026
rect 2538 1026 2556 1044
rect 2538 1044 2556 1062
rect 2538 1062 2556 1080
rect 2538 1080 2556 1098
rect 2538 1098 2556 1116
rect 2538 1116 2556 1134
rect 2538 1134 2556 1152
rect 2538 1152 2556 1170
rect 2538 1170 2556 1188
rect 2538 1188 2556 1206
rect 2538 1206 2556 1224
rect 2538 1224 2556 1242
rect 2538 1242 2556 1260
rect 2538 1260 2556 1278
rect 2538 1278 2556 1296
rect 2538 1296 2556 1314
rect 2538 1314 2556 1332
rect 2538 1332 2556 1350
rect 2538 1350 2556 1368
rect 2538 1368 2556 1386
rect 2538 1386 2556 1404
rect 2538 1404 2556 1422
rect 2538 1422 2556 1440
rect 2538 1440 2556 1458
rect 2538 1458 2556 1476
rect 2538 1476 2556 1494
rect 2538 1494 2556 1512
rect 2538 1512 2556 1530
rect 2538 1530 2556 1548
rect 2538 1548 2556 1566
rect 2538 1566 2556 1584
rect 2538 1584 2556 1602
rect 2538 6444 2556 6462
rect 2538 6462 2556 6480
rect 2538 6480 2556 6498
rect 2538 6498 2556 6516
rect 2538 6516 2556 6534
rect 2538 6534 2556 6552
rect 2538 6552 2556 6570
rect 2538 6570 2556 6588
rect 2538 6588 2556 6606
rect 2538 6606 2556 6624
rect 2538 6624 2556 6642
rect 2538 6642 2556 6660
rect 2538 6660 2556 6678
rect 2538 6678 2556 6696
rect 2538 6696 2556 6714
rect 2538 6714 2556 6732
rect 2538 6732 2556 6750
rect 2538 6750 2556 6768
rect 2538 6768 2556 6786
rect 2538 6786 2556 6804
rect 2538 6804 2556 6822
rect 2538 6822 2556 6840
rect 2538 6840 2556 6858
rect 2538 6858 2556 6876
rect 2538 6876 2556 6894
rect 2538 6894 2556 6912
rect 2538 6912 2556 6930
rect 2538 6930 2556 6948
rect 2538 6948 2556 6966
rect 2538 6966 2556 6984
rect 2538 6984 2556 7002
rect 2538 7002 2556 7020
rect 2538 7020 2556 7038
rect 2538 7038 2556 7056
rect 2538 7056 2556 7074
rect 2538 7074 2556 7092
rect 2538 7092 2556 7110
rect 2556 252 2574 270
rect 2556 270 2574 288
rect 2556 288 2574 306
rect 2556 306 2574 324
rect 2556 324 2574 342
rect 2556 342 2574 360
rect 2556 360 2574 378
rect 2556 378 2574 396
rect 2556 882 2574 900
rect 2556 900 2574 918
rect 2556 918 2574 936
rect 2556 936 2574 954
rect 2556 954 2574 972
rect 2556 972 2574 990
rect 2556 990 2574 1008
rect 2556 1008 2574 1026
rect 2556 1026 2574 1044
rect 2556 1044 2574 1062
rect 2556 1062 2574 1080
rect 2556 1080 2574 1098
rect 2556 1098 2574 1116
rect 2556 1116 2574 1134
rect 2556 1134 2574 1152
rect 2556 1152 2574 1170
rect 2556 1170 2574 1188
rect 2556 1188 2574 1206
rect 2556 1206 2574 1224
rect 2556 1224 2574 1242
rect 2556 1242 2574 1260
rect 2556 1260 2574 1278
rect 2556 1278 2574 1296
rect 2556 1296 2574 1314
rect 2556 1314 2574 1332
rect 2556 1332 2574 1350
rect 2556 1350 2574 1368
rect 2556 1368 2574 1386
rect 2556 1386 2574 1404
rect 2556 1404 2574 1422
rect 2556 1422 2574 1440
rect 2556 1440 2574 1458
rect 2556 1458 2574 1476
rect 2556 1476 2574 1494
rect 2556 1494 2574 1512
rect 2556 1512 2574 1530
rect 2556 1530 2574 1548
rect 2556 1548 2574 1566
rect 2556 1566 2574 1584
rect 2556 1584 2574 1602
rect 2556 1602 2574 1620
rect 2556 1620 2574 1638
rect 2556 1638 2574 1656
rect 2556 1656 2574 1674
rect 2556 1674 2574 1692
rect 2556 6444 2574 6462
rect 2556 6462 2574 6480
rect 2556 6480 2574 6498
rect 2556 6498 2574 6516
rect 2556 6516 2574 6534
rect 2556 6534 2574 6552
rect 2556 6552 2574 6570
rect 2556 6570 2574 6588
rect 2556 6588 2574 6606
rect 2556 6606 2574 6624
rect 2556 6624 2574 6642
rect 2556 6642 2574 6660
rect 2556 6660 2574 6678
rect 2556 6678 2574 6696
rect 2556 6696 2574 6714
rect 2556 6714 2574 6732
rect 2556 6732 2574 6750
rect 2556 6750 2574 6768
rect 2556 6768 2574 6786
rect 2556 6786 2574 6804
rect 2556 6804 2574 6822
rect 2556 6822 2574 6840
rect 2556 6840 2574 6858
rect 2556 6858 2574 6876
rect 2556 6876 2574 6894
rect 2556 6894 2574 6912
rect 2556 6912 2574 6930
rect 2556 6930 2574 6948
rect 2556 6948 2574 6966
rect 2556 6966 2574 6984
rect 2556 6984 2574 7002
rect 2556 7002 2574 7020
rect 2556 7020 2574 7038
rect 2556 7038 2574 7056
rect 2556 7056 2574 7074
rect 2556 7074 2574 7092
rect 2556 7092 2574 7110
rect 2574 270 2592 288
rect 2574 288 2592 306
rect 2574 306 2592 324
rect 2574 324 2592 342
rect 2574 342 2592 360
rect 2574 360 2592 378
rect 2574 378 2592 396
rect 2574 396 2592 414
rect 2574 414 2592 432
rect 2574 918 2592 936
rect 2574 936 2592 954
rect 2574 954 2592 972
rect 2574 972 2592 990
rect 2574 990 2592 1008
rect 2574 1008 2592 1026
rect 2574 1026 2592 1044
rect 2574 1044 2592 1062
rect 2574 1062 2592 1080
rect 2574 1080 2592 1098
rect 2574 1098 2592 1116
rect 2574 1116 2592 1134
rect 2574 1134 2592 1152
rect 2574 1152 2592 1170
rect 2574 1170 2592 1188
rect 2574 1188 2592 1206
rect 2574 1206 2592 1224
rect 2574 1224 2592 1242
rect 2574 1242 2592 1260
rect 2574 1260 2592 1278
rect 2574 1278 2592 1296
rect 2574 1296 2592 1314
rect 2574 1314 2592 1332
rect 2574 1332 2592 1350
rect 2574 1350 2592 1368
rect 2574 1368 2592 1386
rect 2574 1386 2592 1404
rect 2574 1404 2592 1422
rect 2574 1422 2592 1440
rect 2574 1440 2592 1458
rect 2574 1458 2592 1476
rect 2574 1476 2592 1494
rect 2574 1494 2592 1512
rect 2574 1512 2592 1530
rect 2574 1530 2592 1548
rect 2574 1548 2592 1566
rect 2574 1566 2592 1584
rect 2574 1584 2592 1602
rect 2574 1602 2592 1620
rect 2574 1620 2592 1638
rect 2574 1638 2592 1656
rect 2574 1656 2592 1674
rect 2574 1674 2592 1692
rect 2574 1692 2592 1710
rect 2574 1710 2592 1728
rect 2574 1728 2592 1746
rect 2574 1746 2592 1764
rect 2574 6462 2592 6480
rect 2574 6480 2592 6498
rect 2574 6498 2592 6516
rect 2574 6516 2592 6534
rect 2574 6534 2592 6552
rect 2574 6552 2592 6570
rect 2574 6570 2592 6588
rect 2574 6588 2592 6606
rect 2574 6606 2592 6624
rect 2574 6624 2592 6642
rect 2574 6642 2592 6660
rect 2574 6660 2592 6678
rect 2574 6678 2592 6696
rect 2574 6696 2592 6714
rect 2574 6714 2592 6732
rect 2574 6732 2592 6750
rect 2574 6750 2592 6768
rect 2574 6768 2592 6786
rect 2574 6786 2592 6804
rect 2574 6804 2592 6822
rect 2574 6822 2592 6840
rect 2574 6840 2592 6858
rect 2574 6858 2592 6876
rect 2574 6876 2592 6894
rect 2574 6894 2592 6912
rect 2574 6912 2592 6930
rect 2574 6930 2592 6948
rect 2574 6948 2592 6966
rect 2574 6966 2592 6984
rect 2574 6984 2592 7002
rect 2574 7002 2592 7020
rect 2574 7020 2592 7038
rect 2574 7038 2592 7056
rect 2574 7056 2592 7074
rect 2574 7074 2592 7092
rect 2574 7092 2592 7110
rect 2592 270 2610 288
rect 2592 288 2610 306
rect 2592 306 2610 324
rect 2592 324 2610 342
rect 2592 342 2610 360
rect 2592 360 2610 378
rect 2592 378 2610 396
rect 2592 396 2610 414
rect 2592 414 2610 432
rect 2592 432 2610 450
rect 2592 954 2610 972
rect 2592 972 2610 990
rect 2592 990 2610 1008
rect 2592 1008 2610 1026
rect 2592 1026 2610 1044
rect 2592 1044 2610 1062
rect 2592 1062 2610 1080
rect 2592 1080 2610 1098
rect 2592 1098 2610 1116
rect 2592 1116 2610 1134
rect 2592 1134 2610 1152
rect 2592 1152 2610 1170
rect 2592 1170 2610 1188
rect 2592 1188 2610 1206
rect 2592 1206 2610 1224
rect 2592 1224 2610 1242
rect 2592 1242 2610 1260
rect 2592 1260 2610 1278
rect 2592 1278 2610 1296
rect 2592 1296 2610 1314
rect 2592 1314 2610 1332
rect 2592 1332 2610 1350
rect 2592 1350 2610 1368
rect 2592 1368 2610 1386
rect 2592 1386 2610 1404
rect 2592 1404 2610 1422
rect 2592 1422 2610 1440
rect 2592 1440 2610 1458
rect 2592 1458 2610 1476
rect 2592 1476 2610 1494
rect 2592 1494 2610 1512
rect 2592 1512 2610 1530
rect 2592 1530 2610 1548
rect 2592 1548 2610 1566
rect 2592 1566 2610 1584
rect 2592 1584 2610 1602
rect 2592 1602 2610 1620
rect 2592 1620 2610 1638
rect 2592 1638 2610 1656
rect 2592 1656 2610 1674
rect 2592 1674 2610 1692
rect 2592 1692 2610 1710
rect 2592 1710 2610 1728
rect 2592 1728 2610 1746
rect 2592 1746 2610 1764
rect 2592 1764 2610 1782
rect 2592 1782 2610 1800
rect 2592 1800 2610 1818
rect 2592 1818 2610 1836
rect 2592 1836 2610 1854
rect 2592 6462 2610 6480
rect 2592 6480 2610 6498
rect 2592 6498 2610 6516
rect 2592 6516 2610 6534
rect 2592 6534 2610 6552
rect 2592 6552 2610 6570
rect 2592 6570 2610 6588
rect 2592 6588 2610 6606
rect 2592 6606 2610 6624
rect 2592 6624 2610 6642
rect 2592 6642 2610 6660
rect 2592 6660 2610 6678
rect 2592 6678 2610 6696
rect 2592 6696 2610 6714
rect 2592 6714 2610 6732
rect 2592 6732 2610 6750
rect 2592 6750 2610 6768
rect 2592 6768 2610 6786
rect 2592 6786 2610 6804
rect 2592 6804 2610 6822
rect 2592 6822 2610 6840
rect 2592 6840 2610 6858
rect 2592 6858 2610 6876
rect 2592 6876 2610 6894
rect 2592 6894 2610 6912
rect 2592 6912 2610 6930
rect 2592 6930 2610 6948
rect 2592 6948 2610 6966
rect 2592 6966 2610 6984
rect 2592 6984 2610 7002
rect 2592 7002 2610 7020
rect 2592 7020 2610 7038
rect 2592 7038 2610 7056
rect 2592 7056 2610 7074
rect 2592 7074 2610 7092
rect 2592 7092 2610 7110
rect 2592 7110 2610 7128
rect 2610 288 2628 306
rect 2610 306 2628 324
rect 2610 324 2628 342
rect 2610 342 2628 360
rect 2610 360 2628 378
rect 2610 378 2628 396
rect 2610 396 2628 414
rect 2610 414 2628 432
rect 2610 432 2628 450
rect 2610 450 2628 468
rect 2610 468 2628 486
rect 2610 990 2628 1008
rect 2610 1008 2628 1026
rect 2610 1026 2628 1044
rect 2610 1044 2628 1062
rect 2610 1062 2628 1080
rect 2610 1080 2628 1098
rect 2610 1098 2628 1116
rect 2610 1116 2628 1134
rect 2610 1134 2628 1152
rect 2610 1152 2628 1170
rect 2610 1170 2628 1188
rect 2610 1188 2628 1206
rect 2610 1206 2628 1224
rect 2610 1224 2628 1242
rect 2610 1242 2628 1260
rect 2610 1260 2628 1278
rect 2610 1278 2628 1296
rect 2610 1296 2628 1314
rect 2610 1314 2628 1332
rect 2610 1332 2628 1350
rect 2610 1350 2628 1368
rect 2610 1368 2628 1386
rect 2610 1386 2628 1404
rect 2610 1404 2628 1422
rect 2610 1422 2628 1440
rect 2610 1440 2628 1458
rect 2610 1458 2628 1476
rect 2610 1476 2628 1494
rect 2610 1494 2628 1512
rect 2610 1512 2628 1530
rect 2610 1530 2628 1548
rect 2610 1548 2628 1566
rect 2610 1566 2628 1584
rect 2610 1584 2628 1602
rect 2610 1602 2628 1620
rect 2610 1620 2628 1638
rect 2610 1638 2628 1656
rect 2610 1656 2628 1674
rect 2610 1674 2628 1692
rect 2610 1692 2628 1710
rect 2610 1710 2628 1728
rect 2610 1728 2628 1746
rect 2610 1746 2628 1764
rect 2610 1764 2628 1782
rect 2610 1782 2628 1800
rect 2610 1800 2628 1818
rect 2610 1818 2628 1836
rect 2610 1836 2628 1854
rect 2610 1854 2628 1872
rect 2610 1872 2628 1890
rect 2610 1890 2628 1908
rect 2610 1908 2628 1926
rect 2610 6462 2628 6480
rect 2610 6480 2628 6498
rect 2610 6498 2628 6516
rect 2610 6516 2628 6534
rect 2610 6534 2628 6552
rect 2610 6552 2628 6570
rect 2610 6570 2628 6588
rect 2610 6588 2628 6606
rect 2610 6606 2628 6624
rect 2610 6624 2628 6642
rect 2610 6642 2628 6660
rect 2610 6660 2628 6678
rect 2610 6678 2628 6696
rect 2610 6696 2628 6714
rect 2610 6714 2628 6732
rect 2610 6732 2628 6750
rect 2610 6750 2628 6768
rect 2610 6768 2628 6786
rect 2610 6786 2628 6804
rect 2610 6804 2628 6822
rect 2610 6822 2628 6840
rect 2610 6840 2628 6858
rect 2610 6858 2628 6876
rect 2610 6876 2628 6894
rect 2610 6894 2628 6912
rect 2610 6912 2628 6930
rect 2610 6930 2628 6948
rect 2610 6948 2628 6966
rect 2610 6966 2628 6984
rect 2610 6984 2628 7002
rect 2610 7002 2628 7020
rect 2610 7020 2628 7038
rect 2610 7038 2628 7056
rect 2610 7056 2628 7074
rect 2610 7074 2628 7092
rect 2610 7092 2628 7110
rect 2610 7110 2628 7128
rect 2628 306 2646 324
rect 2628 324 2646 342
rect 2628 342 2646 360
rect 2628 360 2646 378
rect 2628 378 2646 396
rect 2628 396 2646 414
rect 2628 414 2646 432
rect 2628 432 2646 450
rect 2628 450 2646 468
rect 2628 468 2646 486
rect 2628 486 2646 504
rect 2628 1026 2646 1044
rect 2628 1044 2646 1062
rect 2628 1062 2646 1080
rect 2628 1080 2646 1098
rect 2628 1098 2646 1116
rect 2628 1116 2646 1134
rect 2628 1134 2646 1152
rect 2628 1152 2646 1170
rect 2628 1170 2646 1188
rect 2628 1188 2646 1206
rect 2628 1206 2646 1224
rect 2628 1224 2646 1242
rect 2628 1242 2646 1260
rect 2628 1260 2646 1278
rect 2628 1278 2646 1296
rect 2628 1296 2646 1314
rect 2628 1314 2646 1332
rect 2628 1332 2646 1350
rect 2628 1350 2646 1368
rect 2628 1368 2646 1386
rect 2628 1386 2646 1404
rect 2628 1404 2646 1422
rect 2628 1422 2646 1440
rect 2628 1440 2646 1458
rect 2628 1458 2646 1476
rect 2628 1476 2646 1494
rect 2628 1494 2646 1512
rect 2628 1512 2646 1530
rect 2628 1530 2646 1548
rect 2628 1548 2646 1566
rect 2628 1566 2646 1584
rect 2628 1584 2646 1602
rect 2628 1602 2646 1620
rect 2628 1620 2646 1638
rect 2628 1638 2646 1656
rect 2628 1656 2646 1674
rect 2628 1674 2646 1692
rect 2628 1692 2646 1710
rect 2628 1710 2646 1728
rect 2628 1728 2646 1746
rect 2628 1746 2646 1764
rect 2628 1764 2646 1782
rect 2628 1782 2646 1800
rect 2628 1800 2646 1818
rect 2628 1818 2646 1836
rect 2628 1836 2646 1854
rect 2628 1854 2646 1872
rect 2628 1872 2646 1890
rect 2628 1890 2646 1908
rect 2628 1908 2646 1926
rect 2628 1926 2646 1944
rect 2628 1944 2646 1962
rect 2628 1962 2646 1980
rect 2628 1980 2646 1998
rect 2628 6480 2646 6498
rect 2628 6498 2646 6516
rect 2628 6516 2646 6534
rect 2628 6534 2646 6552
rect 2628 6552 2646 6570
rect 2628 6570 2646 6588
rect 2628 6588 2646 6606
rect 2628 6606 2646 6624
rect 2628 6624 2646 6642
rect 2628 6642 2646 6660
rect 2628 6660 2646 6678
rect 2628 6678 2646 6696
rect 2628 6696 2646 6714
rect 2628 6714 2646 6732
rect 2628 6732 2646 6750
rect 2628 6750 2646 6768
rect 2628 6768 2646 6786
rect 2628 6786 2646 6804
rect 2628 6804 2646 6822
rect 2628 6822 2646 6840
rect 2628 6840 2646 6858
rect 2628 6858 2646 6876
rect 2628 6876 2646 6894
rect 2628 6894 2646 6912
rect 2628 6912 2646 6930
rect 2628 6930 2646 6948
rect 2628 6948 2646 6966
rect 2628 6966 2646 6984
rect 2628 6984 2646 7002
rect 2628 7002 2646 7020
rect 2628 7020 2646 7038
rect 2628 7038 2646 7056
rect 2628 7056 2646 7074
rect 2628 7074 2646 7092
rect 2628 7092 2646 7110
rect 2628 7110 2646 7128
rect 2646 306 2664 324
rect 2646 324 2664 342
rect 2646 342 2664 360
rect 2646 360 2664 378
rect 2646 378 2664 396
rect 2646 396 2664 414
rect 2646 414 2664 432
rect 2646 432 2664 450
rect 2646 450 2664 468
rect 2646 468 2664 486
rect 2646 486 2664 504
rect 2646 504 2664 522
rect 2646 522 2664 540
rect 2646 1062 2664 1080
rect 2646 1080 2664 1098
rect 2646 1098 2664 1116
rect 2646 1116 2664 1134
rect 2646 1134 2664 1152
rect 2646 1152 2664 1170
rect 2646 1170 2664 1188
rect 2646 1188 2664 1206
rect 2646 1206 2664 1224
rect 2646 1224 2664 1242
rect 2646 1242 2664 1260
rect 2646 1260 2664 1278
rect 2646 1278 2664 1296
rect 2646 1296 2664 1314
rect 2646 1314 2664 1332
rect 2646 1332 2664 1350
rect 2646 1350 2664 1368
rect 2646 1368 2664 1386
rect 2646 1386 2664 1404
rect 2646 1404 2664 1422
rect 2646 1422 2664 1440
rect 2646 1440 2664 1458
rect 2646 1458 2664 1476
rect 2646 1476 2664 1494
rect 2646 1494 2664 1512
rect 2646 1512 2664 1530
rect 2646 1530 2664 1548
rect 2646 1548 2664 1566
rect 2646 1566 2664 1584
rect 2646 1584 2664 1602
rect 2646 1602 2664 1620
rect 2646 1620 2664 1638
rect 2646 1638 2664 1656
rect 2646 1656 2664 1674
rect 2646 1674 2664 1692
rect 2646 1692 2664 1710
rect 2646 1710 2664 1728
rect 2646 1728 2664 1746
rect 2646 1746 2664 1764
rect 2646 1764 2664 1782
rect 2646 1782 2664 1800
rect 2646 1800 2664 1818
rect 2646 1818 2664 1836
rect 2646 1836 2664 1854
rect 2646 1854 2664 1872
rect 2646 1872 2664 1890
rect 2646 1890 2664 1908
rect 2646 1908 2664 1926
rect 2646 1926 2664 1944
rect 2646 1944 2664 1962
rect 2646 1962 2664 1980
rect 2646 1980 2664 1998
rect 2646 1998 2664 2016
rect 2646 2016 2664 2034
rect 2646 2034 2664 2052
rect 2646 2052 2664 2070
rect 2646 6480 2664 6498
rect 2646 6498 2664 6516
rect 2646 6516 2664 6534
rect 2646 6534 2664 6552
rect 2646 6552 2664 6570
rect 2646 6570 2664 6588
rect 2646 6588 2664 6606
rect 2646 6606 2664 6624
rect 2646 6624 2664 6642
rect 2646 6642 2664 6660
rect 2646 6660 2664 6678
rect 2646 6678 2664 6696
rect 2646 6696 2664 6714
rect 2646 6714 2664 6732
rect 2646 6732 2664 6750
rect 2646 6750 2664 6768
rect 2646 6768 2664 6786
rect 2646 6786 2664 6804
rect 2646 6804 2664 6822
rect 2646 6822 2664 6840
rect 2646 6840 2664 6858
rect 2646 6858 2664 6876
rect 2646 6876 2664 6894
rect 2646 6894 2664 6912
rect 2646 6912 2664 6930
rect 2646 6930 2664 6948
rect 2646 6948 2664 6966
rect 2646 6966 2664 6984
rect 2646 6984 2664 7002
rect 2646 7002 2664 7020
rect 2646 7020 2664 7038
rect 2646 7038 2664 7056
rect 2646 7056 2664 7074
rect 2646 7074 2664 7092
rect 2646 7092 2664 7110
rect 2646 7110 2664 7128
rect 2664 324 2682 342
rect 2664 342 2682 360
rect 2664 360 2682 378
rect 2664 378 2682 396
rect 2664 396 2682 414
rect 2664 414 2682 432
rect 2664 432 2682 450
rect 2664 450 2682 468
rect 2664 468 2682 486
rect 2664 486 2682 504
rect 2664 504 2682 522
rect 2664 522 2682 540
rect 2664 540 2682 558
rect 2664 1098 2682 1116
rect 2664 1116 2682 1134
rect 2664 1134 2682 1152
rect 2664 1152 2682 1170
rect 2664 1170 2682 1188
rect 2664 1188 2682 1206
rect 2664 1206 2682 1224
rect 2664 1224 2682 1242
rect 2664 1242 2682 1260
rect 2664 1260 2682 1278
rect 2664 1278 2682 1296
rect 2664 1296 2682 1314
rect 2664 1314 2682 1332
rect 2664 1332 2682 1350
rect 2664 1350 2682 1368
rect 2664 1368 2682 1386
rect 2664 1386 2682 1404
rect 2664 1404 2682 1422
rect 2664 1422 2682 1440
rect 2664 1440 2682 1458
rect 2664 1458 2682 1476
rect 2664 1476 2682 1494
rect 2664 1494 2682 1512
rect 2664 1512 2682 1530
rect 2664 1530 2682 1548
rect 2664 1548 2682 1566
rect 2664 1566 2682 1584
rect 2664 1584 2682 1602
rect 2664 1602 2682 1620
rect 2664 1620 2682 1638
rect 2664 1638 2682 1656
rect 2664 1656 2682 1674
rect 2664 1674 2682 1692
rect 2664 1692 2682 1710
rect 2664 1710 2682 1728
rect 2664 1728 2682 1746
rect 2664 1746 2682 1764
rect 2664 1764 2682 1782
rect 2664 1782 2682 1800
rect 2664 1800 2682 1818
rect 2664 1818 2682 1836
rect 2664 1836 2682 1854
rect 2664 1854 2682 1872
rect 2664 1872 2682 1890
rect 2664 1890 2682 1908
rect 2664 1908 2682 1926
rect 2664 1926 2682 1944
rect 2664 1944 2682 1962
rect 2664 1962 2682 1980
rect 2664 1980 2682 1998
rect 2664 1998 2682 2016
rect 2664 2016 2682 2034
rect 2664 2034 2682 2052
rect 2664 2052 2682 2070
rect 2664 2070 2682 2088
rect 2664 2088 2682 2106
rect 2664 2106 2682 2124
rect 2664 2124 2682 2142
rect 2664 6480 2682 6498
rect 2664 6498 2682 6516
rect 2664 6516 2682 6534
rect 2664 6534 2682 6552
rect 2664 6552 2682 6570
rect 2664 6570 2682 6588
rect 2664 6588 2682 6606
rect 2664 6606 2682 6624
rect 2664 6624 2682 6642
rect 2664 6642 2682 6660
rect 2664 6660 2682 6678
rect 2664 6678 2682 6696
rect 2664 6696 2682 6714
rect 2664 6714 2682 6732
rect 2664 6732 2682 6750
rect 2664 6750 2682 6768
rect 2664 6768 2682 6786
rect 2664 6786 2682 6804
rect 2664 6804 2682 6822
rect 2664 6822 2682 6840
rect 2664 6840 2682 6858
rect 2664 6858 2682 6876
rect 2664 6876 2682 6894
rect 2664 6894 2682 6912
rect 2664 6912 2682 6930
rect 2664 6930 2682 6948
rect 2664 6948 2682 6966
rect 2664 6966 2682 6984
rect 2664 6984 2682 7002
rect 2664 7002 2682 7020
rect 2664 7020 2682 7038
rect 2664 7038 2682 7056
rect 2664 7056 2682 7074
rect 2664 7074 2682 7092
rect 2664 7092 2682 7110
rect 2664 7110 2682 7128
rect 2664 7128 2682 7146
rect 2682 126 2700 144
rect 2682 342 2700 360
rect 2682 360 2700 378
rect 2682 378 2700 396
rect 2682 396 2700 414
rect 2682 414 2700 432
rect 2682 432 2700 450
rect 2682 450 2700 468
rect 2682 468 2700 486
rect 2682 486 2700 504
rect 2682 504 2700 522
rect 2682 522 2700 540
rect 2682 540 2700 558
rect 2682 558 2700 576
rect 2682 1134 2700 1152
rect 2682 1152 2700 1170
rect 2682 1170 2700 1188
rect 2682 1188 2700 1206
rect 2682 1206 2700 1224
rect 2682 1224 2700 1242
rect 2682 1242 2700 1260
rect 2682 1260 2700 1278
rect 2682 1278 2700 1296
rect 2682 1296 2700 1314
rect 2682 1314 2700 1332
rect 2682 1332 2700 1350
rect 2682 1350 2700 1368
rect 2682 1368 2700 1386
rect 2682 1386 2700 1404
rect 2682 1404 2700 1422
rect 2682 1422 2700 1440
rect 2682 1440 2700 1458
rect 2682 1458 2700 1476
rect 2682 1476 2700 1494
rect 2682 1494 2700 1512
rect 2682 1512 2700 1530
rect 2682 1530 2700 1548
rect 2682 1548 2700 1566
rect 2682 1566 2700 1584
rect 2682 1584 2700 1602
rect 2682 1602 2700 1620
rect 2682 1620 2700 1638
rect 2682 1638 2700 1656
rect 2682 1656 2700 1674
rect 2682 1674 2700 1692
rect 2682 1692 2700 1710
rect 2682 1710 2700 1728
rect 2682 1728 2700 1746
rect 2682 1746 2700 1764
rect 2682 1764 2700 1782
rect 2682 1782 2700 1800
rect 2682 1800 2700 1818
rect 2682 1818 2700 1836
rect 2682 1836 2700 1854
rect 2682 1854 2700 1872
rect 2682 1872 2700 1890
rect 2682 1890 2700 1908
rect 2682 1908 2700 1926
rect 2682 1926 2700 1944
rect 2682 1944 2700 1962
rect 2682 1962 2700 1980
rect 2682 1980 2700 1998
rect 2682 1998 2700 2016
rect 2682 2016 2700 2034
rect 2682 2034 2700 2052
rect 2682 2052 2700 2070
rect 2682 2070 2700 2088
rect 2682 2088 2700 2106
rect 2682 2106 2700 2124
rect 2682 2124 2700 2142
rect 2682 2142 2700 2160
rect 2682 2160 2700 2178
rect 2682 2178 2700 2196
rect 2682 2196 2700 2214
rect 2682 6498 2700 6516
rect 2682 6516 2700 6534
rect 2682 6534 2700 6552
rect 2682 6552 2700 6570
rect 2682 6570 2700 6588
rect 2682 6588 2700 6606
rect 2682 6606 2700 6624
rect 2682 6624 2700 6642
rect 2682 6642 2700 6660
rect 2682 6660 2700 6678
rect 2682 6678 2700 6696
rect 2682 6696 2700 6714
rect 2682 6714 2700 6732
rect 2682 6732 2700 6750
rect 2682 6750 2700 6768
rect 2682 6768 2700 6786
rect 2682 6786 2700 6804
rect 2682 6804 2700 6822
rect 2682 6822 2700 6840
rect 2682 6840 2700 6858
rect 2682 6858 2700 6876
rect 2682 6876 2700 6894
rect 2682 6894 2700 6912
rect 2682 6912 2700 6930
rect 2682 6930 2700 6948
rect 2682 6948 2700 6966
rect 2682 6966 2700 6984
rect 2682 6984 2700 7002
rect 2682 7002 2700 7020
rect 2682 7020 2700 7038
rect 2682 7038 2700 7056
rect 2682 7056 2700 7074
rect 2682 7074 2700 7092
rect 2682 7092 2700 7110
rect 2682 7110 2700 7128
rect 2682 7128 2700 7146
rect 2700 126 2718 144
rect 2700 144 2718 162
rect 2700 342 2718 360
rect 2700 360 2718 378
rect 2700 378 2718 396
rect 2700 396 2718 414
rect 2700 414 2718 432
rect 2700 432 2718 450
rect 2700 450 2718 468
rect 2700 468 2718 486
rect 2700 486 2718 504
rect 2700 504 2718 522
rect 2700 522 2718 540
rect 2700 540 2718 558
rect 2700 558 2718 576
rect 2700 576 2718 594
rect 2700 1170 2718 1188
rect 2700 1188 2718 1206
rect 2700 1206 2718 1224
rect 2700 1224 2718 1242
rect 2700 1242 2718 1260
rect 2700 1260 2718 1278
rect 2700 1278 2718 1296
rect 2700 1296 2718 1314
rect 2700 1314 2718 1332
rect 2700 1332 2718 1350
rect 2700 1350 2718 1368
rect 2700 1368 2718 1386
rect 2700 1386 2718 1404
rect 2700 1404 2718 1422
rect 2700 1422 2718 1440
rect 2700 1440 2718 1458
rect 2700 1458 2718 1476
rect 2700 1476 2718 1494
rect 2700 1494 2718 1512
rect 2700 1512 2718 1530
rect 2700 1530 2718 1548
rect 2700 1548 2718 1566
rect 2700 1566 2718 1584
rect 2700 1584 2718 1602
rect 2700 1602 2718 1620
rect 2700 1620 2718 1638
rect 2700 1638 2718 1656
rect 2700 1656 2718 1674
rect 2700 1674 2718 1692
rect 2700 1692 2718 1710
rect 2700 1710 2718 1728
rect 2700 1728 2718 1746
rect 2700 1746 2718 1764
rect 2700 1764 2718 1782
rect 2700 1782 2718 1800
rect 2700 1800 2718 1818
rect 2700 1818 2718 1836
rect 2700 1836 2718 1854
rect 2700 1854 2718 1872
rect 2700 1872 2718 1890
rect 2700 1890 2718 1908
rect 2700 1908 2718 1926
rect 2700 1926 2718 1944
rect 2700 1944 2718 1962
rect 2700 1962 2718 1980
rect 2700 1980 2718 1998
rect 2700 1998 2718 2016
rect 2700 2016 2718 2034
rect 2700 2034 2718 2052
rect 2700 2052 2718 2070
rect 2700 2070 2718 2088
rect 2700 2088 2718 2106
rect 2700 2106 2718 2124
rect 2700 2124 2718 2142
rect 2700 2142 2718 2160
rect 2700 2160 2718 2178
rect 2700 2178 2718 2196
rect 2700 2196 2718 2214
rect 2700 2214 2718 2232
rect 2700 2232 2718 2250
rect 2700 2250 2718 2268
rect 2700 2268 2718 2286
rect 2700 6498 2718 6516
rect 2700 6516 2718 6534
rect 2700 6534 2718 6552
rect 2700 6552 2718 6570
rect 2700 6570 2718 6588
rect 2700 6588 2718 6606
rect 2700 6606 2718 6624
rect 2700 6624 2718 6642
rect 2700 6642 2718 6660
rect 2700 6660 2718 6678
rect 2700 6678 2718 6696
rect 2700 6696 2718 6714
rect 2700 6714 2718 6732
rect 2700 6732 2718 6750
rect 2700 6750 2718 6768
rect 2700 6768 2718 6786
rect 2700 6786 2718 6804
rect 2700 6804 2718 6822
rect 2700 6822 2718 6840
rect 2700 6840 2718 6858
rect 2700 6858 2718 6876
rect 2700 6876 2718 6894
rect 2700 6894 2718 6912
rect 2700 6912 2718 6930
rect 2700 6930 2718 6948
rect 2700 6948 2718 6966
rect 2700 6966 2718 6984
rect 2700 6984 2718 7002
rect 2700 7002 2718 7020
rect 2700 7020 2718 7038
rect 2700 7038 2718 7056
rect 2700 7056 2718 7074
rect 2700 7074 2718 7092
rect 2700 7092 2718 7110
rect 2700 7110 2718 7128
rect 2700 7128 2718 7146
rect 2718 126 2736 144
rect 2718 144 2736 162
rect 2718 162 2736 180
rect 2718 360 2736 378
rect 2718 378 2736 396
rect 2718 396 2736 414
rect 2718 414 2736 432
rect 2718 432 2736 450
rect 2718 450 2736 468
rect 2718 468 2736 486
rect 2718 486 2736 504
rect 2718 504 2736 522
rect 2718 522 2736 540
rect 2718 540 2736 558
rect 2718 558 2736 576
rect 2718 576 2736 594
rect 2718 594 2736 612
rect 2718 1206 2736 1224
rect 2718 1224 2736 1242
rect 2718 1242 2736 1260
rect 2718 1260 2736 1278
rect 2718 1278 2736 1296
rect 2718 1296 2736 1314
rect 2718 1314 2736 1332
rect 2718 1332 2736 1350
rect 2718 1350 2736 1368
rect 2718 1368 2736 1386
rect 2718 1386 2736 1404
rect 2718 1404 2736 1422
rect 2718 1422 2736 1440
rect 2718 1440 2736 1458
rect 2718 1458 2736 1476
rect 2718 1476 2736 1494
rect 2718 1494 2736 1512
rect 2718 1512 2736 1530
rect 2718 1530 2736 1548
rect 2718 1548 2736 1566
rect 2718 1566 2736 1584
rect 2718 1584 2736 1602
rect 2718 1602 2736 1620
rect 2718 1620 2736 1638
rect 2718 1638 2736 1656
rect 2718 1656 2736 1674
rect 2718 1674 2736 1692
rect 2718 1692 2736 1710
rect 2718 1710 2736 1728
rect 2718 1728 2736 1746
rect 2718 1746 2736 1764
rect 2718 1764 2736 1782
rect 2718 1782 2736 1800
rect 2718 1800 2736 1818
rect 2718 1818 2736 1836
rect 2718 1836 2736 1854
rect 2718 1854 2736 1872
rect 2718 1872 2736 1890
rect 2718 1890 2736 1908
rect 2718 1908 2736 1926
rect 2718 1926 2736 1944
rect 2718 1944 2736 1962
rect 2718 1962 2736 1980
rect 2718 1980 2736 1998
rect 2718 1998 2736 2016
rect 2718 2016 2736 2034
rect 2718 2034 2736 2052
rect 2718 2052 2736 2070
rect 2718 2070 2736 2088
rect 2718 2088 2736 2106
rect 2718 2106 2736 2124
rect 2718 2124 2736 2142
rect 2718 2142 2736 2160
rect 2718 2160 2736 2178
rect 2718 2178 2736 2196
rect 2718 2196 2736 2214
rect 2718 2214 2736 2232
rect 2718 2232 2736 2250
rect 2718 2250 2736 2268
rect 2718 2268 2736 2286
rect 2718 2286 2736 2304
rect 2718 2304 2736 2322
rect 2718 2322 2736 2340
rect 2718 6498 2736 6516
rect 2718 6516 2736 6534
rect 2718 6534 2736 6552
rect 2718 6552 2736 6570
rect 2718 6570 2736 6588
rect 2718 6588 2736 6606
rect 2718 6606 2736 6624
rect 2718 6624 2736 6642
rect 2718 6642 2736 6660
rect 2718 6660 2736 6678
rect 2718 6678 2736 6696
rect 2718 6696 2736 6714
rect 2718 6714 2736 6732
rect 2718 6732 2736 6750
rect 2718 6750 2736 6768
rect 2718 6768 2736 6786
rect 2718 6786 2736 6804
rect 2718 6804 2736 6822
rect 2718 6822 2736 6840
rect 2718 6840 2736 6858
rect 2718 6858 2736 6876
rect 2718 6876 2736 6894
rect 2718 6894 2736 6912
rect 2718 6912 2736 6930
rect 2718 6930 2736 6948
rect 2718 6948 2736 6966
rect 2718 6966 2736 6984
rect 2718 6984 2736 7002
rect 2718 7002 2736 7020
rect 2718 7020 2736 7038
rect 2718 7038 2736 7056
rect 2718 7056 2736 7074
rect 2718 7074 2736 7092
rect 2718 7092 2736 7110
rect 2718 7110 2736 7128
rect 2718 7128 2736 7146
rect 2718 7146 2736 7164
rect 2736 126 2754 144
rect 2736 144 2754 162
rect 2736 162 2754 180
rect 2736 378 2754 396
rect 2736 396 2754 414
rect 2736 414 2754 432
rect 2736 432 2754 450
rect 2736 450 2754 468
rect 2736 468 2754 486
rect 2736 486 2754 504
rect 2736 504 2754 522
rect 2736 522 2754 540
rect 2736 540 2754 558
rect 2736 558 2754 576
rect 2736 576 2754 594
rect 2736 594 2754 612
rect 2736 612 2754 630
rect 2736 846 2754 864
rect 2736 1242 2754 1260
rect 2736 1260 2754 1278
rect 2736 1278 2754 1296
rect 2736 1296 2754 1314
rect 2736 1314 2754 1332
rect 2736 1332 2754 1350
rect 2736 1350 2754 1368
rect 2736 1368 2754 1386
rect 2736 1386 2754 1404
rect 2736 1404 2754 1422
rect 2736 1422 2754 1440
rect 2736 1440 2754 1458
rect 2736 1458 2754 1476
rect 2736 1476 2754 1494
rect 2736 1494 2754 1512
rect 2736 1512 2754 1530
rect 2736 1530 2754 1548
rect 2736 1548 2754 1566
rect 2736 1566 2754 1584
rect 2736 1584 2754 1602
rect 2736 1602 2754 1620
rect 2736 1620 2754 1638
rect 2736 1638 2754 1656
rect 2736 1656 2754 1674
rect 2736 1674 2754 1692
rect 2736 1692 2754 1710
rect 2736 1710 2754 1728
rect 2736 1728 2754 1746
rect 2736 1746 2754 1764
rect 2736 1764 2754 1782
rect 2736 1782 2754 1800
rect 2736 1800 2754 1818
rect 2736 1818 2754 1836
rect 2736 1836 2754 1854
rect 2736 1854 2754 1872
rect 2736 1872 2754 1890
rect 2736 1890 2754 1908
rect 2736 1908 2754 1926
rect 2736 1926 2754 1944
rect 2736 1944 2754 1962
rect 2736 1962 2754 1980
rect 2736 1980 2754 1998
rect 2736 1998 2754 2016
rect 2736 2016 2754 2034
rect 2736 2034 2754 2052
rect 2736 2052 2754 2070
rect 2736 2070 2754 2088
rect 2736 2088 2754 2106
rect 2736 2106 2754 2124
rect 2736 2124 2754 2142
rect 2736 2142 2754 2160
rect 2736 2160 2754 2178
rect 2736 2178 2754 2196
rect 2736 2196 2754 2214
rect 2736 2214 2754 2232
rect 2736 2232 2754 2250
rect 2736 2250 2754 2268
rect 2736 2268 2754 2286
rect 2736 2286 2754 2304
rect 2736 2304 2754 2322
rect 2736 2322 2754 2340
rect 2736 2340 2754 2358
rect 2736 2358 2754 2376
rect 2736 2376 2754 2394
rect 2736 2394 2754 2412
rect 2736 6516 2754 6534
rect 2736 6534 2754 6552
rect 2736 6552 2754 6570
rect 2736 6570 2754 6588
rect 2736 6588 2754 6606
rect 2736 6606 2754 6624
rect 2736 6624 2754 6642
rect 2736 6642 2754 6660
rect 2736 6660 2754 6678
rect 2736 6678 2754 6696
rect 2736 6696 2754 6714
rect 2736 6714 2754 6732
rect 2736 6732 2754 6750
rect 2736 6750 2754 6768
rect 2736 6768 2754 6786
rect 2736 6786 2754 6804
rect 2736 6804 2754 6822
rect 2736 6822 2754 6840
rect 2736 6840 2754 6858
rect 2736 6858 2754 6876
rect 2736 6876 2754 6894
rect 2736 6894 2754 6912
rect 2736 6912 2754 6930
rect 2736 6930 2754 6948
rect 2736 6948 2754 6966
rect 2736 6966 2754 6984
rect 2736 6984 2754 7002
rect 2736 7002 2754 7020
rect 2736 7020 2754 7038
rect 2736 7038 2754 7056
rect 2736 7056 2754 7074
rect 2736 7074 2754 7092
rect 2736 7092 2754 7110
rect 2736 7110 2754 7128
rect 2736 7128 2754 7146
rect 2736 7146 2754 7164
rect 2754 108 2772 126
rect 2754 126 2772 144
rect 2754 144 2772 162
rect 2754 162 2772 180
rect 2754 180 2772 198
rect 2754 378 2772 396
rect 2754 396 2772 414
rect 2754 414 2772 432
rect 2754 432 2772 450
rect 2754 450 2772 468
rect 2754 468 2772 486
rect 2754 486 2772 504
rect 2754 504 2772 522
rect 2754 522 2772 540
rect 2754 540 2772 558
rect 2754 558 2772 576
rect 2754 576 2772 594
rect 2754 594 2772 612
rect 2754 612 2772 630
rect 2754 630 2772 648
rect 2754 846 2772 864
rect 2754 864 2772 882
rect 2754 882 2772 900
rect 2754 1278 2772 1296
rect 2754 1296 2772 1314
rect 2754 1314 2772 1332
rect 2754 1332 2772 1350
rect 2754 1350 2772 1368
rect 2754 1368 2772 1386
rect 2754 1386 2772 1404
rect 2754 1404 2772 1422
rect 2754 1422 2772 1440
rect 2754 1440 2772 1458
rect 2754 1458 2772 1476
rect 2754 1476 2772 1494
rect 2754 1494 2772 1512
rect 2754 1512 2772 1530
rect 2754 1530 2772 1548
rect 2754 1548 2772 1566
rect 2754 1566 2772 1584
rect 2754 1584 2772 1602
rect 2754 1602 2772 1620
rect 2754 1620 2772 1638
rect 2754 1638 2772 1656
rect 2754 1656 2772 1674
rect 2754 1674 2772 1692
rect 2754 1692 2772 1710
rect 2754 1710 2772 1728
rect 2754 1728 2772 1746
rect 2754 1746 2772 1764
rect 2754 1764 2772 1782
rect 2754 1782 2772 1800
rect 2754 1800 2772 1818
rect 2754 1818 2772 1836
rect 2754 1836 2772 1854
rect 2754 1854 2772 1872
rect 2754 1872 2772 1890
rect 2754 1890 2772 1908
rect 2754 1908 2772 1926
rect 2754 1926 2772 1944
rect 2754 1944 2772 1962
rect 2754 1962 2772 1980
rect 2754 1980 2772 1998
rect 2754 1998 2772 2016
rect 2754 2016 2772 2034
rect 2754 2034 2772 2052
rect 2754 2052 2772 2070
rect 2754 2070 2772 2088
rect 2754 2088 2772 2106
rect 2754 2106 2772 2124
rect 2754 2124 2772 2142
rect 2754 2142 2772 2160
rect 2754 2160 2772 2178
rect 2754 2178 2772 2196
rect 2754 2196 2772 2214
rect 2754 2214 2772 2232
rect 2754 2232 2772 2250
rect 2754 2250 2772 2268
rect 2754 2268 2772 2286
rect 2754 2286 2772 2304
rect 2754 2304 2772 2322
rect 2754 2322 2772 2340
rect 2754 2340 2772 2358
rect 2754 2358 2772 2376
rect 2754 2376 2772 2394
rect 2754 2394 2772 2412
rect 2754 2412 2772 2430
rect 2754 2430 2772 2448
rect 2754 2448 2772 2466
rect 2754 2466 2772 2484
rect 2754 6516 2772 6534
rect 2754 6534 2772 6552
rect 2754 6552 2772 6570
rect 2754 6570 2772 6588
rect 2754 6588 2772 6606
rect 2754 6606 2772 6624
rect 2754 6624 2772 6642
rect 2754 6642 2772 6660
rect 2754 6660 2772 6678
rect 2754 6678 2772 6696
rect 2754 6696 2772 6714
rect 2754 6714 2772 6732
rect 2754 6732 2772 6750
rect 2754 6750 2772 6768
rect 2754 6768 2772 6786
rect 2754 6786 2772 6804
rect 2754 6804 2772 6822
rect 2754 6822 2772 6840
rect 2754 6840 2772 6858
rect 2754 6858 2772 6876
rect 2754 6876 2772 6894
rect 2754 6894 2772 6912
rect 2754 6912 2772 6930
rect 2754 6930 2772 6948
rect 2754 6948 2772 6966
rect 2754 6966 2772 6984
rect 2754 6984 2772 7002
rect 2754 7002 2772 7020
rect 2754 7020 2772 7038
rect 2754 7038 2772 7056
rect 2754 7056 2772 7074
rect 2754 7074 2772 7092
rect 2754 7092 2772 7110
rect 2754 7110 2772 7128
rect 2754 7128 2772 7146
rect 2754 7146 2772 7164
rect 2772 108 2790 126
rect 2772 126 2790 144
rect 2772 144 2790 162
rect 2772 162 2790 180
rect 2772 180 2790 198
rect 2772 198 2790 216
rect 2772 396 2790 414
rect 2772 414 2790 432
rect 2772 432 2790 450
rect 2772 450 2790 468
rect 2772 468 2790 486
rect 2772 486 2790 504
rect 2772 504 2790 522
rect 2772 522 2790 540
rect 2772 540 2790 558
rect 2772 558 2790 576
rect 2772 576 2790 594
rect 2772 594 2790 612
rect 2772 612 2790 630
rect 2772 630 2790 648
rect 2772 648 2790 666
rect 2772 864 2790 882
rect 2772 882 2790 900
rect 2772 900 2790 918
rect 2772 918 2790 936
rect 2772 936 2790 954
rect 2772 1314 2790 1332
rect 2772 1332 2790 1350
rect 2772 1350 2790 1368
rect 2772 1368 2790 1386
rect 2772 1386 2790 1404
rect 2772 1404 2790 1422
rect 2772 1422 2790 1440
rect 2772 1440 2790 1458
rect 2772 1458 2790 1476
rect 2772 1476 2790 1494
rect 2772 1494 2790 1512
rect 2772 1512 2790 1530
rect 2772 1530 2790 1548
rect 2772 1548 2790 1566
rect 2772 1566 2790 1584
rect 2772 1584 2790 1602
rect 2772 1602 2790 1620
rect 2772 1620 2790 1638
rect 2772 1638 2790 1656
rect 2772 1656 2790 1674
rect 2772 1674 2790 1692
rect 2772 1692 2790 1710
rect 2772 1710 2790 1728
rect 2772 1728 2790 1746
rect 2772 1746 2790 1764
rect 2772 1764 2790 1782
rect 2772 1782 2790 1800
rect 2772 1800 2790 1818
rect 2772 1818 2790 1836
rect 2772 1836 2790 1854
rect 2772 1854 2790 1872
rect 2772 1872 2790 1890
rect 2772 1890 2790 1908
rect 2772 1908 2790 1926
rect 2772 1926 2790 1944
rect 2772 1944 2790 1962
rect 2772 1962 2790 1980
rect 2772 1980 2790 1998
rect 2772 1998 2790 2016
rect 2772 2016 2790 2034
rect 2772 2034 2790 2052
rect 2772 2052 2790 2070
rect 2772 2070 2790 2088
rect 2772 2088 2790 2106
rect 2772 2106 2790 2124
rect 2772 2124 2790 2142
rect 2772 2142 2790 2160
rect 2772 2160 2790 2178
rect 2772 2178 2790 2196
rect 2772 2196 2790 2214
rect 2772 2214 2790 2232
rect 2772 2232 2790 2250
rect 2772 2250 2790 2268
rect 2772 2268 2790 2286
rect 2772 2286 2790 2304
rect 2772 2304 2790 2322
rect 2772 2322 2790 2340
rect 2772 2340 2790 2358
rect 2772 2358 2790 2376
rect 2772 2376 2790 2394
rect 2772 2394 2790 2412
rect 2772 2412 2790 2430
rect 2772 2430 2790 2448
rect 2772 2448 2790 2466
rect 2772 2466 2790 2484
rect 2772 2484 2790 2502
rect 2772 2502 2790 2520
rect 2772 2520 2790 2538
rect 2772 2538 2790 2556
rect 2772 6516 2790 6534
rect 2772 6534 2790 6552
rect 2772 6552 2790 6570
rect 2772 6570 2790 6588
rect 2772 6588 2790 6606
rect 2772 6606 2790 6624
rect 2772 6624 2790 6642
rect 2772 6642 2790 6660
rect 2772 6660 2790 6678
rect 2772 6678 2790 6696
rect 2772 6696 2790 6714
rect 2772 6714 2790 6732
rect 2772 6732 2790 6750
rect 2772 6750 2790 6768
rect 2772 6768 2790 6786
rect 2772 6786 2790 6804
rect 2772 6804 2790 6822
rect 2772 6822 2790 6840
rect 2772 6840 2790 6858
rect 2772 6858 2790 6876
rect 2772 6876 2790 6894
rect 2772 6894 2790 6912
rect 2772 6912 2790 6930
rect 2772 6930 2790 6948
rect 2772 6948 2790 6966
rect 2772 6966 2790 6984
rect 2772 6984 2790 7002
rect 2772 7002 2790 7020
rect 2772 7020 2790 7038
rect 2772 7038 2790 7056
rect 2772 7056 2790 7074
rect 2772 7074 2790 7092
rect 2772 7092 2790 7110
rect 2772 7110 2790 7128
rect 2772 7128 2790 7146
rect 2772 7146 2790 7164
rect 2790 108 2808 126
rect 2790 126 2808 144
rect 2790 144 2808 162
rect 2790 162 2808 180
rect 2790 180 2808 198
rect 2790 198 2808 216
rect 2790 216 2808 234
rect 2790 414 2808 432
rect 2790 432 2808 450
rect 2790 450 2808 468
rect 2790 468 2808 486
rect 2790 486 2808 504
rect 2790 504 2808 522
rect 2790 522 2808 540
rect 2790 540 2808 558
rect 2790 558 2808 576
rect 2790 576 2808 594
rect 2790 594 2808 612
rect 2790 612 2808 630
rect 2790 630 2808 648
rect 2790 648 2808 666
rect 2790 666 2808 684
rect 2790 882 2808 900
rect 2790 900 2808 918
rect 2790 918 2808 936
rect 2790 936 2808 954
rect 2790 954 2808 972
rect 2790 972 2808 990
rect 2790 990 2808 1008
rect 2790 1350 2808 1368
rect 2790 1368 2808 1386
rect 2790 1386 2808 1404
rect 2790 1404 2808 1422
rect 2790 1422 2808 1440
rect 2790 1440 2808 1458
rect 2790 1458 2808 1476
rect 2790 1476 2808 1494
rect 2790 1494 2808 1512
rect 2790 1512 2808 1530
rect 2790 1530 2808 1548
rect 2790 1548 2808 1566
rect 2790 1566 2808 1584
rect 2790 1584 2808 1602
rect 2790 1602 2808 1620
rect 2790 1620 2808 1638
rect 2790 1638 2808 1656
rect 2790 1656 2808 1674
rect 2790 1674 2808 1692
rect 2790 1692 2808 1710
rect 2790 1710 2808 1728
rect 2790 1728 2808 1746
rect 2790 1746 2808 1764
rect 2790 1764 2808 1782
rect 2790 1782 2808 1800
rect 2790 1800 2808 1818
rect 2790 1818 2808 1836
rect 2790 1836 2808 1854
rect 2790 1854 2808 1872
rect 2790 1872 2808 1890
rect 2790 1890 2808 1908
rect 2790 1908 2808 1926
rect 2790 1926 2808 1944
rect 2790 1944 2808 1962
rect 2790 1962 2808 1980
rect 2790 1980 2808 1998
rect 2790 1998 2808 2016
rect 2790 2016 2808 2034
rect 2790 2034 2808 2052
rect 2790 2052 2808 2070
rect 2790 2070 2808 2088
rect 2790 2088 2808 2106
rect 2790 2106 2808 2124
rect 2790 2124 2808 2142
rect 2790 2142 2808 2160
rect 2790 2160 2808 2178
rect 2790 2178 2808 2196
rect 2790 2196 2808 2214
rect 2790 2214 2808 2232
rect 2790 2232 2808 2250
rect 2790 2250 2808 2268
rect 2790 2268 2808 2286
rect 2790 2286 2808 2304
rect 2790 2304 2808 2322
rect 2790 2322 2808 2340
rect 2790 2340 2808 2358
rect 2790 2358 2808 2376
rect 2790 2376 2808 2394
rect 2790 2394 2808 2412
rect 2790 2412 2808 2430
rect 2790 2430 2808 2448
rect 2790 2448 2808 2466
rect 2790 2466 2808 2484
rect 2790 2484 2808 2502
rect 2790 2502 2808 2520
rect 2790 2520 2808 2538
rect 2790 2538 2808 2556
rect 2790 2556 2808 2574
rect 2790 2574 2808 2592
rect 2790 2592 2808 2610
rect 2790 6534 2808 6552
rect 2790 6552 2808 6570
rect 2790 6570 2808 6588
rect 2790 6588 2808 6606
rect 2790 6606 2808 6624
rect 2790 6624 2808 6642
rect 2790 6642 2808 6660
rect 2790 6660 2808 6678
rect 2790 6678 2808 6696
rect 2790 6696 2808 6714
rect 2790 6714 2808 6732
rect 2790 6732 2808 6750
rect 2790 6750 2808 6768
rect 2790 6768 2808 6786
rect 2790 6786 2808 6804
rect 2790 6804 2808 6822
rect 2790 6822 2808 6840
rect 2790 6840 2808 6858
rect 2790 6858 2808 6876
rect 2790 6876 2808 6894
rect 2790 6894 2808 6912
rect 2790 6912 2808 6930
rect 2790 6930 2808 6948
rect 2790 6948 2808 6966
rect 2790 6966 2808 6984
rect 2790 6984 2808 7002
rect 2790 7002 2808 7020
rect 2790 7020 2808 7038
rect 2790 7038 2808 7056
rect 2790 7056 2808 7074
rect 2790 7074 2808 7092
rect 2790 7092 2808 7110
rect 2790 7110 2808 7128
rect 2790 7128 2808 7146
rect 2790 7146 2808 7164
rect 2790 7164 2808 7182
rect 2808 108 2826 126
rect 2808 126 2826 144
rect 2808 144 2826 162
rect 2808 162 2826 180
rect 2808 180 2826 198
rect 2808 198 2826 216
rect 2808 216 2826 234
rect 2808 234 2826 252
rect 2808 432 2826 450
rect 2808 450 2826 468
rect 2808 468 2826 486
rect 2808 486 2826 504
rect 2808 504 2826 522
rect 2808 522 2826 540
rect 2808 540 2826 558
rect 2808 558 2826 576
rect 2808 576 2826 594
rect 2808 594 2826 612
rect 2808 612 2826 630
rect 2808 630 2826 648
rect 2808 648 2826 666
rect 2808 666 2826 684
rect 2808 684 2826 702
rect 2808 900 2826 918
rect 2808 918 2826 936
rect 2808 936 2826 954
rect 2808 954 2826 972
rect 2808 972 2826 990
rect 2808 990 2826 1008
rect 2808 1008 2826 1026
rect 2808 1026 2826 1044
rect 2808 1386 2826 1404
rect 2808 1404 2826 1422
rect 2808 1422 2826 1440
rect 2808 1440 2826 1458
rect 2808 1458 2826 1476
rect 2808 1476 2826 1494
rect 2808 1494 2826 1512
rect 2808 1512 2826 1530
rect 2808 1530 2826 1548
rect 2808 1548 2826 1566
rect 2808 1566 2826 1584
rect 2808 1584 2826 1602
rect 2808 1602 2826 1620
rect 2808 1620 2826 1638
rect 2808 1638 2826 1656
rect 2808 1656 2826 1674
rect 2808 1674 2826 1692
rect 2808 1692 2826 1710
rect 2808 1710 2826 1728
rect 2808 1728 2826 1746
rect 2808 1746 2826 1764
rect 2808 1764 2826 1782
rect 2808 1782 2826 1800
rect 2808 1800 2826 1818
rect 2808 1818 2826 1836
rect 2808 1836 2826 1854
rect 2808 1854 2826 1872
rect 2808 1872 2826 1890
rect 2808 1890 2826 1908
rect 2808 1908 2826 1926
rect 2808 1926 2826 1944
rect 2808 1944 2826 1962
rect 2808 1962 2826 1980
rect 2808 1980 2826 1998
rect 2808 1998 2826 2016
rect 2808 2016 2826 2034
rect 2808 2034 2826 2052
rect 2808 2052 2826 2070
rect 2808 2070 2826 2088
rect 2808 2088 2826 2106
rect 2808 2106 2826 2124
rect 2808 2124 2826 2142
rect 2808 2142 2826 2160
rect 2808 2160 2826 2178
rect 2808 2178 2826 2196
rect 2808 2196 2826 2214
rect 2808 2214 2826 2232
rect 2808 2232 2826 2250
rect 2808 2250 2826 2268
rect 2808 2268 2826 2286
rect 2808 2286 2826 2304
rect 2808 2304 2826 2322
rect 2808 2322 2826 2340
rect 2808 2340 2826 2358
rect 2808 2358 2826 2376
rect 2808 2376 2826 2394
rect 2808 2394 2826 2412
rect 2808 2412 2826 2430
rect 2808 2430 2826 2448
rect 2808 2448 2826 2466
rect 2808 2466 2826 2484
rect 2808 2484 2826 2502
rect 2808 2502 2826 2520
rect 2808 2520 2826 2538
rect 2808 2538 2826 2556
rect 2808 2556 2826 2574
rect 2808 2574 2826 2592
rect 2808 2592 2826 2610
rect 2808 2610 2826 2628
rect 2808 2628 2826 2646
rect 2808 2646 2826 2664
rect 2808 2664 2826 2682
rect 2808 6534 2826 6552
rect 2808 6552 2826 6570
rect 2808 6570 2826 6588
rect 2808 6588 2826 6606
rect 2808 6606 2826 6624
rect 2808 6624 2826 6642
rect 2808 6642 2826 6660
rect 2808 6660 2826 6678
rect 2808 6678 2826 6696
rect 2808 6696 2826 6714
rect 2808 6714 2826 6732
rect 2808 6732 2826 6750
rect 2808 6750 2826 6768
rect 2808 6768 2826 6786
rect 2808 6786 2826 6804
rect 2808 6804 2826 6822
rect 2808 6822 2826 6840
rect 2808 6840 2826 6858
rect 2808 6858 2826 6876
rect 2808 6876 2826 6894
rect 2808 6894 2826 6912
rect 2808 6912 2826 6930
rect 2808 6930 2826 6948
rect 2808 6948 2826 6966
rect 2808 6966 2826 6984
rect 2808 6984 2826 7002
rect 2808 7002 2826 7020
rect 2808 7020 2826 7038
rect 2808 7038 2826 7056
rect 2808 7056 2826 7074
rect 2808 7074 2826 7092
rect 2808 7092 2826 7110
rect 2808 7110 2826 7128
rect 2808 7128 2826 7146
rect 2808 7146 2826 7164
rect 2808 7164 2826 7182
rect 2826 108 2844 126
rect 2826 126 2844 144
rect 2826 144 2844 162
rect 2826 162 2844 180
rect 2826 180 2844 198
rect 2826 198 2844 216
rect 2826 216 2844 234
rect 2826 234 2844 252
rect 2826 432 2844 450
rect 2826 450 2844 468
rect 2826 468 2844 486
rect 2826 486 2844 504
rect 2826 504 2844 522
rect 2826 522 2844 540
rect 2826 540 2844 558
rect 2826 558 2844 576
rect 2826 576 2844 594
rect 2826 594 2844 612
rect 2826 612 2844 630
rect 2826 630 2844 648
rect 2826 648 2844 666
rect 2826 666 2844 684
rect 2826 684 2844 702
rect 2826 702 2844 720
rect 2826 900 2844 918
rect 2826 918 2844 936
rect 2826 936 2844 954
rect 2826 954 2844 972
rect 2826 972 2844 990
rect 2826 990 2844 1008
rect 2826 1008 2844 1026
rect 2826 1026 2844 1044
rect 2826 1044 2844 1062
rect 2826 1062 2844 1080
rect 2826 1080 2844 1098
rect 2826 1422 2844 1440
rect 2826 1440 2844 1458
rect 2826 1458 2844 1476
rect 2826 1476 2844 1494
rect 2826 1494 2844 1512
rect 2826 1512 2844 1530
rect 2826 1530 2844 1548
rect 2826 1548 2844 1566
rect 2826 1566 2844 1584
rect 2826 1584 2844 1602
rect 2826 1602 2844 1620
rect 2826 1620 2844 1638
rect 2826 1638 2844 1656
rect 2826 1656 2844 1674
rect 2826 1674 2844 1692
rect 2826 1692 2844 1710
rect 2826 1710 2844 1728
rect 2826 1728 2844 1746
rect 2826 1746 2844 1764
rect 2826 1764 2844 1782
rect 2826 1782 2844 1800
rect 2826 1800 2844 1818
rect 2826 1818 2844 1836
rect 2826 1836 2844 1854
rect 2826 1854 2844 1872
rect 2826 1872 2844 1890
rect 2826 1890 2844 1908
rect 2826 1908 2844 1926
rect 2826 1926 2844 1944
rect 2826 1944 2844 1962
rect 2826 1962 2844 1980
rect 2826 1980 2844 1998
rect 2826 1998 2844 2016
rect 2826 2016 2844 2034
rect 2826 2034 2844 2052
rect 2826 2052 2844 2070
rect 2826 2070 2844 2088
rect 2826 2088 2844 2106
rect 2826 2106 2844 2124
rect 2826 2124 2844 2142
rect 2826 2142 2844 2160
rect 2826 2160 2844 2178
rect 2826 2178 2844 2196
rect 2826 2196 2844 2214
rect 2826 2214 2844 2232
rect 2826 2232 2844 2250
rect 2826 2250 2844 2268
rect 2826 2268 2844 2286
rect 2826 2286 2844 2304
rect 2826 2304 2844 2322
rect 2826 2322 2844 2340
rect 2826 2340 2844 2358
rect 2826 2358 2844 2376
rect 2826 2376 2844 2394
rect 2826 2394 2844 2412
rect 2826 2412 2844 2430
rect 2826 2430 2844 2448
rect 2826 2448 2844 2466
rect 2826 2466 2844 2484
rect 2826 2484 2844 2502
rect 2826 2502 2844 2520
rect 2826 2520 2844 2538
rect 2826 2538 2844 2556
rect 2826 2556 2844 2574
rect 2826 2574 2844 2592
rect 2826 2592 2844 2610
rect 2826 2610 2844 2628
rect 2826 2628 2844 2646
rect 2826 2646 2844 2664
rect 2826 2664 2844 2682
rect 2826 2682 2844 2700
rect 2826 2700 2844 2718
rect 2826 2718 2844 2736
rect 2826 6534 2844 6552
rect 2826 6552 2844 6570
rect 2826 6570 2844 6588
rect 2826 6588 2844 6606
rect 2826 6606 2844 6624
rect 2826 6624 2844 6642
rect 2826 6642 2844 6660
rect 2826 6660 2844 6678
rect 2826 6678 2844 6696
rect 2826 6696 2844 6714
rect 2826 6714 2844 6732
rect 2826 6732 2844 6750
rect 2826 6750 2844 6768
rect 2826 6768 2844 6786
rect 2826 6786 2844 6804
rect 2826 6804 2844 6822
rect 2826 6822 2844 6840
rect 2826 6840 2844 6858
rect 2826 6858 2844 6876
rect 2826 6876 2844 6894
rect 2826 6894 2844 6912
rect 2826 6912 2844 6930
rect 2826 6930 2844 6948
rect 2826 6948 2844 6966
rect 2826 6966 2844 6984
rect 2826 6984 2844 7002
rect 2826 7002 2844 7020
rect 2826 7020 2844 7038
rect 2826 7038 2844 7056
rect 2826 7056 2844 7074
rect 2826 7074 2844 7092
rect 2826 7092 2844 7110
rect 2826 7110 2844 7128
rect 2826 7128 2844 7146
rect 2826 7146 2844 7164
rect 2826 7164 2844 7182
rect 2844 108 2862 126
rect 2844 126 2862 144
rect 2844 144 2862 162
rect 2844 162 2862 180
rect 2844 180 2862 198
rect 2844 198 2862 216
rect 2844 216 2862 234
rect 2844 234 2862 252
rect 2844 252 2862 270
rect 2844 450 2862 468
rect 2844 468 2862 486
rect 2844 486 2862 504
rect 2844 504 2862 522
rect 2844 522 2862 540
rect 2844 540 2862 558
rect 2844 558 2862 576
rect 2844 576 2862 594
rect 2844 594 2862 612
rect 2844 612 2862 630
rect 2844 630 2862 648
rect 2844 648 2862 666
rect 2844 666 2862 684
rect 2844 684 2862 702
rect 2844 702 2862 720
rect 2844 720 2862 738
rect 2844 918 2862 936
rect 2844 936 2862 954
rect 2844 954 2862 972
rect 2844 972 2862 990
rect 2844 990 2862 1008
rect 2844 1008 2862 1026
rect 2844 1026 2862 1044
rect 2844 1044 2862 1062
rect 2844 1062 2862 1080
rect 2844 1080 2862 1098
rect 2844 1098 2862 1116
rect 2844 1116 2862 1134
rect 2844 1458 2862 1476
rect 2844 1476 2862 1494
rect 2844 1494 2862 1512
rect 2844 1512 2862 1530
rect 2844 1530 2862 1548
rect 2844 1548 2862 1566
rect 2844 1566 2862 1584
rect 2844 1584 2862 1602
rect 2844 1602 2862 1620
rect 2844 1620 2862 1638
rect 2844 1638 2862 1656
rect 2844 1656 2862 1674
rect 2844 1674 2862 1692
rect 2844 1692 2862 1710
rect 2844 1710 2862 1728
rect 2844 1728 2862 1746
rect 2844 1746 2862 1764
rect 2844 1764 2862 1782
rect 2844 1782 2862 1800
rect 2844 1800 2862 1818
rect 2844 1818 2862 1836
rect 2844 1836 2862 1854
rect 2844 1854 2862 1872
rect 2844 1872 2862 1890
rect 2844 1890 2862 1908
rect 2844 1908 2862 1926
rect 2844 1926 2862 1944
rect 2844 1944 2862 1962
rect 2844 1962 2862 1980
rect 2844 1980 2862 1998
rect 2844 1998 2862 2016
rect 2844 2016 2862 2034
rect 2844 2034 2862 2052
rect 2844 2052 2862 2070
rect 2844 2070 2862 2088
rect 2844 2088 2862 2106
rect 2844 2106 2862 2124
rect 2844 2124 2862 2142
rect 2844 2142 2862 2160
rect 2844 2160 2862 2178
rect 2844 2178 2862 2196
rect 2844 2196 2862 2214
rect 2844 2214 2862 2232
rect 2844 2232 2862 2250
rect 2844 2250 2862 2268
rect 2844 2268 2862 2286
rect 2844 2286 2862 2304
rect 2844 2304 2862 2322
rect 2844 2322 2862 2340
rect 2844 2340 2862 2358
rect 2844 2358 2862 2376
rect 2844 2376 2862 2394
rect 2844 2394 2862 2412
rect 2844 2412 2862 2430
rect 2844 2430 2862 2448
rect 2844 2448 2862 2466
rect 2844 2466 2862 2484
rect 2844 2484 2862 2502
rect 2844 2502 2862 2520
rect 2844 2520 2862 2538
rect 2844 2538 2862 2556
rect 2844 2556 2862 2574
rect 2844 2574 2862 2592
rect 2844 2592 2862 2610
rect 2844 2610 2862 2628
rect 2844 2628 2862 2646
rect 2844 2646 2862 2664
rect 2844 2664 2862 2682
rect 2844 2682 2862 2700
rect 2844 2700 2862 2718
rect 2844 2718 2862 2736
rect 2844 2736 2862 2754
rect 2844 2754 2862 2772
rect 2844 2772 2862 2790
rect 2844 2790 2862 2808
rect 2844 6534 2862 6552
rect 2844 6552 2862 6570
rect 2844 6570 2862 6588
rect 2844 6588 2862 6606
rect 2844 6606 2862 6624
rect 2844 6624 2862 6642
rect 2844 6642 2862 6660
rect 2844 6660 2862 6678
rect 2844 6678 2862 6696
rect 2844 6696 2862 6714
rect 2844 6714 2862 6732
rect 2844 6732 2862 6750
rect 2844 6750 2862 6768
rect 2844 6768 2862 6786
rect 2844 6786 2862 6804
rect 2844 6804 2862 6822
rect 2844 6822 2862 6840
rect 2844 6840 2862 6858
rect 2844 6858 2862 6876
rect 2844 6876 2862 6894
rect 2844 6894 2862 6912
rect 2844 6912 2862 6930
rect 2844 6930 2862 6948
rect 2844 6948 2862 6966
rect 2844 6966 2862 6984
rect 2844 6984 2862 7002
rect 2844 7002 2862 7020
rect 2844 7020 2862 7038
rect 2844 7038 2862 7056
rect 2844 7056 2862 7074
rect 2844 7074 2862 7092
rect 2844 7092 2862 7110
rect 2844 7110 2862 7128
rect 2844 7128 2862 7146
rect 2844 7146 2862 7164
rect 2844 7164 2862 7182
rect 2862 90 2880 108
rect 2862 108 2880 126
rect 2862 126 2880 144
rect 2862 144 2880 162
rect 2862 162 2880 180
rect 2862 180 2880 198
rect 2862 198 2880 216
rect 2862 216 2880 234
rect 2862 234 2880 252
rect 2862 252 2880 270
rect 2862 270 2880 288
rect 2862 468 2880 486
rect 2862 486 2880 504
rect 2862 504 2880 522
rect 2862 522 2880 540
rect 2862 540 2880 558
rect 2862 558 2880 576
rect 2862 576 2880 594
rect 2862 594 2880 612
rect 2862 612 2880 630
rect 2862 630 2880 648
rect 2862 648 2880 666
rect 2862 666 2880 684
rect 2862 684 2880 702
rect 2862 702 2880 720
rect 2862 720 2880 738
rect 2862 936 2880 954
rect 2862 954 2880 972
rect 2862 972 2880 990
rect 2862 990 2880 1008
rect 2862 1008 2880 1026
rect 2862 1026 2880 1044
rect 2862 1044 2880 1062
rect 2862 1062 2880 1080
rect 2862 1080 2880 1098
rect 2862 1098 2880 1116
rect 2862 1116 2880 1134
rect 2862 1134 2880 1152
rect 2862 1152 2880 1170
rect 2862 1170 2880 1188
rect 2862 1494 2880 1512
rect 2862 1512 2880 1530
rect 2862 1530 2880 1548
rect 2862 1548 2880 1566
rect 2862 1566 2880 1584
rect 2862 1584 2880 1602
rect 2862 1602 2880 1620
rect 2862 1620 2880 1638
rect 2862 1638 2880 1656
rect 2862 1656 2880 1674
rect 2862 1674 2880 1692
rect 2862 1692 2880 1710
rect 2862 1710 2880 1728
rect 2862 1728 2880 1746
rect 2862 1746 2880 1764
rect 2862 1764 2880 1782
rect 2862 1782 2880 1800
rect 2862 1800 2880 1818
rect 2862 1818 2880 1836
rect 2862 1836 2880 1854
rect 2862 1854 2880 1872
rect 2862 1872 2880 1890
rect 2862 1890 2880 1908
rect 2862 1908 2880 1926
rect 2862 1926 2880 1944
rect 2862 1944 2880 1962
rect 2862 1962 2880 1980
rect 2862 1980 2880 1998
rect 2862 1998 2880 2016
rect 2862 2016 2880 2034
rect 2862 2034 2880 2052
rect 2862 2052 2880 2070
rect 2862 2070 2880 2088
rect 2862 2088 2880 2106
rect 2862 2106 2880 2124
rect 2862 2124 2880 2142
rect 2862 2142 2880 2160
rect 2862 2160 2880 2178
rect 2862 2178 2880 2196
rect 2862 2196 2880 2214
rect 2862 2214 2880 2232
rect 2862 2232 2880 2250
rect 2862 2250 2880 2268
rect 2862 2268 2880 2286
rect 2862 2286 2880 2304
rect 2862 2304 2880 2322
rect 2862 2322 2880 2340
rect 2862 2340 2880 2358
rect 2862 2358 2880 2376
rect 2862 2376 2880 2394
rect 2862 2394 2880 2412
rect 2862 2412 2880 2430
rect 2862 2430 2880 2448
rect 2862 2448 2880 2466
rect 2862 2466 2880 2484
rect 2862 2484 2880 2502
rect 2862 2502 2880 2520
rect 2862 2520 2880 2538
rect 2862 2538 2880 2556
rect 2862 2556 2880 2574
rect 2862 2574 2880 2592
rect 2862 2592 2880 2610
rect 2862 2610 2880 2628
rect 2862 2628 2880 2646
rect 2862 2646 2880 2664
rect 2862 2664 2880 2682
rect 2862 2682 2880 2700
rect 2862 2700 2880 2718
rect 2862 2718 2880 2736
rect 2862 2736 2880 2754
rect 2862 2754 2880 2772
rect 2862 2772 2880 2790
rect 2862 2790 2880 2808
rect 2862 2808 2880 2826
rect 2862 2826 2880 2844
rect 2862 2844 2880 2862
rect 2862 6552 2880 6570
rect 2862 6570 2880 6588
rect 2862 6588 2880 6606
rect 2862 6606 2880 6624
rect 2862 6624 2880 6642
rect 2862 6642 2880 6660
rect 2862 6660 2880 6678
rect 2862 6678 2880 6696
rect 2862 6696 2880 6714
rect 2862 6714 2880 6732
rect 2862 6732 2880 6750
rect 2862 6750 2880 6768
rect 2862 6768 2880 6786
rect 2862 6786 2880 6804
rect 2862 6804 2880 6822
rect 2862 6822 2880 6840
rect 2862 6840 2880 6858
rect 2862 6858 2880 6876
rect 2862 6876 2880 6894
rect 2862 6894 2880 6912
rect 2862 6912 2880 6930
rect 2862 6930 2880 6948
rect 2862 6948 2880 6966
rect 2862 6966 2880 6984
rect 2862 6984 2880 7002
rect 2862 7002 2880 7020
rect 2862 7020 2880 7038
rect 2862 7038 2880 7056
rect 2862 7056 2880 7074
rect 2862 7074 2880 7092
rect 2862 7092 2880 7110
rect 2862 7110 2880 7128
rect 2862 7128 2880 7146
rect 2862 7146 2880 7164
rect 2862 7164 2880 7182
rect 2880 90 2898 108
rect 2880 108 2898 126
rect 2880 126 2898 144
rect 2880 144 2898 162
rect 2880 162 2898 180
rect 2880 180 2898 198
rect 2880 198 2898 216
rect 2880 216 2898 234
rect 2880 234 2898 252
rect 2880 252 2898 270
rect 2880 270 2898 288
rect 2880 288 2898 306
rect 2880 486 2898 504
rect 2880 504 2898 522
rect 2880 522 2898 540
rect 2880 540 2898 558
rect 2880 558 2898 576
rect 2880 576 2898 594
rect 2880 594 2898 612
rect 2880 612 2898 630
rect 2880 630 2898 648
rect 2880 648 2898 666
rect 2880 666 2898 684
rect 2880 684 2898 702
rect 2880 702 2898 720
rect 2880 720 2898 738
rect 2880 738 2898 756
rect 2880 954 2898 972
rect 2880 972 2898 990
rect 2880 990 2898 1008
rect 2880 1008 2898 1026
rect 2880 1026 2898 1044
rect 2880 1044 2898 1062
rect 2880 1062 2898 1080
rect 2880 1080 2898 1098
rect 2880 1098 2898 1116
rect 2880 1116 2898 1134
rect 2880 1134 2898 1152
rect 2880 1152 2898 1170
rect 2880 1170 2898 1188
rect 2880 1188 2898 1206
rect 2880 1206 2898 1224
rect 2880 1530 2898 1548
rect 2880 1548 2898 1566
rect 2880 1566 2898 1584
rect 2880 1584 2898 1602
rect 2880 1602 2898 1620
rect 2880 1620 2898 1638
rect 2880 1638 2898 1656
rect 2880 1656 2898 1674
rect 2880 1674 2898 1692
rect 2880 1692 2898 1710
rect 2880 1710 2898 1728
rect 2880 1728 2898 1746
rect 2880 1746 2898 1764
rect 2880 1764 2898 1782
rect 2880 1782 2898 1800
rect 2880 1800 2898 1818
rect 2880 1818 2898 1836
rect 2880 1836 2898 1854
rect 2880 1854 2898 1872
rect 2880 1872 2898 1890
rect 2880 1890 2898 1908
rect 2880 1908 2898 1926
rect 2880 1926 2898 1944
rect 2880 1944 2898 1962
rect 2880 1962 2898 1980
rect 2880 1980 2898 1998
rect 2880 1998 2898 2016
rect 2880 2016 2898 2034
rect 2880 2034 2898 2052
rect 2880 2052 2898 2070
rect 2880 2070 2898 2088
rect 2880 2088 2898 2106
rect 2880 2106 2898 2124
rect 2880 2124 2898 2142
rect 2880 2142 2898 2160
rect 2880 2160 2898 2178
rect 2880 2178 2898 2196
rect 2880 2196 2898 2214
rect 2880 2214 2898 2232
rect 2880 2232 2898 2250
rect 2880 2250 2898 2268
rect 2880 2268 2898 2286
rect 2880 2286 2898 2304
rect 2880 2304 2898 2322
rect 2880 2322 2898 2340
rect 2880 2340 2898 2358
rect 2880 2358 2898 2376
rect 2880 2376 2898 2394
rect 2880 2394 2898 2412
rect 2880 2412 2898 2430
rect 2880 2430 2898 2448
rect 2880 2448 2898 2466
rect 2880 2466 2898 2484
rect 2880 2484 2898 2502
rect 2880 2502 2898 2520
rect 2880 2520 2898 2538
rect 2880 2538 2898 2556
rect 2880 2556 2898 2574
rect 2880 2574 2898 2592
rect 2880 2592 2898 2610
rect 2880 2610 2898 2628
rect 2880 2628 2898 2646
rect 2880 2646 2898 2664
rect 2880 2664 2898 2682
rect 2880 2682 2898 2700
rect 2880 2700 2898 2718
rect 2880 2718 2898 2736
rect 2880 2736 2898 2754
rect 2880 2754 2898 2772
rect 2880 2772 2898 2790
rect 2880 2790 2898 2808
rect 2880 2808 2898 2826
rect 2880 2826 2898 2844
rect 2880 2844 2898 2862
rect 2880 2862 2898 2880
rect 2880 2880 2898 2898
rect 2880 2898 2898 2916
rect 2880 2916 2898 2934
rect 2880 6552 2898 6570
rect 2880 6570 2898 6588
rect 2880 6588 2898 6606
rect 2880 6606 2898 6624
rect 2880 6624 2898 6642
rect 2880 6642 2898 6660
rect 2880 6660 2898 6678
rect 2880 6678 2898 6696
rect 2880 6696 2898 6714
rect 2880 6714 2898 6732
rect 2880 6732 2898 6750
rect 2880 6750 2898 6768
rect 2880 6768 2898 6786
rect 2880 6786 2898 6804
rect 2880 6804 2898 6822
rect 2880 6822 2898 6840
rect 2880 6840 2898 6858
rect 2880 6858 2898 6876
rect 2880 6876 2898 6894
rect 2880 6894 2898 6912
rect 2880 6912 2898 6930
rect 2880 6930 2898 6948
rect 2880 6948 2898 6966
rect 2880 6966 2898 6984
rect 2880 6984 2898 7002
rect 2880 7002 2898 7020
rect 2880 7020 2898 7038
rect 2880 7038 2898 7056
rect 2880 7056 2898 7074
rect 2880 7074 2898 7092
rect 2880 7092 2898 7110
rect 2880 7110 2898 7128
rect 2880 7128 2898 7146
rect 2880 7146 2898 7164
rect 2880 7164 2898 7182
rect 2880 7182 2898 7200
rect 2898 90 2916 108
rect 2898 108 2916 126
rect 2898 126 2916 144
rect 2898 144 2916 162
rect 2898 162 2916 180
rect 2898 180 2916 198
rect 2898 198 2916 216
rect 2898 216 2916 234
rect 2898 234 2916 252
rect 2898 252 2916 270
rect 2898 270 2916 288
rect 2898 288 2916 306
rect 2898 306 2916 324
rect 2898 486 2916 504
rect 2898 504 2916 522
rect 2898 522 2916 540
rect 2898 540 2916 558
rect 2898 558 2916 576
rect 2898 576 2916 594
rect 2898 594 2916 612
rect 2898 612 2916 630
rect 2898 630 2916 648
rect 2898 648 2916 666
rect 2898 666 2916 684
rect 2898 684 2916 702
rect 2898 702 2916 720
rect 2898 720 2916 738
rect 2898 738 2916 756
rect 2898 756 2916 774
rect 2898 954 2916 972
rect 2898 972 2916 990
rect 2898 990 2916 1008
rect 2898 1008 2916 1026
rect 2898 1026 2916 1044
rect 2898 1044 2916 1062
rect 2898 1062 2916 1080
rect 2898 1080 2916 1098
rect 2898 1098 2916 1116
rect 2898 1116 2916 1134
rect 2898 1134 2916 1152
rect 2898 1152 2916 1170
rect 2898 1170 2916 1188
rect 2898 1188 2916 1206
rect 2898 1206 2916 1224
rect 2898 1224 2916 1242
rect 2898 1242 2916 1260
rect 2898 1566 2916 1584
rect 2898 1584 2916 1602
rect 2898 1602 2916 1620
rect 2898 1620 2916 1638
rect 2898 1638 2916 1656
rect 2898 1656 2916 1674
rect 2898 1674 2916 1692
rect 2898 1692 2916 1710
rect 2898 1710 2916 1728
rect 2898 1728 2916 1746
rect 2898 1746 2916 1764
rect 2898 1764 2916 1782
rect 2898 1782 2916 1800
rect 2898 1800 2916 1818
rect 2898 1818 2916 1836
rect 2898 1836 2916 1854
rect 2898 1854 2916 1872
rect 2898 1872 2916 1890
rect 2898 1890 2916 1908
rect 2898 1908 2916 1926
rect 2898 1926 2916 1944
rect 2898 1944 2916 1962
rect 2898 1962 2916 1980
rect 2898 1980 2916 1998
rect 2898 1998 2916 2016
rect 2898 2016 2916 2034
rect 2898 2034 2916 2052
rect 2898 2052 2916 2070
rect 2898 2070 2916 2088
rect 2898 2088 2916 2106
rect 2898 2106 2916 2124
rect 2898 2124 2916 2142
rect 2898 2142 2916 2160
rect 2898 2160 2916 2178
rect 2898 2178 2916 2196
rect 2898 2196 2916 2214
rect 2898 2214 2916 2232
rect 2898 2232 2916 2250
rect 2898 2250 2916 2268
rect 2898 2268 2916 2286
rect 2898 2286 2916 2304
rect 2898 2304 2916 2322
rect 2898 2322 2916 2340
rect 2898 2340 2916 2358
rect 2898 2358 2916 2376
rect 2898 2376 2916 2394
rect 2898 2394 2916 2412
rect 2898 2412 2916 2430
rect 2898 2430 2916 2448
rect 2898 2448 2916 2466
rect 2898 2466 2916 2484
rect 2898 2484 2916 2502
rect 2898 2502 2916 2520
rect 2898 2520 2916 2538
rect 2898 2538 2916 2556
rect 2898 2556 2916 2574
rect 2898 2574 2916 2592
rect 2898 2592 2916 2610
rect 2898 2610 2916 2628
rect 2898 2628 2916 2646
rect 2898 2646 2916 2664
rect 2898 2664 2916 2682
rect 2898 2682 2916 2700
rect 2898 2700 2916 2718
rect 2898 2718 2916 2736
rect 2898 2736 2916 2754
rect 2898 2754 2916 2772
rect 2898 2772 2916 2790
rect 2898 2790 2916 2808
rect 2898 2808 2916 2826
rect 2898 2826 2916 2844
rect 2898 2844 2916 2862
rect 2898 2862 2916 2880
rect 2898 2880 2916 2898
rect 2898 2898 2916 2916
rect 2898 2916 2916 2934
rect 2898 2934 2916 2952
rect 2898 2952 2916 2970
rect 2898 2970 2916 2988
rect 2898 6552 2916 6570
rect 2898 6570 2916 6588
rect 2898 6588 2916 6606
rect 2898 6606 2916 6624
rect 2898 6624 2916 6642
rect 2898 6642 2916 6660
rect 2898 6660 2916 6678
rect 2898 6678 2916 6696
rect 2898 6696 2916 6714
rect 2898 6714 2916 6732
rect 2898 6732 2916 6750
rect 2898 6750 2916 6768
rect 2898 6768 2916 6786
rect 2898 6786 2916 6804
rect 2898 6804 2916 6822
rect 2898 6822 2916 6840
rect 2898 6840 2916 6858
rect 2898 6858 2916 6876
rect 2898 6876 2916 6894
rect 2898 6894 2916 6912
rect 2898 6912 2916 6930
rect 2898 6930 2916 6948
rect 2898 6948 2916 6966
rect 2898 6966 2916 6984
rect 2898 6984 2916 7002
rect 2898 7002 2916 7020
rect 2898 7020 2916 7038
rect 2898 7038 2916 7056
rect 2898 7056 2916 7074
rect 2898 7074 2916 7092
rect 2898 7092 2916 7110
rect 2898 7110 2916 7128
rect 2898 7128 2916 7146
rect 2898 7146 2916 7164
rect 2898 7164 2916 7182
rect 2898 7182 2916 7200
rect 2916 90 2934 108
rect 2916 108 2934 126
rect 2916 126 2934 144
rect 2916 144 2934 162
rect 2916 162 2934 180
rect 2916 180 2934 198
rect 2916 198 2934 216
rect 2916 216 2934 234
rect 2916 234 2934 252
rect 2916 252 2934 270
rect 2916 270 2934 288
rect 2916 288 2934 306
rect 2916 306 2934 324
rect 2916 324 2934 342
rect 2916 504 2934 522
rect 2916 522 2934 540
rect 2916 540 2934 558
rect 2916 558 2934 576
rect 2916 576 2934 594
rect 2916 594 2934 612
rect 2916 612 2934 630
rect 2916 630 2934 648
rect 2916 648 2934 666
rect 2916 666 2934 684
rect 2916 684 2934 702
rect 2916 702 2934 720
rect 2916 720 2934 738
rect 2916 738 2934 756
rect 2916 756 2934 774
rect 2916 774 2934 792
rect 2916 972 2934 990
rect 2916 990 2934 1008
rect 2916 1008 2934 1026
rect 2916 1026 2934 1044
rect 2916 1044 2934 1062
rect 2916 1062 2934 1080
rect 2916 1080 2934 1098
rect 2916 1098 2934 1116
rect 2916 1116 2934 1134
rect 2916 1134 2934 1152
rect 2916 1152 2934 1170
rect 2916 1170 2934 1188
rect 2916 1188 2934 1206
rect 2916 1206 2934 1224
rect 2916 1224 2934 1242
rect 2916 1242 2934 1260
rect 2916 1260 2934 1278
rect 2916 1278 2934 1296
rect 2916 1296 2934 1314
rect 2916 1602 2934 1620
rect 2916 1620 2934 1638
rect 2916 1638 2934 1656
rect 2916 1656 2934 1674
rect 2916 1674 2934 1692
rect 2916 1692 2934 1710
rect 2916 1710 2934 1728
rect 2916 1728 2934 1746
rect 2916 1746 2934 1764
rect 2916 1764 2934 1782
rect 2916 1782 2934 1800
rect 2916 1800 2934 1818
rect 2916 1818 2934 1836
rect 2916 1836 2934 1854
rect 2916 1854 2934 1872
rect 2916 1872 2934 1890
rect 2916 1890 2934 1908
rect 2916 1908 2934 1926
rect 2916 1926 2934 1944
rect 2916 1944 2934 1962
rect 2916 1962 2934 1980
rect 2916 1980 2934 1998
rect 2916 1998 2934 2016
rect 2916 2016 2934 2034
rect 2916 2034 2934 2052
rect 2916 2052 2934 2070
rect 2916 2070 2934 2088
rect 2916 2088 2934 2106
rect 2916 2106 2934 2124
rect 2916 2124 2934 2142
rect 2916 2142 2934 2160
rect 2916 2160 2934 2178
rect 2916 2178 2934 2196
rect 2916 2196 2934 2214
rect 2916 2214 2934 2232
rect 2916 2232 2934 2250
rect 2916 2250 2934 2268
rect 2916 2268 2934 2286
rect 2916 2286 2934 2304
rect 2916 2304 2934 2322
rect 2916 2322 2934 2340
rect 2916 2340 2934 2358
rect 2916 2358 2934 2376
rect 2916 2376 2934 2394
rect 2916 2394 2934 2412
rect 2916 2412 2934 2430
rect 2916 2430 2934 2448
rect 2916 2448 2934 2466
rect 2916 2466 2934 2484
rect 2916 2484 2934 2502
rect 2916 2502 2934 2520
rect 2916 2520 2934 2538
rect 2916 2538 2934 2556
rect 2916 2556 2934 2574
rect 2916 2574 2934 2592
rect 2916 2592 2934 2610
rect 2916 2610 2934 2628
rect 2916 2628 2934 2646
rect 2916 2646 2934 2664
rect 2916 2664 2934 2682
rect 2916 2682 2934 2700
rect 2916 2700 2934 2718
rect 2916 2718 2934 2736
rect 2916 2736 2934 2754
rect 2916 2754 2934 2772
rect 2916 2772 2934 2790
rect 2916 2790 2934 2808
rect 2916 2808 2934 2826
rect 2916 2826 2934 2844
rect 2916 2844 2934 2862
rect 2916 2862 2934 2880
rect 2916 2880 2934 2898
rect 2916 2898 2934 2916
rect 2916 2916 2934 2934
rect 2916 2934 2934 2952
rect 2916 2952 2934 2970
rect 2916 2970 2934 2988
rect 2916 2988 2934 3006
rect 2916 3006 2934 3024
rect 2916 3024 2934 3042
rect 2916 3042 2934 3060
rect 2916 6552 2934 6570
rect 2916 6570 2934 6588
rect 2916 6588 2934 6606
rect 2916 6606 2934 6624
rect 2916 6624 2934 6642
rect 2916 6642 2934 6660
rect 2916 6660 2934 6678
rect 2916 6678 2934 6696
rect 2916 6696 2934 6714
rect 2916 6714 2934 6732
rect 2916 6732 2934 6750
rect 2916 6750 2934 6768
rect 2916 6768 2934 6786
rect 2916 6786 2934 6804
rect 2916 6804 2934 6822
rect 2916 6822 2934 6840
rect 2916 6840 2934 6858
rect 2916 6858 2934 6876
rect 2916 6876 2934 6894
rect 2916 6894 2934 6912
rect 2916 6912 2934 6930
rect 2916 6930 2934 6948
rect 2916 6948 2934 6966
rect 2916 6966 2934 6984
rect 2916 6984 2934 7002
rect 2916 7002 2934 7020
rect 2916 7020 2934 7038
rect 2916 7038 2934 7056
rect 2916 7056 2934 7074
rect 2916 7074 2934 7092
rect 2916 7092 2934 7110
rect 2916 7110 2934 7128
rect 2916 7128 2934 7146
rect 2916 7146 2934 7164
rect 2916 7164 2934 7182
rect 2916 7182 2934 7200
rect 2934 90 2952 108
rect 2934 108 2952 126
rect 2934 126 2952 144
rect 2934 144 2952 162
rect 2934 162 2952 180
rect 2934 180 2952 198
rect 2934 198 2952 216
rect 2934 216 2952 234
rect 2934 234 2952 252
rect 2934 252 2952 270
rect 2934 270 2952 288
rect 2934 288 2952 306
rect 2934 306 2952 324
rect 2934 324 2952 342
rect 2934 522 2952 540
rect 2934 540 2952 558
rect 2934 558 2952 576
rect 2934 576 2952 594
rect 2934 594 2952 612
rect 2934 612 2952 630
rect 2934 630 2952 648
rect 2934 648 2952 666
rect 2934 666 2952 684
rect 2934 684 2952 702
rect 2934 702 2952 720
rect 2934 720 2952 738
rect 2934 738 2952 756
rect 2934 756 2952 774
rect 2934 774 2952 792
rect 2934 792 2952 810
rect 2934 990 2952 1008
rect 2934 1008 2952 1026
rect 2934 1026 2952 1044
rect 2934 1044 2952 1062
rect 2934 1062 2952 1080
rect 2934 1080 2952 1098
rect 2934 1098 2952 1116
rect 2934 1116 2952 1134
rect 2934 1134 2952 1152
rect 2934 1152 2952 1170
rect 2934 1170 2952 1188
rect 2934 1188 2952 1206
rect 2934 1206 2952 1224
rect 2934 1224 2952 1242
rect 2934 1242 2952 1260
rect 2934 1260 2952 1278
rect 2934 1278 2952 1296
rect 2934 1296 2952 1314
rect 2934 1314 2952 1332
rect 2934 1332 2952 1350
rect 2934 1638 2952 1656
rect 2934 1656 2952 1674
rect 2934 1674 2952 1692
rect 2934 1692 2952 1710
rect 2934 1710 2952 1728
rect 2934 1728 2952 1746
rect 2934 1746 2952 1764
rect 2934 1764 2952 1782
rect 2934 1782 2952 1800
rect 2934 1800 2952 1818
rect 2934 1818 2952 1836
rect 2934 1836 2952 1854
rect 2934 1854 2952 1872
rect 2934 1872 2952 1890
rect 2934 1890 2952 1908
rect 2934 1908 2952 1926
rect 2934 1926 2952 1944
rect 2934 1944 2952 1962
rect 2934 1962 2952 1980
rect 2934 1980 2952 1998
rect 2934 1998 2952 2016
rect 2934 2016 2952 2034
rect 2934 2034 2952 2052
rect 2934 2052 2952 2070
rect 2934 2070 2952 2088
rect 2934 2088 2952 2106
rect 2934 2106 2952 2124
rect 2934 2124 2952 2142
rect 2934 2142 2952 2160
rect 2934 2160 2952 2178
rect 2934 2178 2952 2196
rect 2934 2196 2952 2214
rect 2934 2214 2952 2232
rect 2934 2232 2952 2250
rect 2934 2250 2952 2268
rect 2934 2268 2952 2286
rect 2934 2286 2952 2304
rect 2934 2304 2952 2322
rect 2934 2322 2952 2340
rect 2934 2340 2952 2358
rect 2934 2358 2952 2376
rect 2934 2376 2952 2394
rect 2934 2394 2952 2412
rect 2934 2412 2952 2430
rect 2934 2430 2952 2448
rect 2934 2448 2952 2466
rect 2934 2466 2952 2484
rect 2934 2484 2952 2502
rect 2934 2502 2952 2520
rect 2934 2520 2952 2538
rect 2934 2538 2952 2556
rect 2934 2556 2952 2574
rect 2934 2574 2952 2592
rect 2934 2592 2952 2610
rect 2934 2610 2952 2628
rect 2934 2628 2952 2646
rect 2934 2646 2952 2664
rect 2934 2664 2952 2682
rect 2934 2682 2952 2700
rect 2934 2700 2952 2718
rect 2934 2718 2952 2736
rect 2934 2736 2952 2754
rect 2934 2754 2952 2772
rect 2934 2772 2952 2790
rect 2934 2790 2952 2808
rect 2934 2808 2952 2826
rect 2934 2826 2952 2844
rect 2934 2844 2952 2862
rect 2934 2862 2952 2880
rect 2934 2880 2952 2898
rect 2934 2898 2952 2916
rect 2934 2916 2952 2934
rect 2934 2934 2952 2952
rect 2934 2952 2952 2970
rect 2934 2970 2952 2988
rect 2934 2988 2952 3006
rect 2934 3006 2952 3024
rect 2934 3024 2952 3042
rect 2934 3042 2952 3060
rect 2934 3060 2952 3078
rect 2934 3078 2952 3096
rect 2934 3096 2952 3114
rect 2934 6570 2952 6588
rect 2934 6588 2952 6606
rect 2934 6606 2952 6624
rect 2934 6624 2952 6642
rect 2934 6642 2952 6660
rect 2934 6660 2952 6678
rect 2934 6678 2952 6696
rect 2934 6696 2952 6714
rect 2934 6714 2952 6732
rect 2934 6732 2952 6750
rect 2934 6750 2952 6768
rect 2934 6768 2952 6786
rect 2934 6786 2952 6804
rect 2934 6804 2952 6822
rect 2934 6822 2952 6840
rect 2934 6840 2952 6858
rect 2934 6858 2952 6876
rect 2934 6876 2952 6894
rect 2934 6894 2952 6912
rect 2934 6912 2952 6930
rect 2934 6930 2952 6948
rect 2934 6948 2952 6966
rect 2934 6966 2952 6984
rect 2934 6984 2952 7002
rect 2934 7002 2952 7020
rect 2934 7020 2952 7038
rect 2934 7038 2952 7056
rect 2934 7056 2952 7074
rect 2934 7074 2952 7092
rect 2934 7092 2952 7110
rect 2934 7110 2952 7128
rect 2934 7128 2952 7146
rect 2934 7146 2952 7164
rect 2934 7164 2952 7182
rect 2934 7182 2952 7200
rect 2952 90 2970 108
rect 2952 108 2970 126
rect 2952 126 2970 144
rect 2952 144 2970 162
rect 2952 162 2970 180
rect 2952 180 2970 198
rect 2952 198 2970 216
rect 2952 216 2970 234
rect 2952 234 2970 252
rect 2952 252 2970 270
rect 2952 270 2970 288
rect 2952 288 2970 306
rect 2952 306 2970 324
rect 2952 324 2970 342
rect 2952 342 2970 360
rect 2952 540 2970 558
rect 2952 558 2970 576
rect 2952 576 2970 594
rect 2952 594 2970 612
rect 2952 612 2970 630
rect 2952 630 2970 648
rect 2952 648 2970 666
rect 2952 666 2970 684
rect 2952 684 2970 702
rect 2952 702 2970 720
rect 2952 720 2970 738
rect 2952 738 2970 756
rect 2952 756 2970 774
rect 2952 774 2970 792
rect 2952 792 2970 810
rect 2952 810 2970 828
rect 2952 1008 2970 1026
rect 2952 1026 2970 1044
rect 2952 1044 2970 1062
rect 2952 1062 2970 1080
rect 2952 1080 2970 1098
rect 2952 1098 2970 1116
rect 2952 1116 2970 1134
rect 2952 1134 2970 1152
rect 2952 1152 2970 1170
rect 2952 1170 2970 1188
rect 2952 1188 2970 1206
rect 2952 1206 2970 1224
rect 2952 1224 2970 1242
rect 2952 1242 2970 1260
rect 2952 1260 2970 1278
rect 2952 1278 2970 1296
rect 2952 1296 2970 1314
rect 2952 1314 2970 1332
rect 2952 1332 2970 1350
rect 2952 1350 2970 1368
rect 2952 1368 2970 1386
rect 2952 1674 2970 1692
rect 2952 1692 2970 1710
rect 2952 1710 2970 1728
rect 2952 1728 2970 1746
rect 2952 1746 2970 1764
rect 2952 1764 2970 1782
rect 2952 1782 2970 1800
rect 2952 1800 2970 1818
rect 2952 1818 2970 1836
rect 2952 1836 2970 1854
rect 2952 1854 2970 1872
rect 2952 1872 2970 1890
rect 2952 1890 2970 1908
rect 2952 1908 2970 1926
rect 2952 1926 2970 1944
rect 2952 1944 2970 1962
rect 2952 1962 2970 1980
rect 2952 1980 2970 1998
rect 2952 1998 2970 2016
rect 2952 2016 2970 2034
rect 2952 2034 2970 2052
rect 2952 2052 2970 2070
rect 2952 2070 2970 2088
rect 2952 2088 2970 2106
rect 2952 2106 2970 2124
rect 2952 2124 2970 2142
rect 2952 2142 2970 2160
rect 2952 2160 2970 2178
rect 2952 2178 2970 2196
rect 2952 2196 2970 2214
rect 2952 2214 2970 2232
rect 2952 2232 2970 2250
rect 2952 2250 2970 2268
rect 2952 2268 2970 2286
rect 2952 2286 2970 2304
rect 2952 2304 2970 2322
rect 2952 2322 2970 2340
rect 2952 2340 2970 2358
rect 2952 2358 2970 2376
rect 2952 2376 2970 2394
rect 2952 2394 2970 2412
rect 2952 2412 2970 2430
rect 2952 2430 2970 2448
rect 2952 2448 2970 2466
rect 2952 2466 2970 2484
rect 2952 2484 2970 2502
rect 2952 2502 2970 2520
rect 2952 2520 2970 2538
rect 2952 2538 2970 2556
rect 2952 2556 2970 2574
rect 2952 2574 2970 2592
rect 2952 2592 2970 2610
rect 2952 2610 2970 2628
rect 2952 2628 2970 2646
rect 2952 2646 2970 2664
rect 2952 2664 2970 2682
rect 2952 2682 2970 2700
rect 2952 2700 2970 2718
rect 2952 2718 2970 2736
rect 2952 2736 2970 2754
rect 2952 2754 2970 2772
rect 2952 2772 2970 2790
rect 2952 2790 2970 2808
rect 2952 2808 2970 2826
rect 2952 2826 2970 2844
rect 2952 2844 2970 2862
rect 2952 2862 2970 2880
rect 2952 2880 2970 2898
rect 2952 2898 2970 2916
rect 2952 2916 2970 2934
rect 2952 2934 2970 2952
rect 2952 2952 2970 2970
rect 2952 2970 2970 2988
rect 2952 2988 2970 3006
rect 2952 3006 2970 3024
rect 2952 3024 2970 3042
rect 2952 3042 2970 3060
rect 2952 3060 2970 3078
rect 2952 3078 2970 3096
rect 2952 3096 2970 3114
rect 2952 3114 2970 3132
rect 2952 3132 2970 3150
rect 2952 3150 2970 3168
rect 2952 3168 2970 3186
rect 2952 6570 2970 6588
rect 2952 6588 2970 6606
rect 2952 6606 2970 6624
rect 2952 6624 2970 6642
rect 2952 6642 2970 6660
rect 2952 6660 2970 6678
rect 2952 6678 2970 6696
rect 2952 6696 2970 6714
rect 2952 6714 2970 6732
rect 2952 6732 2970 6750
rect 2952 6750 2970 6768
rect 2952 6768 2970 6786
rect 2952 6786 2970 6804
rect 2952 6804 2970 6822
rect 2952 6822 2970 6840
rect 2952 6840 2970 6858
rect 2952 6858 2970 6876
rect 2952 6876 2970 6894
rect 2952 6894 2970 6912
rect 2952 6912 2970 6930
rect 2952 6930 2970 6948
rect 2952 6948 2970 6966
rect 2952 6966 2970 6984
rect 2952 6984 2970 7002
rect 2952 7002 2970 7020
rect 2952 7020 2970 7038
rect 2952 7038 2970 7056
rect 2952 7056 2970 7074
rect 2952 7074 2970 7092
rect 2952 7092 2970 7110
rect 2952 7110 2970 7128
rect 2952 7128 2970 7146
rect 2952 7146 2970 7164
rect 2952 7164 2970 7182
rect 2952 7182 2970 7200
rect 2970 90 2988 108
rect 2970 108 2988 126
rect 2970 126 2988 144
rect 2970 144 2988 162
rect 2970 162 2988 180
rect 2970 180 2988 198
rect 2970 198 2988 216
rect 2970 216 2988 234
rect 2970 234 2988 252
rect 2970 252 2988 270
rect 2970 270 2988 288
rect 2970 288 2988 306
rect 2970 306 2988 324
rect 2970 324 2988 342
rect 2970 342 2988 360
rect 2970 360 2988 378
rect 2970 540 2988 558
rect 2970 558 2988 576
rect 2970 576 2988 594
rect 2970 594 2988 612
rect 2970 612 2988 630
rect 2970 630 2988 648
rect 2970 648 2988 666
rect 2970 666 2988 684
rect 2970 684 2988 702
rect 2970 702 2988 720
rect 2970 720 2988 738
rect 2970 738 2988 756
rect 2970 756 2988 774
rect 2970 774 2988 792
rect 2970 792 2988 810
rect 2970 810 2988 828
rect 2970 1008 2988 1026
rect 2970 1026 2988 1044
rect 2970 1044 2988 1062
rect 2970 1062 2988 1080
rect 2970 1080 2988 1098
rect 2970 1098 2988 1116
rect 2970 1116 2988 1134
rect 2970 1134 2988 1152
rect 2970 1152 2988 1170
rect 2970 1170 2988 1188
rect 2970 1188 2988 1206
rect 2970 1206 2988 1224
rect 2970 1224 2988 1242
rect 2970 1242 2988 1260
rect 2970 1260 2988 1278
rect 2970 1278 2988 1296
rect 2970 1296 2988 1314
rect 2970 1314 2988 1332
rect 2970 1332 2988 1350
rect 2970 1350 2988 1368
rect 2970 1368 2988 1386
rect 2970 1386 2988 1404
rect 2970 1404 2988 1422
rect 2970 1710 2988 1728
rect 2970 1728 2988 1746
rect 2970 1746 2988 1764
rect 2970 1764 2988 1782
rect 2970 1782 2988 1800
rect 2970 1800 2988 1818
rect 2970 1818 2988 1836
rect 2970 1836 2988 1854
rect 2970 1854 2988 1872
rect 2970 1872 2988 1890
rect 2970 1890 2988 1908
rect 2970 1908 2988 1926
rect 2970 1926 2988 1944
rect 2970 1944 2988 1962
rect 2970 1962 2988 1980
rect 2970 1980 2988 1998
rect 2970 1998 2988 2016
rect 2970 2016 2988 2034
rect 2970 2034 2988 2052
rect 2970 2052 2988 2070
rect 2970 2070 2988 2088
rect 2970 2088 2988 2106
rect 2970 2106 2988 2124
rect 2970 2124 2988 2142
rect 2970 2142 2988 2160
rect 2970 2160 2988 2178
rect 2970 2178 2988 2196
rect 2970 2196 2988 2214
rect 2970 2214 2988 2232
rect 2970 2232 2988 2250
rect 2970 2250 2988 2268
rect 2970 2268 2988 2286
rect 2970 2286 2988 2304
rect 2970 2304 2988 2322
rect 2970 2322 2988 2340
rect 2970 2340 2988 2358
rect 2970 2358 2988 2376
rect 2970 2376 2988 2394
rect 2970 2394 2988 2412
rect 2970 2412 2988 2430
rect 2970 2430 2988 2448
rect 2970 2448 2988 2466
rect 2970 2466 2988 2484
rect 2970 2484 2988 2502
rect 2970 2502 2988 2520
rect 2970 2520 2988 2538
rect 2970 2538 2988 2556
rect 2970 2556 2988 2574
rect 2970 2574 2988 2592
rect 2970 2592 2988 2610
rect 2970 2610 2988 2628
rect 2970 2628 2988 2646
rect 2970 2646 2988 2664
rect 2970 2664 2988 2682
rect 2970 2682 2988 2700
rect 2970 2700 2988 2718
rect 2970 2718 2988 2736
rect 2970 2736 2988 2754
rect 2970 2754 2988 2772
rect 2970 2772 2988 2790
rect 2970 2790 2988 2808
rect 2970 2808 2988 2826
rect 2970 2826 2988 2844
rect 2970 2844 2988 2862
rect 2970 2862 2988 2880
rect 2970 2880 2988 2898
rect 2970 2898 2988 2916
rect 2970 2916 2988 2934
rect 2970 2934 2988 2952
rect 2970 2952 2988 2970
rect 2970 2970 2988 2988
rect 2970 2988 2988 3006
rect 2970 3006 2988 3024
rect 2970 3024 2988 3042
rect 2970 3042 2988 3060
rect 2970 3060 2988 3078
rect 2970 3078 2988 3096
rect 2970 3096 2988 3114
rect 2970 3114 2988 3132
rect 2970 3132 2988 3150
rect 2970 3150 2988 3168
rect 2970 3168 2988 3186
rect 2970 3186 2988 3204
rect 2970 3204 2988 3222
rect 2970 3222 2988 3240
rect 2970 6570 2988 6588
rect 2970 6588 2988 6606
rect 2970 6606 2988 6624
rect 2970 6624 2988 6642
rect 2970 6642 2988 6660
rect 2970 6660 2988 6678
rect 2970 6678 2988 6696
rect 2970 6696 2988 6714
rect 2970 6714 2988 6732
rect 2970 6732 2988 6750
rect 2970 6750 2988 6768
rect 2970 6768 2988 6786
rect 2970 6786 2988 6804
rect 2970 6804 2988 6822
rect 2970 6822 2988 6840
rect 2970 6840 2988 6858
rect 2970 6858 2988 6876
rect 2970 6876 2988 6894
rect 2970 6894 2988 6912
rect 2970 6912 2988 6930
rect 2970 6930 2988 6948
rect 2970 6948 2988 6966
rect 2970 6966 2988 6984
rect 2970 6984 2988 7002
rect 2970 7002 2988 7020
rect 2970 7020 2988 7038
rect 2970 7038 2988 7056
rect 2970 7056 2988 7074
rect 2970 7074 2988 7092
rect 2970 7092 2988 7110
rect 2970 7110 2988 7128
rect 2970 7128 2988 7146
rect 2970 7146 2988 7164
rect 2970 7164 2988 7182
rect 2970 7182 2988 7200
rect 2970 7200 2988 7218
rect 2988 72 3006 90
rect 2988 90 3006 108
rect 2988 108 3006 126
rect 2988 126 3006 144
rect 2988 144 3006 162
rect 2988 162 3006 180
rect 2988 180 3006 198
rect 2988 198 3006 216
rect 2988 216 3006 234
rect 2988 234 3006 252
rect 2988 252 3006 270
rect 2988 270 3006 288
rect 2988 288 3006 306
rect 2988 306 3006 324
rect 2988 324 3006 342
rect 2988 342 3006 360
rect 2988 360 3006 378
rect 2988 378 3006 396
rect 2988 558 3006 576
rect 2988 576 3006 594
rect 2988 594 3006 612
rect 2988 612 3006 630
rect 2988 630 3006 648
rect 2988 648 3006 666
rect 2988 666 3006 684
rect 2988 684 3006 702
rect 2988 702 3006 720
rect 2988 720 3006 738
rect 2988 738 3006 756
rect 2988 756 3006 774
rect 2988 774 3006 792
rect 2988 792 3006 810
rect 2988 810 3006 828
rect 2988 828 3006 846
rect 2988 1026 3006 1044
rect 2988 1044 3006 1062
rect 2988 1062 3006 1080
rect 2988 1080 3006 1098
rect 2988 1098 3006 1116
rect 2988 1116 3006 1134
rect 2988 1134 3006 1152
rect 2988 1152 3006 1170
rect 2988 1170 3006 1188
rect 2988 1188 3006 1206
rect 2988 1206 3006 1224
rect 2988 1224 3006 1242
rect 2988 1242 3006 1260
rect 2988 1260 3006 1278
rect 2988 1278 3006 1296
rect 2988 1296 3006 1314
rect 2988 1314 3006 1332
rect 2988 1332 3006 1350
rect 2988 1350 3006 1368
rect 2988 1368 3006 1386
rect 2988 1386 3006 1404
rect 2988 1404 3006 1422
rect 2988 1422 3006 1440
rect 2988 1440 3006 1458
rect 2988 1746 3006 1764
rect 2988 1764 3006 1782
rect 2988 1782 3006 1800
rect 2988 1800 3006 1818
rect 2988 1818 3006 1836
rect 2988 1836 3006 1854
rect 2988 1854 3006 1872
rect 2988 1872 3006 1890
rect 2988 1890 3006 1908
rect 2988 1908 3006 1926
rect 2988 1926 3006 1944
rect 2988 1944 3006 1962
rect 2988 1962 3006 1980
rect 2988 1980 3006 1998
rect 2988 1998 3006 2016
rect 2988 2016 3006 2034
rect 2988 2034 3006 2052
rect 2988 2052 3006 2070
rect 2988 2070 3006 2088
rect 2988 2088 3006 2106
rect 2988 2106 3006 2124
rect 2988 2124 3006 2142
rect 2988 2142 3006 2160
rect 2988 2160 3006 2178
rect 2988 2178 3006 2196
rect 2988 2196 3006 2214
rect 2988 2214 3006 2232
rect 2988 2232 3006 2250
rect 2988 2250 3006 2268
rect 2988 2268 3006 2286
rect 2988 2286 3006 2304
rect 2988 2304 3006 2322
rect 2988 2322 3006 2340
rect 2988 2340 3006 2358
rect 2988 2358 3006 2376
rect 2988 2376 3006 2394
rect 2988 2394 3006 2412
rect 2988 2412 3006 2430
rect 2988 2430 3006 2448
rect 2988 2448 3006 2466
rect 2988 2466 3006 2484
rect 2988 2484 3006 2502
rect 2988 2502 3006 2520
rect 2988 2520 3006 2538
rect 2988 2538 3006 2556
rect 2988 2556 3006 2574
rect 2988 2574 3006 2592
rect 2988 2592 3006 2610
rect 2988 2610 3006 2628
rect 2988 2628 3006 2646
rect 2988 2646 3006 2664
rect 2988 2664 3006 2682
rect 2988 2682 3006 2700
rect 2988 2700 3006 2718
rect 2988 2718 3006 2736
rect 2988 2736 3006 2754
rect 2988 2754 3006 2772
rect 2988 2772 3006 2790
rect 2988 2790 3006 2808
rect 2988 2808 3006 2826
rect 2988 2826 3006 2844
rect 2988 2844 3006 2862
rect 2988 2862 3006 2880
rect 2988 2880 3006 2898
rect 2988 2898 3006 2916
rect 2988 2916 3006 2934
rect 2988 2934 3006 2952
rect 2988 2952 3006 2970
rect 2988 2970 3006 2988
rect 2988 2988 3006 3006
rect 2988 3006 3006 3024
rect 2988 3024 3006 3042
rect 2988 3042 3006 3060
rect 2988 3060 3006 3078
rect 2988 3078 3006 3096
rect 2988 3096 3006 3114
rect 2988 3114 3006 3132
rect 2988 3132 3006 3150
rect 2988 3150 3006 3168
rect 2988 3168 3006 3186
rect 2988 3186 3006 3204
rect 2988 3204 3006 3222
rect 2988 3222 3006 3240
rect 2988 3240 3006 3258
rect 2988 3258 3006 3276
rect 2988 3276 3006 3294
rect 2988 3294 3006 3312
rect 2988 6570 3006 6588
rect 2988 6588 3006 6606
rect 2988 6606 3006 6624
rect 2988 6624 3006 6642
rect 2988 6642 3006 6660
rect 2988 6660 3006 6678
rect 2988 6678 3006 6696
rect 2988 6696 3006 6714
rect 2988 6714 3006 6732
rect 2988 6732 3006 6750
rect 2988 6750 3006 6768
rect 2988 6768 3006 6786
rect 2988 6786 3006 6804
rect 2988 6804 3006 6822
rect 2988 6822 3006 6840
rect 2988 6840 3006 6858
rect 2988 6858 3006 6876
rect 2988 6876 3006 6894
rect 2988 6894 3006 6912
rect 2988 6912 3006 6930
rect 2988 6930 3006 6948
rect 2988 6948 3006 6966
rect 2988 6966 3006 6984
rect 2988 6984 3006 7002
rect 2988 7002 3006 7020
rect 2988 7020 3006 7038
rect 2988 7038 3006 7056
rect 2988 7056 3006 7074
rect 2988 7074 3006 7092
rect 2988 7092 3006 7110
rect 2988 7110 3006 7128
rect 2988 7128 3006 7146
rect 2988 7146 3006 7164
rect 2988 7164 3006 7182
rect 2988 7182 3006 7200
rect 2988 7200 3006 7218
rect 3006 72 3024 90
rect 3006 90 3024 108
rect 3006 108 3024 126
rect 3006 126 3024 144
rect 3006 144 3024 162
rect 3006 162 3024 180
rect 3006 180 3024 198
rect 3006 198 3024 216
rect 3006 216 3024 234
rect 3006 234 3024 252
rect 3006 252 3024 270
rect 3006 270 3024 288
rect 3006 288 3024 306
rect 3006 306 3024 324
rect 3006 324 3024 342
rect 3006 342 3024 360
rect 3006 360 3024 378
rect 3006 378 3024 396
rect 3006 396 3024 414
rect 3006 576 3024 594
rect 3006 594 3024 612
rect 3006 612 3024 630
rect 3006 630 3024 648
rect 3006 648 3024 666
rect 3006 666 3024 684
rect 3006 684 3024 702
rect 3006 702 3024 720
rect 3006 720 3024 738
rect 3006 738 3024 756
rect 3006 756 3024 774
rect 3006 774 3024 792
rect 3006 792 3024 810
rect 3006 810 3024 828
rect 3006 828 3024 846
rect 3006 846 3024 864
rect 3006 1044 3024 1062
rect 3006 1062 3024 1080
rect 3006 1080 3024 1098
rect 3006 1098 3024 1116
rect 3006 1116 3024 1134
rect 3006 1134 3024 1152
rect 3006 1152 3024 1170
rect 3006 1170 3024 1188
rect 3006 1188 3024 1206
rect 3006 1206 3024 1224
rect 3006 1224 3024 1242
rect 3006 1242 3024 1260
rect 3006 1260 3024 1278
rect 3006 1278 3024 1296
rect 3006 1296 3024 1314
rect 3006 1314 3024 1332
rect 3006 1332 3024 1350
rect 3006 1350 3024 1368
rect 3006 1368 3024 1386
rect 3006 1386 3024 1404
rect 3006 1404 3024 1422
rect 3006 1422 3024 1440
rect 3006 1440 3024 1458
rect 3006 1458 3024 1476
rect 3006 1476 3024 1494
rect 3006 1764 3024 1782
rect 3006 1782 3024 1800
rect 3006 1800 3024 1818
rect 3006 1818 3024 1836
rect 3006 1836 3024 1854
rect 3006 1854 3024 1872
rect 3006 1872 3024 1890
rect 3006 1890 3024 1908
rect 3006 1908 3024 1926
rect 3006 1926 3024 1944
rect 3006 1944 3024 1962
rect 3006 1962 3024 1980
rect 3006 1980 3024 1998
rect 3006 1998 3024 2016
rect 3006 2016 3024 2034
rect 3006 2034 3024 2052
rect 3006 2052 3024 2070
rect 3006 2070 3024 2088
rect 3006 2088 3024 2106
rect 3006 2106 3024 2124
rect 3006 2124 3024 2142
rect 3006 2142 3024 2160
rect 3006 2160 3024 2178
rect 3006 2178 3024 2196
rect 3006 2196 3024 2214
rect 3006 2214 3024 2232
rect 3006 2232 3024 2250
rect 3006 2250 3024 2268
rect 3006 2268 3024 2286
rect 3006 2286 3024 2304
rect 3006 2304 3024 2322
rect 3006 2322 3024 2340
rect 3006 2340 3024 2358
rect 3006 2358 3024 2376
rect 3006 2376 3024 2394
rect 3006 2394 3024 2412
rect 3006 2412 3024 2430
rect 3006 2430 3024 2448
rect 3006 2448 3024 2466
rect 3006 2466 3024 2484
rect 3006 2484 3024 2502
rect 3006 2502 3024 2520
rect 3006 2520 3024 2538
rect 3006 2538 3024 2556
rect 3006 2556 3024 2574
rect 3006 2574 3024 2592
rect 3006 2592 3024 2610
rect 3006 2610 3024 2628
rect 3006 2628 3024 2646
rect 3006 2646 3024 2664
rect 3006 2664 3024 2682
rect 3006 2682 3024 2700
rect 3006 2700 3024 2718
rect 3006 2718 3024 2736
rect 3006 2736 3024 2754
rect 3006 2754 3024 2772
rect 3006 2772 3024 2790
rect 3006 2790 3024 2808
rect 3006 2808 3024 2826
rect 3006 2826 3024 2844
rect 3006 2844 3024 2862
rect 3006 2862 3024 2880
rect 3006 2880 3024 2898
rect 3006 2898 3024 2916
rect 3006 2916 3024 2934
rect 3006 2934 3024 2952
rect 3006 2952 3024 2970
rect 3006 2970 3024 2988
rect 3006 2988 3024 3006
rect 3006 3006 3024 3024
rect 3006 3024 3024 3042
rect 3006 3042 3024 3060
rect 3006 3060 3024 3078
rect 3006 3078 3024 3096
rect 3006 3096 3024 3114
rect 3006 3114 3024 3132
rect 3006 3132 3024 3150
rect 3006 3150 3024 3168
rect 3006 3168 3024 3186
rect 3006 3186 3024 3204
rect 3006 3204 3024 3222
rect 3006 3222 3024 3240
rect 3006 3240 3024 3258
rect 3006 3258 3024 3276
rect 3006 3276 3024 3294
rect 3006 3294 3024 3312
rect 3006 3312 3024 3330
rect 3006 3330 3024 3348
rect 3006 3348 3024 3366
rect 3006 6588 3024 6606
rect 3006 6606 3024 6624
rect 3006 6624 3024 6642
rect 3006 6642 3024 6660
rect 3006 6660 3024 6678
rect 3006 6678 3024 6696
rect 3006 6696 3024 6714
rect 3006 6714 3024 6732
rect 3006 6732 3024 6750
rect 3006 6750 3024 6768
rect 3006 6768 3024 6786
rect 3006 6786 3024 6804
rect 3006 6804 3024 6822
rect 3006 6822 3024 6840
rect 3006 6840 3024 6858
rect 3006 6858 3024 6876
rect 3006 6876 3024 6894
rect 3006 6894 3024 6912
rect 3006 6912 3024 6930
rect 3006 6930 3024 6948
rect 3006 6948 3024 6966
rect 3006 6966 3024 6984
rect 3006 6984 3024 7002
rect 3006 7002 3024 7020
rect 3006 7020 3024 7038
rect 3006 7038 3024 7056
rect 3006 7056 3024 7074
rect 3006 7074 3024 7092
rect 3006 7092 3024 7110
rect 3006 7110 3024 7128
rect 3006 7128 3024 7146
rect 3006 7146 3024 7164
rect 3006 7164 3024 7182
rect 3006 7182 3024 7200
rect 3006 7200 3024 7218
rect 3024 72 3042 90
rect 3024 90 3042 108
rect 3024 108 3042 126
rect 3024 126 3042 144
rect 3024 144 3042 162
rect 3024 162 3042 180
rect 3024 180 3042 198
rect 3024 198 3042 216
rect 3024 216 3042 234
rect 3024 234 3042 252
rect 3024 252 3042 270
rect 3024 270 3042 288
rect 3024 288 3042 306
rect 3024 306 3042 324
rect 3024 324 3042 342
rect 3024 342 3042 360
rect 3024 360 3042 378
rect 3024 378 3042 396
rect 3024 396 3042 414
rect 3024 576 3042 594
rect 3024 594 3042 612
rect 3024 612 3042 630
rect 3024 630 3042 648
rect 3024 648 3042 666
rect 3024 666 3042 684
rect 3024 684 3042 702
rect 3024 702 3042 720
rect 3024 720 3042 738
rect 3024 738 3042 756
rect 3024 756 3042 774
rect 3024 774 3042 792
rect 3024 792 3042 810
rect 3024 810 3042 828
rect 3024 828 3042 846
rect 3024 846 3042 864
rect 3024 864 3042 882
rect 3024 1062 3042 1080
rect 3024 1080 3042 1098
rect 3024 1098 3042 1116
rect 3024 1116 3042 1134
rect 3024 1134 3042 1152
rect 3024 1152 3042 1170
rect 3024 1170 3042 1188
rect 3024 1188 3042 1206
rect 3024 1206 3042 1224
rect 3024 1224 3042 1242
rect 3024 1242 3042 1260
rect 3024 1260 3042 1278
rect 3024 1278 3042 1296
rect 3024 1296 3042 1314
rect 3024 1314 3042 1332
rect 3024 1332 3042 1350
rect 3024 1350 3042 1368
rect 3024 1368 3042 1386
rect 3024 1386 3042 1404
rect 3024 1404 3042 1422
rect 3024 1422 3042 1440
rect 3024 1440 3042 1458
rect 3024 1458 3042 1476
rect 3024 1476 3042 1494
rect 3024 1494 3042 1512
rect 3024 1512 3042 1530
rect 3024 1800 3042 1818
rect 3024 1818 3042 1836
rect 3024 1836 3042 1854
rect 3024 1854 3042 1872
rect 3024 1872 3042 1890
rect 3024 1890 3042 1908
rect 3024 1908 3042 1926
rect 3024 1926 3042 1944
rect 3024 1944 3042 1962
rect 3024 1962 3042 1980
rect 3024 1980 3042 1998
rect 3024 1998 3042 2016
rect 3024 2016 3042 2034
rect 3024 2034 3042 2052
rect 3024 2052 3042 2070
rect 3024 2070 3042 2088
rect 3024 2088 3042 2106
rect 3024 2106 3042 2124
rect 3024 2124 3042 2142
rect 3024 2142 3042 2160
rect 3024 2160 3042 2178
rect 3024 2178 3042 2196
rect 3024 2196 3042 2214
rect 3024 2214 3042 2232
rect 3024 2232 3042 2250
rect 3024 2250 3042 2268
rect 3024 2268 3042 2286
rect 3024 2286 3042 2304
rect 3024 2304 3042 2322
rect 3024 2322 3042 2340
rect 3024 2340 3042 2358
rect 3024 2358 3042 2376
rect 3024 2376 3042 2394
rect 3024 2394 3042 2412
rect 3024 2412 3042 2430
rect 3024 2430 3042 2448
rect 3024 2448 3042 2466
rect 3024 2466 3042 2484
rect 3024 2484 3042 2502
rect 3024 2502 3042 2520
rect 3024 2520 3042 2538
rect 3024 2538 3042 2556
rect 3024 2556 3042 2574
rect 3024 2574 3042 2592
rect 3024 2592 3042 2610
rect 3024 2610 3042 2628
rect 3024 2628 3042 2646
rect 3024 2646 3042 2664
rect 3024 2664 3042 2682
rect 3024 2682 3042 2700
rect 3024 2700 3042 2718
rect 3024 2718 3042 2736
rect 3024 2736 3042 2754
rect 3024 2754 3042 2772
rect 3024 2772 3042 2790
rect 3024 2790 3042 2808
rect 3024 2808 3042 2826
rect 3024 2826 3042 2844
rect 3024 2844 3042 2862
rect 3024 2862 3042 2880
rect 3024 2880 3042 2898
rect 3024 2898 3042 2916
rect 3024 2916 3042 2934
rect 3024 2934 3042 2952
rect 3024 2952 3042 2970
rect 3024 2970 3042 2988
rect 3024 2988 3042 3006
rect 3024 3006 3042 3024
rect 3024 3024 3042 3042
rect 3024 3042 3042 3060
rect 3024 3060 3042 3078
rect 3024 3078 3042 3096
rect 3024 3096 3042 3114
rect 3024 3114 3042 3132
rect 3024 3132 3042 3150
rect 3024 3150 3042 3168
rect 3024 3168 3042 3186
rect 3024 3186 3042 3204
rect 3024 3204 3042 3222
rect 3024 3222 3042 3240
rect 3024 3240 3042 3258
rect 3024 3258 3042 3276
rect 3024 3276 3042 3294
rect 3024 3294 3042 3312
rect 3024 3312 3042 3330
rect 3024 3330 3042 3348
rect 3024 3348 3042 3366
rect 3024 3366 3042 3384
rect 3024 3384 3042 3402
rect 3024 3402 3042 3420
rect 3024 6588 3042 6606
rect 3024 6606 3042 6624
rect 3024 6624 3042 6642
rect 3024 6642 3042 6660
rect 3024 6660 3042 6678
rect 3024 6678 3042 6696
rect 3024 6696 3042 6714
rect 3024 6714 3042 6732
rect 3024 6732 3042 6750
rect 3024 6750 3042 6768
rect 3024 6768 3042 6786
rect 3024 6786 3042 6804
rect 3024 6804 3042 6822
rect 3024 6822 3042 6840
rect 3024 6840 3042 6858
rect 3024 6858 3042 6876
rect 3024 6876 3042 6894
rect 3024 6894 3042 6912
rect 3024 6912 3042 6930
rect 3024 6930 3042 6948
rect 3024 6948 3042 6966
rect 3024 6966 3042 6984
rect 3024 6984 3042 7002
rect 3024 7002 3042 7020
rect 3024 7020 3042 7038
rect 3024 7038 3042 7056
rect 3024 7056 3042 7074
rect 3024 7074 3042 7092
rect 3024 7092 3042 7110
rect 3024 7110 3042 7128
rect 3024 7128 3042 7146
rect 3024 7146 3042 7164
rect 3024 7164 3042 7182
rect 3024 7182 3042 7200
rect 3024 7200 3042 7218
rect 3042 72 3060 90
rect 3042 90 3060 108
rect 3042 108 3060 126
rect 3042 126 3060 144
rect 3042 144 3060 162
rect 3042 162 3060 180
rect 3042 180 3060 198
rect 3042 198 3060 216
rect 3042 216 3060 234
rect 3042 234 3060 252
rect 3042 252 3060 270
rect 3042 270 3060 288
rect 3042 288 3060 306
rect 3042 306 3060 324
rect 3042 324 3060 342
rect 3042 342 3060 360
rect 3042 360 3060 378
rect 3042 378 3060 396
rect 3042 396 3060 414
rect 3042 414 3060 432
rect 3042 594 3060 612
rect 3042 612 3060 630
rect 3042 630 3060 648
rect 3042 648 3060 666
rect 3042 666 3060 684
rect 3042 684 3060 702
rect 3042 702 3060 720
rect 3042 720 3060 738
rect 3042 738 3060 756
rect 3042 756 3060 774
rect 3042 774 3060 792
rect 3042 792 3060 810
rect 3042 810 3060 828
rect 3042 828 3060 846
rect 3042 846 3060 864
rect 3042 864 3060 882
rect 3042 1062 3060 1080
rect 3042 1080 3060 1098
rect 3042 1098 3060 1116
rect 3042 1116 3060 1134
rect 3042 1134 3060 1152
rect 3042 1152 3060 1170
rect 3042 1170 3060 1188
rect 3042 1188 3060 1206
rect 3042 1206 3060 1224
rect 3042 1224 3060 1242
rect 3042 1242 3060 1260
rect 3042 1260 3060 1278
rect 3042 1278 3060 1296
rect 3042 1296 3060 1314
rect 3042 1314 3060 1332
rect 3042 1332 3060 1350
rect 3042 1350 3060 1368
rect 3042 1368 3060 1386
rect 3042 1386 3060 1404
rect 3042 1404 3060 1422
rect 3042 1422 3060 1440
rect 3042 1440 3060 1458
rect 3042 1458 3060 1476
rect 3042 1476 3060 1494
rect 3042 1494 3060 1512
rect 3042 1512 3060 1530
rect 3042 1530 3060 1548
rect 3042 1836 3060 1854
rect 3042 1854 3060 1872
rect 3042 1872 3060 1890
rect 3042 1890 3060 1908
rect 3042 1908 3060 1926
rect 3042 1926 3060 1944
rect 3042 1944 3060 1962
rect 3042 1962 3060 1980
rect 3042 1980 3060 1998
rect 3042 1998 3060 2016
rect 3042 2016 3060 2034
rect 3042 2034 3060 2052
rect 3042 2052 3060 2070
rect 3042 2070 3060 2088
rect 3042 2088 3060 2106
rect 3042 2106 3060 2124
rect 3042 2124 3060 2142
rect 3042 2142 3060 2160
rect 3042 2160 3060 2178
rect 3042 2178 3060 2196
rect 3042 2196 3060 2214
rect 3042 2214 3060 2232
rect 3042 2232 3060 2250
rect 3042 2250 3060 2268
rect 3042 2268 3060 2286
rect 3042 2286 3060 2304
rect 3042 2304 3060 2322
rect 3042 2322 3060 2340
rect 3042 2340 3060 2358
rect 3042 2358 3060 2376
rect 3042 2376 3060 2394
rect 3042 2394 3060 2412
rect 3042 2412 3060 2430
rect 3042 2430 3060 2448
rect 3042 2448 3060 2466
rect 3042 2466 3060 2484
rect 3042 2484 3060 2502
rect 3042 2502 3060 2520
rect 3042 2520 3060 2538
rect 3042 2538 3060 2556
rect 3042 2556 3060 2574
rect 3042 2574 3060 2592
rect 3042 2592 3060 2610
rect 3042 2610 3060 2628
rect 3042 2628 3060 2646
rect 3042 2646 3060 2664
rect 3042 2664 3060 2682
rect 3042 2682 3060 2700
rect 3042 2700 3060 2718
rect 3042 2718 3060 2736
rect 3042 2736 3060 2754
rect 3042 2754 3060 2772
rect 3042 2772 3060 2790
rect 3042 2790 3060 2808
rect 3042 2808 3060 2826
rect 3042 2826 3060 2844
rect 3042 2844 3060 2862
rect 3042 2862 3060 2880
rect 3042 2880 3060 2898
rect 3042 2898 3060 2916
rect 3042 2916 3060 2934
rect 3042 2934 3060 2952
rect 3042 2952 3060 2970
rect 3042 2970 3060 2988
rect 3042 2988 3060 3006
rect 3042 3006 3060 3024
rect 3042 3024 3060 3042
rect 3042 3042 3060 3060
rect 3042 3060 3060 3078
rect 3042 3078 3060 3096
rect 3042 3096 3060 3114
rect 3042 3114 3060 3132
rect 3042 3132 3060 3150
rect 3042 3150 3060 3168
rect 3042 3168 3060 3186
rect 3042 3186 3060 3204
rect 3042 3204 3060 3222
rect 3042 3222 3060 3240
rect 3042 3240 3060 3258
rect 3042 3258 3060 3276
rect 3042 3276 3060 3294
rect 3042 3294 3060 3312
rect 3042 3312 3060 3330
rect 3042 3330 3060 3348
rect 3042 3348 3060 3366
rect 3042 3366 3060 3384
rect 3042 3384 3060 3402
rect 3042 3402 3060 3420
rect 3042 3420 3060 3438
rect 3042 3438 3060 3456
rect 3042 3456 3060 3474
rect 3042 3474 3060 3492
rect 3042 6588 3060 6606
rect 3042 6606 3060 6624
rect 3042 6624 3060 6642
rect 3042 6642 3060 6660
rect 3042 6660 3060 6678
rect 3042 6678 3060 6696
rect 3042 6696 3060 6714
rect 3042 6714 3060 6732
rect 3042 6732 3060 6750
rect 3042 6750 3060 6768
rect 3042 6768 3060 6786
rect 3042 6786 3060 6804
rect 3042 6804 3060 6822
rect 3042 6822 3060 6840
rect 3042 6840 3060 6858
rect 3042 6858 3060 6876
rect 3042 6876 3060 6894
rect 3042 6894 3060 6912
rect 3042 6912 3060 6930
rect 3042 6930 3060 6948
rect 3042 6948 3060 6966
rect 3042 6966 3060 6984
rect 3042 6984 3060 7002
rect 3042 7002 3060 7020
rect 3042 7020 3060 7038
rect 3042 7038 3060 7056
rect 3042 7056 3060 7074
rect 3042 7074 3060 7092
rect 3042 7092 3060 7110
rect 3042 7110 3060 7128
rect 3042 7128 3060 7146
rect 3042 7146 3060 7164
rect 3042 7164 3060 7182
rect 3042 7182 3060 7200
rect 3042 7200 3060 7218
rect 3060 72 3078 90
rect 3060 90 3078 108
rect 3060 108 3078 126
rect 3060 126 3078 144
rect 3060 144 3078 162
rect 3060 162 3078 180
rect 3060 180 3078 198
rect 3060 198 3078 216
rect 3060 216 3078 234
rect 3060 234 3078 252
rect 3060 252 3078 270
rect 3060 270 3078 288
rect 3060 288 3078 306
rect 3060 306 3078 324
rect 3060 324 3078 342
rect 3060 342 3078 360
rect 3060 360 3078 378
rect 3060 378 3078 396
rect 3060 396 3078 414
rect 3060 414 3078 432
rect 3060 432 3078 450
rect 3060 612 3078 630
rect 3060 630 3078 648
rect 3060 648 3078 666
rect 3060 666 3078 684
rect 3060 684 3078 702
rect 3060 702 3078 720
rect 3060 720 3078 738
rect 3060 738 3078 756
rect 3060 756 3078 774
rect 3060 774 3078 792
rect 3060 792 3078 810
rect 3060 810 3078 828
rect 3060 828 3078 846
rect 3060 846 3078 864
rect 3060 864 3078 882
rect 3060 882 3078 900
rect 3060 1080 3078 1098
rect 3060 1098 3078 1116
rect 3060 1116 3078 1134
rect 3060 1134 3078 1152
rect 3060 1152 3078 1170
rect 3060 1170 3078 1188
rect 3060 1188 3078 1206
rect 3060 1206 3078 1224
rect 3060 1224 3078 1242
rect 3060 1242 3078 1260
rect 3060 1260 3078 1278
rect 3060 1278 3078 1296
rect 3060 1296 3078 1314
rect 3060 1314 3078 1332
rect 3060 1332 3078 1350
rect 3060 1350 3078 1368
rect 3060 1368 3078 1386
rect 3060 1386 3078 1404
rect 3060 1404 3078 1422
rect 3060 1422 3078 1440
rect 3060 1440 3078 1458
rect 3060 1458 3078 1476
rect 3060 1476 3078 1494
rect 3060 1494 3078 1512
rect 3060 1512 3078 1530
rect 3060 1530 3078 1548
rect 3060 1548 3078 1566
rect 3060 1566 3078 1584
rect 3060 1872 3078 1890
rect 3060 1890 3078 1908
rect 3060 1908 3078 1926
rect 3060 1926 3078 1944
rect 3060 1944 3078 1962
rect 3060 1962 3078 1980
rect 3060 1980 3078 1998
rect 3060 1998 3078 2016
rect 3060 2016 3078 2034
rect 3060 2034 3078 2052
rect 3060 2052 3078 2070
rect 3060 2070 3078 2088
rect 3060 2088 3078 2106
rect 3060 2106 3078 2124
rect 3060 2124 3078 2142
rect 3060 2142 3078 2160
rect 3060 2160 3078 2178
rect 3060 2178 3078 2196
rect 3060 2196 3078 2214
rect 3060 2214 3078 2232
rect 3060 2232 3078 2250
rect 3060 2250 3078 2268
rect 3060 2268 3078 2286
rect 3060 2286 3078 2304
rect 3060 2304 3078 2322
rect 3060 2322 3078 2340
rect 3060 2340 3078 2358
rect 3060 2358 3078 2376
rect 3060 2376 3078 2394
rect 3060 2394 3078 2412
rect 3060 2412 3078 2430
rect 3060 2430 3078 2448
rect 3060 2448 3078 2466
rect 3060 2466 3078 2484
rect 3060 2484 3078 2502
rect 3060 2502 3078 2520
rect 3060 2520 3078 2538
rect 3060 2538 3078 2556
rect 3060 2556 3078 2574
rect 3060 2574 3078 2592
rect 3060 2592 3078 2610
rect 3060 2610 3078 2628
rect 3060 2628 3078 2646
rect 3060 2646 3078 2664
rect 3060 2664 3078 2682
rect 3060 2682 3078 2700
rect 3060 2700 3078 2718
rect 3060 2718 3078 2736
rect 3060 2736 3078 2754
rect 3060 2754 3078 2772
rect 3060 2772 3078 2790
rect 3060 2790 3078 2808
rect 3060 2808 3078 2826
rect 3060 2826 3078 2844
rect 3060 2844 3078 2862
rect 3060 2862 3078 2880
rect 3060 2880 3078 2898
rect 3060 2898 3078 2916
rect 3060 2916 3078 2934
rect 3060 2934 3078 2952
rect 3060 2952 3078 2970
rect 3060 2970 3078 2988
rect 3060 2988 3078 3006
rect 3060 3006 3078 3024
rect 3060 3024 3078 3042
rect 3060 3042 3078 3060
rect 3060 3060 3078 3078
rect 3060 3078 3078 3096
rect 3060 3096 3078 3114
rect 3060 3114 3078 3132
rect 3060 3132 3078 3150
rect 3060 3150 3078 3168
rect 3060 3168 3078 3186
rect 3060 3186 3078 3204
rect 3060 3204 3078 3222
rect 3060 3222 3078 3240
rect 3060 3240 3078 3258
rect 3060 3258 3078 3276
rect 3060 3276 3078 3294
rect 3060 3294 3078 3312
rect 3060 3312 3078 3330
rect 3060 3330 3078 3348
rect 3060 3348 3078 3366
rect 3060 3366 3078 3384
rect 3060 3384 3078 3402
rect 3060 3402 3078 3420
rect 3060 3420 3078 3438
rect 3060 3438 3078 3456
rect 3060 3456 3078 3474
rect 3060 3474 3078 3492
rect 3060 3492 3078 3510
rect 3060 3510 3078 3528
rect 3060 3528 3078 3546
rect 3060 6588 3078 6606
rect 3060 6606 3078 6624
rect 3060 6624 3078 6642
rect 3060 6642 3078 6660
rect 3060 6660 3078 6678
rect 3060 6678 3078 6696
rect 3060 6696 3078 6714
rect 3060 6714 3078 6732
rect 3060 6732 3078 6750
rect 3060 6750 3078 6768
rect 3060 6768 3078 6786
rect 3060 6786 3078 6804
rect 3060 6804 3078 6822
rect 3060 6822 3078 6840
rect 3060 6840 3078 6858
rect 3060 6858 3078 6876
rect 3060 6876 3078 6894
rect 3060 6894 3078 6912
rect 3060 6912 3078 6930
rect 3060 6930 3078 6948
rect 3060 6948 3078 6966
rect 3060 6966 3078 6984
rect 3060 6984 3078 7002
rect 3060 7002 3078 7020
rect 3060 7020 3078 7038
rect 3060 7038 3078 7056
rect 3060 7056 3078 7074
rect 3060 7074 3078 7092
rect 3060 7092 3078 7110
rect 3060 7110 3078 7128
rect 3060 7128 3078 7146
rect 3060 7146 3078 7164
rect 3060 7164 3078 7182
rect 3060 7182 3078 7200
rect 3060 7200 3078 7218
rect 3060 7218 3078 7236
rect 3078 72 3096 90
rect 3078 90 3096 108
rect 3078 108 3096 126
rect 3078 126 3096 144
rect 3078 144 3096 162
rect 3078 162 3096 180
rect 3078 180 3096 198
rect 3078 198 3096 216
rect 3078 216 3096 234
rect 3078 234 3096 252
rect 3078 252 3096 270
rect 3078 270 3096 288
rect 3078 288 3096 306
rect 3078 306 3096 324
rect 3078 324 3096 342
rect 3078 342 3096 360
rect 3078 360 3096 378
rect 3078 378 3096 396
rect 3078 396 3096 414
rect 3078 414 3096 432
rect 3078 432 3096 450
rect 3078 450 3096 468
rect 3078 612 3096 630
rect 3078 630 3096 648
rect 3078 648 3096 666
rect 3078 666 3096 684
rect 3078 684 3096 702
rect 3078 702 3096 720
rect 3078 720 3096 738
rect 3078 738 3096 756
rect 3078 756 3096 774
rect 3078 774 3096 792
rect 3078 792 3096 810
rect 3078 810 3096 828
rect 3078 828 3096 846
rect 3078 846 3096 864
rect 3078 864 3096 882
rect 3078 882 3096 900
rect 3078 900 3096 918
rect 3078 1098 3096 1116
rect 3078 1116 3096 1134
rect 3078 1134 3096 1152
rect 3078 1152 3096 1170
rect 3078 1170 3096 1188
rect 3078 1188 3096 1206
rect 3078 1206 3096 1224
rect 3078 1224 3096 1242
rect 3078 1242 3096 1260
rect 3078 1260 3096 1278
rect 3078 1278 3096 1296
rect 3078 1296 3096 1314
rect 3078 1314 3096 1332
rect 3078 1332 3096 1350
rect 3078 1350 3096 1368
rect 3078 1368 3096 1386
rect 3078 1386 3096 1404
rect 3078 1404 3096 1422
rect 3078 1422 3096 1440
rect 3078 1440 3096 1458
rect 3078 1458 3096 1476
rect 3078 1476 3096 1494
rect 3078 1494 3096 1512
rect 3078 1512 3096 1530
rect 3078 1530 3096 1548
rect 3078 1548 3096 1566
rect 3078 1566 3096 1584
rect 3078 1584 3096 1602
rect 3078 1602 3096 1620
rect 3078 1908 3096 1926
rect 3078 1926 3096 1944
rect 3078 1944 3096 1962
rect 3078 1962 3096 1980
rect 3078 1980 3096 1998
rect 3078 1998 3096 2016
rect 3078 2016 3096 2034
rect 3078 2034 3096 2052
rect 3078 2052 3096 2070
rect 3078 2070 3096 2088
rect 3078 2088 3096 2106
rect 3078 2106 3096 2124
rect 3078 2124 3096 2142
rect 3078 2142 3096 2160
rect 3078 2160 3096 2178
rect 3078 2178 3096 2196
rect 3078 2196 3096 2214
rect 3078 2214 3096 2232
rect 3078 2232 3096 2250
rect 3078 2250 3096 2268
rect 3078 2268 3096 2286
rect 3078 2286 3096 2304
rect 3078 2304 3096 2322
rect 3078 2322 3096 2340
rect 3078 2340 3096 2358
rect 3078 2358 3096 2376
rect 3078 2376 3096 2394
rect 3078 2394 3096 2412
rect 3078 2412 3096 2430
rect 3078 2430 3096 2448
rect 3078 2448 3096 2466
rect 3078 2466 3096 2484
rect 3078 2484 3096 2502
rect 3078 2502 3096 2520
rect 3078 2520 3096 2538
rect 3078 2538 3096 2556
rect 3078 2556 3096 2574
rect 3078 2574 3096 2592
rect 3078 2592 3096 2610
rect 3078 2610 3096 2628
rect 3078 2628 3096 2646
rect 3078 2646 3096 2664
rect 3078 2664 3096 2682
rect 3078 2682 3096 2700
rect 3078 2700 3096 2718
rect 3078 2718 3096 2736
rect 3078 2736 3096 2754
rect 3078 2754 3096 2772
rect 3078 2772 3096 2790
rect 3078 2790 3096 2808
rect 3078 2808 3096 2826
rect 3078 2826 3096 2844
rect 3078 2844 3096 2862
rect 3078 2862 3096 2880
rect 3078 2880 3096 2898
rect 3078 2898 3096 2916
rect 3078 2916 3096 2934
rect 3078 2934 3096 2952
rect 3078 2952 3096 2970
rect 3078 2970 3096 2988
rect 3078 2988 3096 3006
rect 3078 3006 3096 3024
rect 3078 3024 3096 3042
rect 3078 3042 3096 3060
rect 3078 3060 3096 3078
rect 3078 3078 3096 3096
rect 3078 3096 3096 3114
rect 3078 3114 3096 3132
rect 3078 3132 3096 3150
rect 3078 3150 3096 3168
rect 3078 3168 3096 3186
rect 3078 3186 3096 3204
rect 3078 3204 3096 3222
rect 3078 3222 3096 3240
rect 3078 3240 3096 3258
rect 3078 3258 3096 3276
rect 3078 3276 3096 3294
rect 3078 3294 3096 3312
rect 3078 3312 3096 3330
rect 3078 3330 3096 3348
rect 3078 3348 3096 3366
rect 3078 3366 3096 3384
rect 3078 3384 3096 3402
rect 3078 3402 3096 3420
rect 3078 3420 3096 3438
rect 3078 3438 3096 3456
rect 3078 3456 3096 3474
rect 3078 3474 3096 3492
rect 3078 3492 3096 3510
rect 3078 3510 3096 3528
rect 3078 3528 3096 3546
rect 3078 3546 3096 3564
rect 3078 3564 3096 3582
rect 3078 3582 3096 3600
rect 3078 3600 3096 3618
rect 3078 6588 3096 6606
rect 3078 6606 3096 6624
rect 3078 6624 3096 6642
rect 3078 6642 3096 6660
rect 3078 6660 3096 6678
rect 3078 6678 3096 6696
rect 3078 6696 3096 6714
rect 3078 6714 3096 6732
rect 3078 6732 3096 6750
rect 3078 6750 3096 6768
rect 3078 6768 3096 6786
rect 3078 6786 3096 6804
rect 3078 6804 3096 6822
rect 3078 6822 3096 6840
rect 3078 6840 3096 6858
rect 3078 6858 3096 6876
rect 3078 6876 3096 6894
rect 3078 6894 3096 6912
rect 3078 6912 3096 6930
rect 3078 6930 3096 6948
rect 3078 6948 3096 6966
rect 3078 6966 3096 6984
rect 3078 6984 3096 7002
rect 3078 7002 3096 7020
rect 3078 7020 3096 7038
rect 3078 7038 3096 7056
rect 3078 7056 3096 7074
rect 3078 7074 3096 7092
rect 3078 7092 3096 7110
rect 3078 7110 3096 7128
rect 3078 7128 3096 7146
rect 3078 7146 3096 7164
rect 3078 7164 3096 7182
rect 3078 7182 3096 7200
rect 3078 7200 3096 7218
rect 3078 7218 3096 7236
rect 3096 54 3114 72
rect 3096 72 3114 90
rect 3096 90 3114 108
rect 3096 108 3114 126
rect 3096 126 3114 144
rect 3096 144 3114 162
rect 3096 162 3114 180
rect 3096 180 3114 198
rect 3096 198 3114 216
rect 3096 216 3114 234
rect 3096 234 3114 252
rect 3096 252 3114 270
rect 3096 270 3114 288
rect 3096 288 3114 306
rect 3096 306 3114 324
rect 3096 324 3114 342
rect 3096 342 3114 360
rect 3096 360 3114 378
rect 3096 378 3114 396
rect 3096 396 3114 414
rect 3096 414 3114 432
rect 3096 432 3114 450
rect 3096 450 3114 468
rect 3096 468 3114 486
rect 3096 630 3114 648
rect 3096 648 3114 666
rect 3096 666 3114 684
rect 3096 684 3114 702
rect 3096 702 3114 720
rect 3096 720 3114 738
rect 3096 738 3114 756
rect 3096 756 3114 774
rect 3096 774 3114 792
rect 3096 792 3114 810
rect 3096 810 3114 828
rect 3096 828 3114 846
rect 3096 846 3114 864
rect 3096 864 3114 882
rect 3096 882 3114 900
rect 3096 900 3114 918
rect 3096 918 3114 936
rect 3096 1116 3114 1134
rect 3096 1134 3114 1152
rect 3096 1152 3114 1170
rect 3096 1170 3114 1188
rect 3096 1188 3114 1206
rect 3096 1206 3114 1224
rect 3096 1224 3114 1242
rect 3096 1242 3114 1260
rect 3096 1260 3114 1278
rect 3096 1278 3114 1296
rect 3096 1296 3114 1314
rect 3096 1314 3114 1332
rect 3096 1332 3114 1350
rect 3096 1350 3114 1368
rect 3096 1368 3114 1386
rect 3096 1386 3114 1404
rect 3096 1404 3114 1422
rect 3096 1422 3114 1440
rect 3096 1440 3114 1458
rect 3096 1458 3114 1476
rect 3096 1476 3114 1494
rect 3096 1494 3114 1512
rect 3096 1512 3114 1530
rect 3096 1530 3114 1548
rect 3096 1548 3114 1566
rect 3096 1566 3114 1584
rect 3096 1584 3114 1602
rect 3096 1602 3114 1620
rect 3096 1620 3114 1638
rect 3096 1638 3114 1656
rect 3096 1944 3114 1962
rect 3096 1962 3114 1980
rect 3096 1980 3114 1998
rect 3096 1998 3114 2016
rect 3096 2016 3114 2034
rect 3096 2034 3114 2052
rect 3096 2052 3114 2070
rect 3096 2070 3114 2088
rect 3096 2088 3114 2106
rect 3096 2106 3114 2124
rect 3096 2124 3114 2142
rect 3096 2142 3114 2160
rect 3096 2160 3114 2178
rect 3096 2178 3114 2196
rect 3096 2196 3114 2214
rect 3096 2214 3114 2232
rect 3096 2232 3114 2250
rect 3096 2250 3114 2268
rect 3096 2268 3114 2286
rect 3096 2286 3114 2304
rect 3096 2304 3114 2322
rect 3096 2322 3114 2340
rect 3096 2340 3114 2358
rect 3096 2358 3114 2376
rect 3096 2376 3114 2394
rect 3096 2394 3114 2412
rect 3096 2412 3114 2430
rect 3096 2430 3114 2448
rect 3096 2448 3114 2466
rect 3096 2466 3114 2484
rect 3096 2484 3114 2502
rect 3096 2502 3114 2520
rect 3096 2520 3114 2538
rect 3096 2538 3114 2556
rect 3096 2556 3114 2574
rect 3096 2574 3114 2592
rect 3096 2592 3114 2610
rect 3096 2610 3114 2628
rect 3096 2628 3114 2646
rect 3096 2646 3114 2664
rect 3096 2664 3114 2682
rect 3096 2682 3114 2700
rect 3096 2700 3114 2718
rect 3096 2718 3114 2736
rect 3096 2736 3114 2754
rect 3096 2754 3114 2772
rect 3096 2772 3114 2790
rect 3096 2790 3114 2808
rect 3096 2808 3114 2826
rect 3096 2826 3114 2844
rect 3096 2844 3114 2862
rect 3096 2862 3114 2880
rect 3096 2880 3114 2898
rect 3096 2898 3114 2916
rect 3096 2916 3114 2934
rect 3096 2934 3114 2952
rect 3096 2952 3114 2970
rect 3096 2970 3114 2988
rect 3096 2988 3114 3006
rect 3096 3006 3114 3024
rect 3096 3024 3114 3042
rect 3096 3042 3114 3060
rect 3096 3060 3114 3078
rect 3096 3078 3114 3096
rect 3096 3096 3114 3114
rect 3096 3114 3114 3132
rect 3096 3132 3114 3150
rect 3096 3150 3114 3168
rect 3096 3168 3114 3186
rect 3096 3186 3114 3204
rect 3096 3204 3114 3222
rect 3096 3222 3114 3240
rect 3096 3240 3114 3258
rect 3096 3258 3114 3276
rect 3096 3276 3114 3294
rect 3096 3294 3114 3312
rect 3096 3312 3114 3330
rect 3096 3330 3114 3348
rect 3096 3348 3114 3366
rect 3096 3366 3114 3384
rect 3096 3384 3114 3402
rect 3096 3402 3114 3420
rect 3096 3420 3114 3438
rect 3096 3438 3114 3456
rect 3096 3456 3114 3474
rect 3096 3474 3114 3492
rect 3096 3492 3114 3510
rect 3096 3510 3114 3528
rect 3096 3528 3114 3546
rect 3096 3546 3114 3564
rect 3096 3564 3114 3582
rect 3096 3582 3114 3600
rect 3096 3600 3114 3618
rect 3096 3618 3114 3636
rect 3096 3636 3114 3654
rect 3096 3654 3114 3672
rect 3096 6606 3114 6624
rect 3096 6624 3114 6642
rect 3096 6642 3114 6660
rect 3096 6660 3114 6678
rect 3096 6678 3114 6696
rect 3096 6696 3114 6714
rect 3096 6714 3114 6732
rect 3096 6732 3114 6750
rect 3096 6750 3114 6768
rect 3096 6768 3114 6786
rect 3096 6786 3114 6804
rect 3096 6804 3114 6822
rect 3096 6822 3114 6840
rect 3096 6840 3114 6858
rect 3096 6858 3114 6876
rect 3096 6876 3114 6894
rect 3096 6894 3114 6912
rect 3096 6912 3114 6930
rect 3096 6930 3114 6948
rect 3096 6948 3114 6966
rect 3096 6966 3114 6984
rect 3096 6984 3114 7002
rect 3096 7002 3114 7020
rect 3096 7020 3114 7038
rect 3096 7038 3114 7056
rect 3096 7056 3114 7074
rect 3096 7074 3114 7092
rect 3096 7092 3114 7110
rect 3096 7110 3114 7128
rect 3096 7128 3114 7146
rect 3096 7146 3114 7164
rect 3096 7164 3114 7182
rect 3096 7182 3114 7200
rect 3096 7200 3114 7218
rect 3096 7218 3114 7236
rect 3114 54 3132 72
rect 3114 72 3132 90
rect 3114 90 3132 108
rect 3114 108 3132 126
rect 3114 126 3132 144
rect 3114 144 3132 162
rect 3114 162 3132 180
rect 3114 180 3132 198
rect 3114 198 3132 216
rect 3114 216 3132 234
rect 3114 234 3132 252
rect 3114 252 3132 270
rect 3114 270 3132 288
rect 3114 288 3132 306
rect 3114 306 3132 324
rect 3114 324 3132 342
rect 3114 342 3132 360
rect 3114 360 3132 378
rect 3114 378 3132 396
rect 3114 396 3132 414
rect 3114 414 3132 432
rect 3114 432 3132 450
rect 3114 450 3132 468
rect 3114 468 3132 486
rect 3114 648 3132 666
rect 3114 666 3132 684
rect 3114 684 3132 702
rect 3114 702 3132 720
rect 3114 720 3132 738
rect 3114 738 3132 756
rect 3114 756 3132 774
rect 3114 774 3132 792
rect 3114 792 3132 810
rect 3114 810 3132 828
rect 3114 828 3132 846
rect 3114 846 3132 864
rect 3114 864 3132 882
rect 3114 882 3132 900
rect 3114 900 3132 918
rect 3114 918 3132 936
rect 3114 1134 3132 1152
rect 3114 1152 3132 1170
rect 3114 1170 3132 1188
rect 3114 1188 3132 1206
rect 3114 1206 3132 1224
rect 3114 1224 3132 1242
rect 3114 1242 3132 1260
rect 3114 1260 3132 1278
rect 3114 1278 3132 1296
rect 3114 1296 3132 1314
rect 3114 1314 3132 1332
rect 3114 1332 3132 1350
rect 3114 1350 3132 1368
rect 3114 1368 3132 1386
rect 3114 1386 3132 1404
rect 3114 1404 3132 1422
rect 3114 1422 3132 1440
rect 3114 1440 3132 1458
rect 3114 1458 3132 1476
rect 3114 1476 3132 1494
rect 3114 1494 3132 1512
rect 3114 1512 3132 1530
rect 3114 1530 3132 1548
rect 3114 1548 3132 1566
rect 3114 1566 3132 1584
rect 3114 1584 3132 1602
rect 3114 1602 3132 1620
rect 3114 1620 3132 1638
rect 3114 1638 3132 1656
rect 3114 1656 3132 1674
rect 3114 1674 3132 1692
rect 3114 1962 3132 1980
rect 3114 1980 3132 1998
rect 3114 1998 3132 2016
rect 3114 2016 3132 2034
rect 3114 2034 3132 2052
rect 3114 2052 3132 2070
rect 3114 2070 3132 2088
rect 3114 2088 3132 2106
rect 3114 2106 3132 2124
rect 3114 2124 3132 2142
rect 3114 2142 3132 2160
rect 3114 2160 3132 2178
rect 3114 2178 3132 2196
rect 3114 2196 3132 2214
rect 3114 2214 3132 2232
rect 3114 2232 3132 2250
rect 3114 2250 3132 2268
rect 3114 2268 3132 2286
rect 3114 2286 3132 2304
rect 3114 2304 3132 2322
rect 3114 2322 3132 2340
rect 3114 2340 3132 2358
rect 3114 2358 3132 2376
rect 3114 2376 3132 2394
rect 3114 2394 3132 2412
rect 3114 2412 3132 2430
rect 3114 2430 3132 2448
rect 3114 2448 3132 2466
rect 3114 2466 3132 2484
rect 3114 2484 3132 2502
rect 3114 2502 3132 2520
rect 3114 2520 3132 2538
rect 3114 2538 3132 2556
rect 3114 2556 3132 2574
rect 3114 2574 3132 2592
rect 3114 2592 3132 2610
rect 3114 2610 3132 2628
rect 3114 2628 3132 2646
rect 3114 2646 3132 2664
rect 3114 2664 3132 2682
rect 3114 2682 3132 2700
rect 3114 2700 3132 2718
rect 3114 2718 3132 2736
rect 3114 2736 3132 2754
rect 3114 2754 3132 2772
rect 3114 2772 3132 2790
rect 3114 2790 3132 2808
rect 3114 2808 3132 2826
rect 3114 2826 3132 2844
rect 3114 2844 3132 2862
rect 3114 2862 3132 2880
rect 3114 2880 3132 2898
rect 3114 2898 3132 2916
rect 3114 2916 3132 2934
rect 3114 2934 3132 2952
rect 3114 2952 3132 2970
rect 3114 2970 3132 2988
rect 3114 2988 3132 3006
rect 3114 3006 3132 3024
rect 3114 3024 3132 3042
rect 3114 3042 3132 3060
rect 3114 3060 3132 3078
rect 3114 3078 3132 3096
rect 3114 3096 3132 3114
rect 3114 3114 3132 3132
rect 3114 3132 3132 3150
rect 3114 3150 3132 3168
rect 3114 3168 3132 3186
rect 3114 3186 3132 3204
rect 3114 3204 3132 3222
rect 3114 3222 3132 3240
rect 3114 3240 3132 3258
rect 3114 3258 3132 3276
rect 3114 3276 3132 3294
rect 3114 3294 3132 3312
rect 3114 3312 3132 3330
rect 3114 3330 3132 3348
rect 3114 3348 3132 3366
rect 3114 3366 3132 3384
rect 3114 3384 3132 3402
rect 3114 3402 3132 3420
rect 3114 3420 3132 3438
rect 3114 3438 3132 3456
rect 3114 3456 3132 3474
rect 3114 3474 3132 3492
rect 3114 3492 3132 3510
rect 3114 3510 3132 3528
rect 3114 3528 3132 3546
rect 3114 3546 3132 3564
rect 3114 3564 3132 3582
rect 3114 3582 3132 3600
rect 3114 3600 3132 3618
rect 3114 3618 3132 3636
rect 3114 3636 3132 3654
rect 3114 3654 3132 3672
rect 3114 3672 3132 3690
rect 3114 3690 3132 3708
rect 3114 3708 3132 3726
rect 3114 6606 3132 6624
rect 3114 6624 3132 6642
rect 3114 6642 3132 6660
rect 3114 6660 3132 6678
rect 3114 6678 3132 6696
rect 3114 6696 3132 6714
rect 3114 6714 3132 6732
rect 3114 6732 3132 6750
rect 3114 6750 3132 6768
rect 3114 6768 3132 6786
rect 3114 6786 3132 6804
rect 3114 6804 3132 6822
rect 3114 6822 3132 6840
rect 3114 6840 3132 6858
rect 3114 6858 3132 6876
rect 3114 6876 3132 6894
rect 3114 6894 3132 6912
rect 3114 6912 3132 6930
rect 3114 6930 3132 6948
rect 3114 6948 3132 6966
rect 3114 6966 3132 6984
rect 3114 6984 3132 7002
rect 3114 7002 3132 7020
rect 3114 7020 3132 7038
rect 3114 7038 3132 7056
rect 3114 7056 3132 7074
rect 3114 7074 3132 7092
rect 3114 7092 3132 7110
rect 3114 7110 3132 7128
rect 3114 7128 3132 7146
rect 3114 7146 3132 7164
rect 3114 7164 3132 7182
rect 3114 7182 3132 7200
rect 3114 7200 3132 7218
rect 3114 7218 3132 7236
rect 3132 54 3150 72
rect 3132 72 3150 90
rect 3132 90 3150 108
rect 3132 108 3150 126
rect 3132 126 3150 144
rect 3132 144 3150 162
rect 3132 162 3150 180
rect 3132 180 3150 198
rect 3132 198 3150 216
rect 3132 216 3150 234
rect 3132 234 3150 252
rect 3132 252 3150 270
rect 3132 270 3150 288
rect 3132 288 3150 306
rect 3132 306 3150 324
rect 3132 324 3150 342
rect 3132 342 3150 360
rect 3132 360 3150 378
rect 3132 378 3150 396
rect 3132 396 3150 414
rect 3132 414 3150 432
rect 3132 432 3150 450
rect 3132 450 3150 468
rect 3132 468 3150 486
rect 3132 486 3150 504
rect 3132 648 3150 666
rect 3132 666 3150 684
rect 3132 684 3150 702
rect 3132 702 3150 720
rect 3132 720 3150 738
rect 3132 738 3150 756
rect 3132 756 3150 774
rect 3132 774 3150 792
rect 3132 792 3150 810
rect 3132 810 3150 828
rect 3132 828 3150 846
rect 3132 846 3150 864
rect 3132 864 3150 882
rect 3132 882 3150 900
rect 3132 900 3150 918
rect 3132 918 3150 936
rect 3132 936 3150 954
rect 3132 1134 3150 1152
rect 3132 1152 3150 1170
rect 3132 1170 3150 1188
rect 3132 1188 3150 1206
rect 3132 1206 3150 1224
rect 3132 1224 3150 1242
rect 3132 1242 3150 1260
rect 3132 1260 3150 1278
rect 3132 1278 3150 1296
rect 3132 1296 3150 1314
rect 3132 1314 3150 1332
rect 3132 1332 3150 1350
rect 3132 1350 3150 1368
rect 3132 1368 3150 1386
rect 3132 1386 3150 1404
rect 3132 1404 3150 1422
rect 3132 1422 3150 1440
rect 3132 1440 3150 1458
rect 3132 1458 3150 1476
rect 3132 1476 3150 1494
rect 3132 1494 3150 1512
rect 3132 1512 3150 1530
rect 3132 1530 3150 1548
rect 3132 1548 3150 1566
rect 3132 1566 3150 1584
rect 3132 1584 3150 1602
rect 3132 1602 3150 1620
rect 3132 1620 3150 1638
rect 3132 1638 3150 1656
rect 3132 1656 3150 1674
rect 3132 1674 3150 1692
rect 3132 1692 3150 1710
rect 3132 1710 3150 1728
rect 3132 1998 3150 2016
rect 3132 2016 3150 2034
rect 3132 2034 3150 2052
rect 3132 2052 3150 2070
rect 3132 2070 3150 2088
rect 3132 2088 3150 2106
rect 3132 2106 3150 2124
rect 3132 2124 3150 2142
rect 3132 2142 3150 2160
rect 3132 2160 3150 2178
rect 3132 2178 3150 2196
rect 3132 2196 3150 2214
rect 3132 2214 3150 2232
rect 3132 2232 3150 2250
rect 3132 2250 3150 2268
rect 3132 2268 3150 2286
rect 3132 2286 3150 2304
rect 3132 2304 3150 2322
rect 3132 2322 3150 2340
rect 3132 2340 3150 2358
rect 3132 2358 3150 2376
rect 3132 2376 3150 2394
rect 3132 2394 3150 2412
rect 3132 2412 3150 2430
rect 3132 2430 3150 2448
rect 3132 2448 3150 2466
rect 3132 2466 3150 2484
rect 3132 2484 3150 2502
rect 3132 2502 3150 2520
rect 3132 2520 3150 2538
rect 3132 2538 3150 2556
rect 3132 2556 3150 2574
rect 3132 2574 3150 2592
rect 3132 2592 3150 2610
rect 3132 2610 3150 2628
rect 3132 2628 3150 2646
rect 3132 2646 3150 2664
rect 3132 2664 3150 2682
rect 3132 2682 3150 2700
rect 3132 2700 3150 2718
rect 3132 2718 3150 2736
rect 3132 2736 3150 2754
rect 3132 2754 3150 2772
rect 3132 2772 3150 2790
rect 3132 2790 3150 2808
rect 3132 2808 3150 2826
rect 3132 2826 3150 2844
rect 3132 2844 3150 2862
rect 3132 2862 3150 2880
rect 3132 2880 3150 2898
rect 3132 2898 3150 2916
rect 3132 2916 3150 2934
rect 3132 2934 3150 2952
rect 3132 2952 3150 2970
rect 3132 2970 3150 2988
rect 3132 2988 3150 3006
rect 3132 3006 3150 3024
rect 3132 3024 3150 3042
rect 3132 3042 3150 3060
rect 3132 3060 3150 3078
rect 3132 3078 3150 3096
rect 3132 3096 3150 3114
rect 3132 3114 3150 3132
rect 3132 3132 3150 3150
rect 3132 3150 3150 3168
rect 3132 3168 3150 3186
rect 3132 3186 3150 3204
rect 3132 3204 3150 3222
rect 3132 3222 3150 3240
rect 3132 3240 3150 3258
rect 3132 3258 3150 3276
rect 3132 3276 3150 3294
rect 3132 3294 3150 3312
rect 3132 3312 3150 3330
rect 3132 3330 3150 3348
rect 3132 3348 3150 3366
rect 3132 3366 3150 3384
rect 3132 3384 3150 3402
rect 3132 3402 3150 3420
rect 3132 3420 3150 3438
rect 3132 3438 3150 3456
rect 3132 3456 3150 3474
rect 3132 3474 3150 3492
rect 3132 3492 3150 3510
rect 3132 3510 3150 3528
rect 3132 3528 3150 3546
rect 3132 3546 3150 3564
rect 3132 3564 3150 3582
rect 3132 3582 3150 3600
rect 3132 3600 3150 3618
rect 3132 3618 3150 3636
rect 3132 3636 3150 3654
rect 3132 3654 3150 3672
rect 3132 3672 3150 3690
rect 3132 3690 3150 3708
rect 3132 3708 3150 3726
rect 3132 3726 3150 3744
rect 3132 3744 3150 3762
rect 3132 3762 3150 3780
rect 3132 3780 3150 3798
rect 3132 6606 3150 6624
rect 3132 6624 3150 6642
rect 3132 6642 3150 6660
rect 3132 6660 3150 6678
rect 3132 6678 3150 6696
rect 3132 6696 3150 6714
rect 3132 6714 3150 6732
rect 3132 6732 3150 6750
rect 3132 6750 3150 6768
rect 3132 6768 3150 6786
rect 3132 6786 3150 6804
rect 3132 6804 3150 6822
rect 3132 6822 3150 6840
rect 3132 6840 3150 6858
rect 3132 6858 3150 6876
rect 3132 6876 3150 6894
rect 3132 6894 3150 6912
rect 3132 6912 3150 6930
rect 3132 6930 3150 6948
rect 3132 6948 3150 6966
rect 3132 6966 3150 6984
rect 3132 6984 3150 7002
rect 3132 7002 3150 7020
rect 3132 7020 3150 7038
rect 3132 7038 3150 7056
rect 3132 7056 3150 7074
rect 3132 7074 3150 7092
rect 3132 7092 3150 7110
rect 3132 7110 3150 7128
rect 3132 7128 3150 7146
rect 3132 7146 3150 7164
rect 3132 7164 3150 7182
rect 3132 7182 3150 7200
rect 3132 7200 3150 7218
rect 3132 7218 3150 7236
rect 3150 54 3168 72
rect 3150 72 3168 90
rect 3150 90 3168 108
rect 3150 108 3168 126
rect 3150 126 3168 144
rect 3150 144 3168 162
rect 3150 162 3168 180
rect 3150 180 3168 198
rect 3150 198 3168 216
rect 3150 216 3168 234
rect 3150 234 3168 252
rect 3150 252 3168 270
rect 3150 270 3168 288
rect 3150 288 3168 306
rect 3150 306 3168 324
rect 3150 324 3168 342
rect 3150 342 3168 360
rect 3150 360 3168 378
rect 3150 378 3168 396
rect 3150 396 3168 414
rect 3150 414 3168 432
rect 3150 432 3168 450
rect 3150 450 3168 468
rect 3150 468 3168 486
rect 3150 486 3168 504
rect 3150 504 3168 522
rect 3150 666 3168 684
rect 3150 684 3168 702
rect 3150 702 3168 720
rect 3150 720 3168 738
rect 3150 738 3168 756
rect 3150 756 3168 774
rect 3150 774 3168 792
rect 3150 792 3168 810
rect 3150 810 3168 828
rect 3150 828 3168 846
rect 3150 846 3168 864
rect 3150 864 3168 882
rect 3150 882 3168 900
rect 3150 900 3168 918
rect 3150 918 3168 936
rect 3150 936 3168 954
rect 3150 954 3168 972
rect 3150 1152 3168 1170
rect 3150 1170 3168 1188
rect 3150 1188 3168 1206
rect 3150 1206 3168 1224
rect 3150 1224 3168 1242
rect 3150 1242 3168 1260
rect 3150 1260 3168 1278
rect 3150 1278 3168 1296
rect 3150 1296 3168 1314
rect 3150 1314 3168 1332
rect 3150 1332 3168 1350
rect 3150 1350 3168 1368
rect 3150 1368 3168 1386
rect 3150 1386 3168 1404
rect 3150 1404 3168 1422
rect 3150 1422 3168 1440
rect 3150 1440 3168 1458
rect 3150 1458 3168 1476
rect 3150 1476 3168 1494
rect 3150 1494 3168 1512
rect 3150 1512 3168 1530
rect 3150 1530 3168 1548
rect 3150 1548 3168 1566
rect 3150 1566 3168 1584
rect 3150 1584 3168 1602
rect 3150 1602 3168 1620
rect 3150 1620 3168 1638
rect 3150 1638 3168 1656
rect 3150 1656 3168 1674
rect 3150 1674 3168 1692
rect 3150 1692 3168 1710
rect 3150 1710 3168 1728
rect 3150 1728 3168 1746
rect 3150 2034 3168 2052
rect 3150 2052 3168 2070
rect 3150 2070 3168 2088
rect 3150 2088 3168 2106
rect 3150 2106 3168 2124
rect 3150 2124 3168 2142
rect 3150 2142 3168 2160
rect 3150 2160 3168 2178
rect 3150 2178 3168 2196
rect 3150 2196 3168 2214
rect 3150 2214 3168 2232
rect 3150 2232 3168 2250
rect 3150 2250 3168 2268
rect 3150 2268 3168 2286
rect 3150 2286 3168 2304
rect 3150 2304 3168 2322
rect 3150 2322 3168 2340
rect 3150 2340 3168 2358
rect 3150 2358 3168 2376
rect 3150 2376 3168 2394
rect 3150 2394 3168 2412
rect 3150 2412 3168 2430
rect 3150 2430 3168 2448
rect 3150 2448 3168 2466
rect 3150 2466 3168 2484
rect 3150 2484 3168 2502
rect 3150 2502 3168 2520
rect 3150 2520 3168 2538
rect 3150 2538 3168 2556
rect 3150 2556 3168 2574
rect 3150 2574 3168 2592
rect 3150 2592 3168 2610
rect 3150 2610 3168 2628
rect 3150 2628 3168 2646
rect 3150 2646 3168 2664
rect 3150 2664 3168 2682
rect 3150 2682 3168 2700
rect 3150 2700 3168 2718
rect 3150 2718 3168 2736
rect 3150 2736 3168 2754
rect 3150 2754 3168 2772
rect 3150 2772 3168 2790
rect 3150 2790 3168 2808
rect 3150 2808 3168 2826
rect 3150 2826 3168 2844
rect 3150 2844 3168 2862
rect 3150 2862 3168 2880
rect 3150 2880 3168 2898
rect 3150 2898 3168 2916
rect 3150 2916 3168 2934
rect 3150 2934 3168 2952
rect 3150 2952 3168 2970
rect 3150 2970 3168 2988
rect 3150 2988 3168 3006
rect 3150 3006 3168 3024
rect 3150 3024 3168 3042
rect 3150 3042 3168 3060
rect 3150 3060 3168 3078
rect 3150 3078 3168 3096
rect 3150 3096 3168 3114
rect 3150 3114 3168 3132
rect 3150 3132 3168 3150
rect 3150 3150 3168 3168
rect 3150 3168 3168 3186
rect 3150 3186 3168 3204
rect 3150 3204 3168 3222
rect 3150 3222 3168 3240
rect 3150 3240 3168 3258
rect 3150 3258 3168 3276
rect 3150 3276 3168 3294
rect 3150 3294 3168 3312
rect 3150 3312 3168 3330
rect 3150 3330 3168 3348
rect 3150 3348 3168 3366
rect 3150 3366 3168 3384
rect 3150 3384 3168 3402
rect 3150 3402 3168 3420
rect 3150 3420 3168 3438
rect 3150 3438 3168 3456
rect 3150 3456 3168 3474
rect 3150 3474 3168 3492
rect 3150 3492 3168 3510
rect 3150 3510 3168 3528
rect 3150 3528 3168 3546
rect 3150 3546 3168 3564
rect 3150 3564 3168 3582
rect 3150 3582 3168 3600
rect 3150 3600 3168 3618
rect 3150 3618 3168 3636
rect 3150 3636 3168 3654
rect 3150 3654 3168 3672
rect 3150 3672 3168 3690
rect 3150 3690 3168 3708
rect 3150 3708 3168 3726
rect 3150 3726 3168 3744
rect 3150 3744 3168 3762
rect 3150 3762 3168 3780
rect 3150 3780 3168 3798
rect 3150 3798 3168 3816
rect 3150 3816 3168 3834
rect 3150 3834 3168 3852
rect 3150 6606 3168 6624
rect 3150 6624 3168 6642
rect 3150 6642 3168 6660
rect 3150 6660 3168 6678
rect 3150 6678 3168 6696
rect 3150 6696 3168 6714
rect 3150 6714 3168 6732
rect 3150 6732 3168 6750
rect 3150 6750 3168 6768
rect 3150 6768 3168 6786
rect 3150 6786 3168 6804
rect 3150 6804 3168 6822
rect 3150 6822 3168 6840
rect 3150 6840 3168 6858
rect 3150 6858 3168 6876
rect 3150 6876 3168 6894
rect 3150 6894 3168 6912
rect 3150 6912 3168 6930
rect 3150 6930 3168 6948
rect 3150 6948 3168 6966
rect 3150 6966 3168 6984
rect 3150 6984 3168 7002
rect 3150 7002 3168 7020
rect 3150 7020 3168 7038
rect 3150 7038 3168 7056
rect 3150 7056 3168 7074
rect 3150 7074 3168 7092
rect 3150 7092 3168 7110
rect 3150 7110 3168 7128
rect 3150 7128 3168 7146
rect 3150 7146 3168 7164
rect 3150 7164 3168 7182
rect 3150 7182 3168 7200
rect 3150 7200 3168 7218
rect 3150 7218 3168 7236
rect 3168 54 3186 72
rect 3168 72 3186 90
rect 3168 90 3186 108
rect 3168 108 3186 126
rect 3168 126 3186 144
rect 3168 144 3186 162
rect 3168 162 3186 180
rect 3168 180 3186 198
rect 3168 198 3186 216
rect 3168 216 3186 234
rect 3168 234 3186 252
rect 3168 252 3186 270
rect 3168 270 3186 288
rect 3168 288 3186 306
rect 3168 306 3186 324
rect 3168 324 3186 342
rect 3168 342 3186 360
rect 3168 360 3186 378
rect 3168 378 3186 396
rect 3168 396 3186 414
rect 3168 414 3186 432
rect 3168 432 3186 450
rect 3168 450 3186 468
rect 3168 468 3186 486
rect 3168 486 3186 504
rect 3168 504 3186 522
rect 3168 522 3186 540
rect 3168 666 3186 684
rect 3168 684 3186 702
rect 3168 702 3186 720
rect 3168 720 3186 738
rect 3168 738 3186 756
rect 3168 756 3186 774
rect 3168 774 3186 792
rect 3168 792 3186 810
rect 3168 810 3186 828
rect 3168 828 3186 846
rect 3168 846 3186 864
rect 3168 864 3186 882
rect 3168 882 3186 900
rect 3168 900 3186 918
rect 3168 918 3186 936
rect 3168 936 3186 954
rect 3168 954 3186 972
rect 3168 972 3186 990
rect 3168 1170 3186 1188
rect 3168 1188 3186 1206
rect 3168 1206 3186 1224
rect 3168 1224 3186 1242
rect 3168 1242 3186 1260
rect 3168 1260 3186 1278
rect 3168 1278 3186 1296
rect 3168 1296 3186 1314
rect 3168 1314 3186 1332
rect 3168 1332 3186 1350
rect 3168 1350 3186 1368
rect 3168 1368 3186 1386
rect 3168 1386 3186 1404
rect 3168 1404 3186 1422
rect 3168 1422 3186 1440
rect 3168 1440 3186 1458
rect 3168 1458 3186 1476
rect 3168 1476 3186 1494
rect 3168 1494 3186 1512
rect 3168 1512 3186 1530
rect 3168 1530 3186 1548
rect 3168 1548 3186 1566
rect 3168 1566 3186 1584
rect 3168 1584 3186 1602
rect 3168 1602 3186 1620
rect 3168 1620 3186 1638
rect 3168 1638 3186 1656
rect 3168 1656 3186 1674
rect 3168 1674 3186 1692
rect 3168 1692 3186 1710
rect 3168 1710 3186 1728
rect 3168 1728 3186 1746
rect 3168 1746 3186 1764
rect 3168 1764 3186 1782
rect 3168 2070 3186 2088
rect 3168 2088 3186 2106
rect 3168 2106 3186 2124
rect 3168 2124 3186 2142
rect 3168 2142 3186 2160
rect 3168 2160 3186 2178
rect 3168 2178 3186 2196
rect 3168 2196 3186 2214
rect 3168 2214 3186 2232
rect 3168 2232 3186 2250
rect 3168 2250 3186 2268
rect 3168 2268 3186 2286
rect 3168 2286 3186 2304
rect 3168 2304 3186 2322
rect 3168 2322 3186 2340
rect 3168 2340 3186 2358
rect 3168 2358 3186 2376
rect 3168 2376 3186 2394
rect 3168 2394 3186 2412
rect 3168 2412 3186 2430
rect 3168 2430 3186 2448
rect 3168 2448 3186 2466
rect 3168 2466 3186 2484
rect 3168 2484 3186 2502
rect 3168 2502 3186 2520
rect 3168 2520 3186 2538
rect 3168 2538 3186 2556
rect 3168 2556 3186 2574
rect 3168 2574 3186 2592
rect 3168 2592 3186 2610
rect 3168 2610 3186 2628
rect 3168 2628 3186 2646
rect 3168 2646 3186 2664
rect 3168 2664 3186 2682
rect 3168 2682 3186 2700
rect 3168 2700 3186 2718
rect 3168 2718 3186 2736
rect 3168 2736 3186 2754
rect 3168 2754 3186 2772
rect 3168 2772 3186 2790
rect 3168 2790 3186 2808
rect 3168 2808 3186 2826
rect 3168 2826 3186 2844
rect 3168 2844 3186 2862
rect 3168 2862 3186 2880
rect 3168 2880 3186 2898
rect 3168 2898 3186 2916
rect 3168 2916 3186 2934
rect 3168 2934 3186 2952
rect 3168 2952 3186 2970
rect 3168 2970 3186 2988
rect 3168 2988 3186 3006
rect 3168 3006 3186 3024
rect 3168 3024 3186 3042
rect 3168 3042 3186 3060
rect 3168 3060 3186 3078
rect 3168 3078 3186 3096
rect 3168 3096 3186 3114
rect 3168 3114 3186 3132
rect 3168 3132 3186 3150
rect 3168 3150 3186 3168
rect 3168 3168 3186 3186
rect 3168 3186 3186 3204
rect 3168 3204 3186 3222
rect 3168 3222 3186 3240
rect 3168 3240 3186 3258
rect 3168 3258 3186 3276
rect 3168 3276 3186 3294
rect 3168 3294 3186 3312
rect 3168 3312 3186 3330
rect 3168 3330 3186 3348
rect 3168 3348 3186 3366
rect 3168 3366 3186 3384
rect 3168 3384 3186 3402
rect 3168 3402 3186 3420
rect 3168 3420 3186 3438
rect 3168 3438 3186 3456
rect 3168 3456 3186 3474
rect 3168 3474 3186 3492
rect 3168 3492 3186 3510
rect 3168 3510 3186 3528
rect 3168 3528 3186 3546
rect 3168 3546 3186 3564
rect 3168 3564 3186 3582
rect 3168 3582 3186 3600
rect 3168 3600 3186 3618
rect 3168 3618 3186 3636
rect 3168 3636 3186 3654
rect 3168 3654 3186 3672
rect 3168 3672 3186 3690
rect 3168 3690 3186 3708
rect 3168 3708 3186 3726
rect 3168 3726 3186 3744
rect 3168 3744 3186 3762
rect 3168 3762 3186 3780
rect 3168 3780 3186 3798
rect 3168 3798 3186 3816
rect 3168 3816 3186 3834
rect 3168 3834 3186 3852
rect 3168 3852 3186 3870
rect 3168 3870 3186 3888
rect 3168 3888 3186 3906
rect 3168 6606 3186 6624
rect 3168 6624 3186 6642
rect 3168 6642 3186 6660
rect 3168 6660 3186 6678
rect 3168 6678 3186 6696
rect 3168 6696 3186 6714
rect 3168 6714 3186 6732
rect 3168 6732 3186 6750
rect 3168 6750 3186 6768
rect 3168 6768 3186 6786
rect 3168 6786 3186 6804
rect 3168 6804 3186 6822
rect 3168 6822 3186 6840
rect 3168 6840 3186 6858
rect 3168 6858 3186 6876
rect 3168 6876 3186 6894
rect 3168 6894 3186 6912
rect 3168 6912 3186 6930
rect 3168 6930 3186 6948
rect 3168 6948 3186 6966
rect 3168 6966 3186 6984
rect 3168 6984 3186 7002
rect 3168 7002 3186 7020
rect 3168 7020 3186 7038
rect 3168 7038 3186 7056
rect 3168 7056 3186 7074
rect 3168 7074 3186 7092
rect 3168 7092 3186 7110
rect 3168 7110 3186 7128
rect 3168 7128 3186 7146
rect 3168 7146 3186 7164
rect 3168 7164 3186 7182
rect 3168 7182 3186 7200
rect 3168 7200 3186 7218
rect 3168 7218 3186 7236
rect 3186 54 3204 72
rect 3186 72 3204 90
rect 3186 90 3204 108
rect 3186 108 3204 126
rect 3186 126 3204 144
rect 3186 144 3204 162
rect 3186 162 3204 180
rect 3186 180 3204 198
rect 3186 198 3204 216
rect 3186 216 3204 234
rect 3186 234 3204 252
rect 3186 252 3204 270
rect 3186 270 3204 288
rect 3186 288 3204 306
rect 3186 306 3204 324
rect 3186 324 3204 342
rect 3186 342 3204 360
rect 3186 360 3204 378
rect 3186 378 3204 396
rect 3186 396 3204 414
rect 3186 414 3204 432
rect 3186 432 3204 450
rect 3186 450 3204 468
rect 3186 468 3204 486
rect 3186 486 3204 504
rect 3186 504 3204 522
rect 3186 522 3204 540
rect 3186 540 3204 558
rect 3186 684 3204 702
rect 3186 702 3204 720
rect 3186 720 3204 738
rect 3186 738 3204 756
rect 3186 756 3204 774
rect 3186 774 3204 792
rect 3186 792 3204 810
rect 3186 810 3204 828
rect 3186 828 3204 846
rect 3186 846 3204 864
rect 3186 864 3204 882
rect 3186 882 3204 900
rect 3186 900 3204 918
rect 3186 918 3204 936
rect 3186 936 3204 954
rect 3186 954 3204 972
rect 3186 972 3204 990
rect 3186 1188 3204 1206
rect 3186 1206 3204 1224
rect 3186 1224 3204 1242
rect 3186 1242 3204 1260
rect 3186 1260 3204 1278
rect 3186 1278 3204 1296
rect 3186 1296 3204 1314
rect 3186 1314 3204 1332
rect 3186 1332 3204 1350
rect 3186 1350 3204 1368
rect 3186 1368 3204 1386
rect 3186 1386 3204 1404
rect 3186 1404 3204 1422
rect 3186 1422 3204 1440
rect 3186 1440 3204 1458
rect 3186 1458 3204 1476
rect 3186 1476 3204 1494
rect 3186 1494 3204 1512
rect 3186 1512 3204 1530
rect 3186 1530 3204 1548
rect 3186 1548 3204 1566
rect 3186 1566 3204 1584
rect 3186 1584 3204 1602
rect 3186 1602 3204 1620
rect 3186 1620 3204 1638
rect 3186 1638 3204 1656
rect 3186 1656 3204 1674
rect 3186 1674 3204 1692
rect 3186 1692 3204 1710
rect 3186 1710 3204 1728
rect 3186 1728 3204 1746
rect 3186 1746 3204 1764
rect 3186 1764 3204 1782
rect 3186 1782 3204 1800
rect 3186 1800 3204 1818
rect 3186 2088 3204 2106
rect 3186 2106 3204 2124
rect 3186 2124 3204 2142
rect 3186 2142 3204 2160
rect 3186 2160 3204 2178
rect 3186 2178 3204 2196
rect 3186 2196 3204 2214
rect 3186 2214 3204 2232
rect 3186 2232 3204 2250
rect 3186 2250 3204 2268
rect 3186 2268 3204 2286
rect 3186 2286 3204 2304
rect 3186 2304 3204 2322
rect 3186 2322 3204 2340
rect 3186 2340 3204 2358
rect 3186 2358 3204 2376
rect 3186 2376 3204 2394
rect 3186 2394 3204 2412
rect 3186 2412 3204 2430
rect 3186 2430 3204 2448
rect 3186 2448 3204 2466
rect 3186 2466 3204 2484
rect 3186 2484 3204 2502
rect 3186 2502 3204 2520
rect 3186 2520 3204 2538
rect 3186 2538 3204 2556
rect 3186 2556 3204 2574
rect 3186 2574 3204 2592
rect 3186 2592 3204 2610
rect 3186 2610 3204 2628
rect 3186 2628 3204 2646
rect 3186 2646 3204 2664
rect 3186 2664 3204 2682
rect 3186 2682 3204 2700
rect 3186 2700 3204 2718
rect 3186 2718 3204 2736
rect 3186 2736 3204 2754
rect 3186 2754 3204 2772
rect 3186 2772 3204 2790
rect 3186 2790 3204 2808
rect 3186 2808 3204 2826
rect 3186 2826 3204 2844
rect 3186 2844 3204 2862
rect 3186 2862 3204 2880
rect 3186 2880 3204 2898
rect 3186 2898 3204 2916
rect 3186 2916 3204 2934
rect 3186 2934 3204 2952
rect 3186 2952 3204 2970
rect 3186 2970 3204 2988
rect 3186 2988 3204 3006
rect 3186 3006 3204 3024
rect 3186 3024 3204 3042
rect 3186 3042 3204 3060
rect 3186 3060 3204 3078
rect 3186 3078 3204 3096
rect 3186 3096 3204 3114
rect 3186 3114 3204 3132
rect 3186 3132 3204 3150
rect 3186 3150 3204 3168
rect 3186 3168 3204 3186
rect 3186 3186 3204 3204
rect 3186 3204 3204 3222
rect 3186 3222 3204 3240
rect 3186 3240 3204 3258
rect 3186 3258 3204 3276
rect 3186 3276 3204 3294
rect 3186 3294 3204 3312
rect 3186 3312 3204 3330
rect 3186 3330 3204 3348
rect 3186 3348 3204 3366
rect 3186 3366 3204 3384
rect 3186 3384 3204 3402
rect 3186 3402 3204 3420
rect 3186 3420 3204 3438
rect 3186 3438 3204 3456
rect 3186 3456 3204 3474
rect 3186 3474 3204 3492
rect 3186 3492 3204 3510
rect 3186 3510 3204 3528
rect 3186 3528 3204 3546
rect 3186 3546 3204 3564
rect 3186 3564 3204 3582
rect 3186 3582 3204 3600
rect 3186 3600 3204 3618
rect 3186 3618 3204 3636
rect 3186 3636 3204 3654
rect 3186 3654 3204 3672
rect 3186 3672 3204 3690
rect 3186 3690 3204 3708
rect 3186 3708 3204 3726
rect 3186 3726 3204 3744
rect 3186 3744 3204 3762
rect 3186 3762 3204 3780
rect 3186 3780 3204 3798
rect 3186 3798 3204 3816
rect 3186 3816 3204 3834
rect 3186 3834 3204 3852
rect 3186 3852 3204 3870
rect 3186 3870 3204 3888
rect 3186 3888 3204 3906
rect 3186 3906 3204 3924
rect 3186 3924 3204 3942
rect 3186 3942 3204 3960
rect 3186 6606 3204 6624
rect 3186 6624 3204 6642
rect 3186 6642 3204 6660
rect 3186 6660 3204 6678
rect 3186 6678 3204 6696
rect 3186 6696 3204 6714
rect 3186 6714 3204 6732
rect 3186 6732 3204 6750
rect 3186 6750 3204 6768
rect 3186 6768 3204 6786
rect 3186 6786 3204 6804
rect 3186 6804 3204 6822
rect 3186 6822 3204 6840
rect 3186 6840 3204 6858
rect 3186 6858 3204 6876
rect 3186 6876 3204 6894
rect 3186 6894 3204 6912
rect 3186 6912 3204 6930
rect 3186 6930 3204 6948
rect 3186 6948 3204 6966
rect 3186 6966 3204 6984
rect 3186 6984 3204 7002
rect 3186 7002 3204 7020
rect 3186 7020 3204 7038
rect 3186 7038 3204 7056
rect 3186 7056 3204 7074
rect 3186 7074 3204 7092
rect 3186 7092 3204 7110
rect 3186 7110 3204 7128
rect 3186 7128 3204 7146
rect 3186 7146 3204 7164
rect 3186 7164 3204 7182
rect 3186 7182 3204 7200
rect 3186 7200 3204 7218
rect 3186 7218 3204 7236
rect 3204 54 3222 72
rect 3204 72 3222 90
rect 3204 90 3222 108
rect 3204 108 3222 126
rect 3204 126 3222 144
rect 3204 144 3222 162
rect 3204 162 3222 180
rect 3204 180 3222 198
rect 3204 198 3222 216
rect 3204 216 3222 234
rect 3204 234 3222 252
rect 3204 252 3222 270
rect 3204 270 3222 288
rect 3204 288 3222 306
rect 3204 306 3222 324
rect 3204 324 3222 342
rect 3204 342 3222 360
rect 3204 360 3222 378
rect 3204 378 3222 396
rect 3204 396 3222 414
rect 3204 414 3222 432
rect 3204 432 3222 450
rect 3204 450 3222 468
rect 3204 468 3222 486
rect 3204 486 3222 504
rect 3204 504 3222 522
rect 3204 522 3222 540
rect 3204 540 3222 558
rect 3204 558 3222 576
rect 3204 684 3222 702
rect 3204 702 3222 720
rect 3204 720 3222 738
rect 3204 738 3222 756
rect 3204 756 3222 774
rect 3204 774 3222 792
rect 3204 792 3222 810
rect 3204 810 3222 828
rect 3204 828 3222 846
rect 3204 846 3222 864
rect 3204 864 3222 882
rect 3204 882 3222 900
rect 3204 900 3222 918
rect 3204 918 3222 936
rect 3204 936 3222 954
rect 3204 954 3222 972
rect 3204 972 3222 990
rect 3204 990 3222 1008
rect 3204 1188 3222 1206
rect 3204 1206 3222 1224
rect 3204 1224 3222 1242
rect 3204 1242 3222 1260
rect 3204 1260 3222 1278
rect 3204 1278 3222 1296
rect 3204 1296 3222 1314
rect 3204 1314 3222 1332
rect 3204 1332 3222 1350
rect 3204 1350 3222 1368
rect 3204 1368 3222 1386
rect 3204 1386 3222 1404
rect 3204 1404 3222 1422
rect 3204 1422 3222 1440
rect 3204 1440 3222 1458
rect 3204 1458 3222 1476
rect 3204 1476 3222 1494
rect 3204 1494 3222 1512
rect 3204 1512 3222 1530
rect 3204 1530 3222 1548
rect 3204 1548 3222 1566
rect 3204 1566 3222 1584
rect 3204 1584 3222 1602
rect 3204 1602 3222 1620
rect 3204 1620 3222 1638
rect 3204 1638 3222 1656
rect 3204 1656 3222 1674
rect 3204 1674 3222 1692
rect 3204 1692 3222 1710
rect 3204 1710 3222 1728
rect 3204 1728 3222 1746
rect 3204 1746 3222 1764
rect 3204 1764 3222 1782
rect 3204 1782 3222 1800
rect 3204 1800 3222 1818
rect 3204 1818 3222 1836
rect 3204 2124 3222 2142
rect 3204 2142 3222 2160
rect 3204 2160 3222 2178
rect 3204 2178 3222 2196
rect 3204 2196 3222 2214
rect 3204 2214 3222 2232
rect 3204 2232 3222 2250
rect 3204 2250 3222 2268
rect 3204 2268 3222 2286
rect 3204 2286 3222 2304
rect 3204 2304 3222 2322
rect 3204 2322 3222 2340
rect 3204 2340 3222 2358
rect 3204 2358 3222 2376
rect 3204 2376 3222 2394
rect 3204 2394 3222 2412
rect 3204 2412 3222 2430
rect 3204 2430 3222 2448
rect 3204 2448 3222 2466
rect 3204 2466 3222 2484
rect 3204 2484 3222 2502
rect 3204 2502 3222 2520
rect 3204 2520 3222 2538
rect 3204 2538 3222 2556
rect 3204 2556 3222 2574
rect 3204 2574 3222 2592
rect 3204 2592 3222 2610
rect 3204 2610 3222 2628
rect 3204 2628 3222 2646
rect 3204 2646 3222 2664
rect 3204 2664 3222 2682
rect 3204 2682 3222 2700
rect 3204 2700 3222 2718
rect 3204 2718 3222 2736
rect 3204 2736 3222 2754
rect 3204 2754 3222 2772
rect 3204 2772 3222 2790
rect 3204 2790 3222 2808
rect 3204 2808 3222 2826
rect 3204 2826 3222 2844
rect 3204 2844 3222 2862
rect 3204 2862 3222 2880
rect 3204 2880 3222 2898
rect 3204 2898 3222 2916
rect 3204 2916 3222 2934
rect 3204 2934 3222 2952
rect 3204 2952 3222 2970
rect 3204 2970 3222 2988
rect 3204 2988 3222 3006
rect 3204 3006 3222 3024
rect 3204 3024 3222 3042
rect 3204 3042 3222 3060
rect 3204 3060 3222 3078
rect 3204 3078 3222 3096
rect 3204 3096 3222 3114
rect 3204 3114 3222 3132
rect 3204 3132 3222 3150
rect 3204 3150 3222 3168
rect 3204 3168 3222 3186
rect 3204 3186 3222 3204
rect 3204 3204 3222 3222
rect 3204 3222 3222 3240
rect 3204 3240 3222 3258
rect 3204 3258 3222 3276
rect 3204 3276 3222 3294
rect 3204 3294 3222 3312
rect 3204 3312 3222 3330
rect 3204 3330 3222 3348
rect 3204 3348 3222 3366
rect 3204 3366 3222 3384
rect 3204 3384 3222 3402
rect 3204 3402 3222 3420
rect 3204 3420 3222 3438
rect 3204 3438 3222 3456
rect 3204 3456 3222 3474
rect 3204 3474 3222 3492
rect 3204 3492 3222 3510
rect 3204 3510 3222 3528
rect 3204 3528 3222 3546
rect 3204 3546 3222 3564
rect 3204 3564 3222 3582
rect 3204 3582 3222 3600
rect 3204 3600 3222 3618
rect 3204 3618 3222 3636
rect 3204 3636 3222 3654
rect 3204 3654 3222 3672
rect 3204 3672 3222 3690
rect 3204 3690 3222 3708
rect 3204 3708 3222 3726
rect 3204 3726 3222 3744
rect 3204 3744 3222 3762
rect 3204 3762 3222 3780
rect 3204 3780 3222 3798
rect 3204 3798 3222 3816
rect 3204 3816 3222 3834
rect 3204 3834 3222 3852
rect 3204 3852 3222 3870
rect 3204 3870 3222 3888
rect 3204 3888 3222 3906
rect 3204 3906 3222 3924
rect 3204 3924 3222 3942
rect 3204 3942 3222 3960
rect 3204 3960 3222 3978
rect 3204 3978 3222 3996
rect 3204 3996 3222 4014
rect 3204 6624 3222 6642
rect 3204 6642 3222 6660
rect 3204 6660 3222 6678
rect 3204 6678 3222 6696
rect 3204 6696 3222 6714
rect 3204 6714 3222 6732
rect 3204 6732 3222 6750
rect 3204 6750 3222 6768
rect 3204 6768 3222 6786
rect 3204 6786 3222 6804
rect 3204 6804 3222 6822
rect 3204 6822 3222 6840
rect 3204 6840 3222 6858
rect 3204 6858 3222 6876
rect 3204 6876 3222 6894
rect 3204 6894 3222 6912
rect 3204 6912 3222 6930
rect 3204 6930 3222 6948
rect 3204 6948 3222 6966
rect 3204 6966 3222 6984
rect 3204 6984 3222 7002
rect 3204 7002 3222 7020
rect 3204 7020 3222 7038
rect 3204 7038 3222 7056
rect 3204 7056 3222 7074
rect 3204 7074 3222 7092
rect 3204 7092 3222 7110
rect 3204 7110 3222 7128
rect 3204 7128 3222 7146
rect 3204 7146 3222 7164
rect 3204 7164 3222 7182
rect 3204 7182 3222 7200
rect 3204 7200 3222 7218
rect 3204 7218 3222 7236
rect 3204 7236 3222 7254
rect 3222 54 3240 72
rect 3222 72 3240 90
rect 3222 90 3240 108
rect 3222 108 3240 126
rect 3222 126 3240 144
rect 3222 144 3240 162
rect 3222 162 3240 180
rect 3222 180 3240 198
rect 3222 198 3240 216
rect 3222 216 3240 234
rect 3222 234 3240 252
rect 3222 252 3240 270
rect 3222 270 3240 288
rect 3222 288 3240 306
rect 3222 306 3240 324
rect 3222 324 3240 342
rect 3222 342 3240 360
rect 3222 360 3240 378
rect 3222 378 3240 396
rect 3222 396 3240 414
rect 3222 414 3240 432
rect 3222 432 3240 450
rect 3222 450 3240 468
rect 3222 468 3240 486
rect 3222 486 3240 504
rect 3222 504 3240 522
rect 3222 522 3240 540
rect 3222 540 3240 558
rect 3222 558 3240 576
rect 3222 702 3240 720
rect 3222 720 3240 738
rect 3222 738 3240 756
rect 3222 756 3240 774
rect 3222 774 3240 792
rect 3222 792 3240 810
rect 3222 810 3240 828
rect 3222 828 3240 846
rect 3222 846 3240 864
rect 3222 864 3240 882
rect 3222 882 3240 900
rect 3222 900 3240 918
rect 3222 918 3240 936
rect 3222 936 3240 954
rect 3222 954 3240 972
rect 3222 972 3240 990
rect 3222 990 3240 1008
rect 3222 1008 3240 1026
rect 3222 1206 3240 1224
rect 3222 1224 3240 1242
rect 3222 1242 3240 1260
rect 3222 1260 3240 1278
rect 3222 1278 3240 1296
rect 3222 1296 3240 1314
rect 3222 1314 3240 1332
rect 3222 1332 3240 1350
rect 3222 1350 3240 1368
rect 3222 1368 3240 1386
rect 3222 1386 3240 1404
rect 3222 1404 3240 1422
rect 3222 1422 3240 1440
rect 3222 1440 3240 1458
rect 3222 1458 3240 1476
rect 3222 1476 3240 1494
rect 3222 1494 3240 1512
rect 3222 1512 3240 1530
rect 3222 1530 3240 1548
rect 3222 1548 3240 1566
rect 3222 1566 3240 1584
rect 3222 1584 3240 1602
rect 3222 1602 3240 1620
rect 3222 1620 3240 1638
rect 3222 1638 3240 1656
rect 3222 1656 3240 1674
rect 3222 1674 3240 1692
rect 3222 1692 3240 1710
rect 3222 1710 3240 1728
rect 3222 1728 3240 1746
rect 3222 1746 3240 1764
rect 3222 1764 3240 1782
rect 3222 1782 3240 1800
rect 3222 1800 3240 1818
rect 3222 1818 3240 1836
rect 3222 1836 3240 1854
rect 3222 1854 3240 1872
rect 3222 2160 3240 2178
rect 3222 2178 3240 2196
rect 3222 2196 3240 2214
rect 3222 2214 3240 2232
rect 3222 2232 3240 2250
rect 3222 2250 3240 2268
rect 3222 2268 3240 2286
rect 3222 2286 3240 2304
rect 3222 2304 3240 2322
rect 3222 2322 3240 2340
rect 3222 2340 3240 2358
rect 3222 2358 3240 2376
rect 3222 2376 3240 2394
rect 3222 2394 3240 2412
rect 3222 2412 3240 2430
rect 3222 2430 3240 2448
rect 3222 2448 3240 2466
rect 3222 2466 3240 2484
rect 3222 2484 3240 2502
rect 3222 2502 3240 2520
rect 3222 2520 3240 2538
rect 3222 2538 3240 2556
rect 3222 2556 3240 2574
rect 3222 2574 3240 2592
rect 3222 2592 3240 2610
rect 3222 2610 3240 2628
rect 3222 2628 3240 2646
rect 3222 2646 3240 2664
rect 3222 2664 3240 2682
rect 3222 2682 3240 2700
rect 3222 2700 3240 2718
rect 3222 2718 3240 2736
rect 3222 2736 3240 2754
rect 3222 2754 3240 2772
rect 3222 2772 3240 2790
rect 3222 2790 3240 2808
rect 3222 2808 3240 2826
rect 3222 2826 3240 2844
rect 3222 2844 3240 2862
rect 3222 2862 3240 2880
rect 3222 2880 3240 2898
rect 3222 2898 3240 2916
rect 3222 2916 3240 2934
rect 3222 2934 3240 2952
rect 3222 2952 3240 2970
rect 3222 2970 3240 2988
rect 3222 2988 3240 3006
rect 3222 3006 3240 3024
rect 3222 3024 3240 3042
rect 3222 3042 3240 3060
rect 3222 3060 3240 3078
rect 3222 3078 3240 3096
rect 3222 3096 3240 3114
rect 3222 3114 3240 3132
rect 3222 3132 3240 3150
rect 3222 3150 3240 3168
rect 3222 3168 3240 3186
rect 3222 3186 3240 3204
rect 3222 3204 3240 3222
rect 3222 3222 3240 3240
rect 3222 3240 3240 3258
rect 3222 3258 3240 3276
rect 3222 3276 3240 3294
rect 3222 3294 3240 3312
rect 3222 3312 3240 3330
rect 3222 3330 3240 3348
rect 3222 3348 3240 3366
rect 3222 3366 3240 3384
rect 3222 3384 3240 3402
rect 3222 3402 3240 3420
rect 3222 3420 3240 3438
rect 3222 3438 3240 3456
rect 3222 3456 3240 3474
rect 3222 3474 3240 3492
rect 3222 3492 3240 3510
rect 3222 3510 3240 3528
rect 3222 3528 3240 3546
rect 3222 3546 3240 3564
rect 3222 3564 3240 3582
rect 3222 3582 3240 3600
rect 3222 3600 3240 3618
rect 3222 3618 3240 3636
rect 3222 3636 3240 3654
rect 3222 3654 3240 3672
rect 3222 3672 3240 3690
rect 3222 3690 3240 3708
rect 3222 3708 3240 3726
rect 3222 3726 3240 3744
rect 3222 3744 3240 3762
rect 3222 3762 3240 3780
rect 3222 3780 3240 3798
rect 3222 3798 3240 3816
rect 3222 3816 3240 3834
rect 3222 3834 3240 3852
rect 3222 3852 3240 3870
rect 3222 3870 3240 3888
rect 3222 3888 3240 3906
rect 3222 3906 3240 3924
rect 3222 3924 3240 3942
rect 3222 3942 3240 3960
rect 3222 3960 3240 3978
rect 3222 3978 3240 3996
rect 3222 3996 3240 4014
rect 3222 4014 3240 4032
rect 3222 4032 3240 4050
rect 3222 4050 3240 4068
rect 3222 4068 3240 4086
rect 3222 6624 3240 6642
rect 3222 6642 3240 6660
rect 3222 6660 3240 6678
rect 3222 6678 3240 6696
rect 3222 6696 3240 6714
rect 3222 6714 3240 6732
rect 3222 6732 3240 6750
rect 3222 6750 3240 6768
rect 3222 6768 3240 6786
rect 3222 6786 3240 6804
rect 3222 6804 3240 6822
rect 3222 6822 3240 6840
rect 3222 6840 3240 6858
rect 3222 6858 3240 6876
rect 3222 6876 3240 6894
rect 3222 6894 3240 6912
rect 3222 6912 3240 6930
rect 3222 6930 3240 6948
rect 3222 6948 3240 6966
rect 3222 6966 3240 6984
rect 3222 6984 3240 7002
rect 3222 7002 3240 7020
rect 3222 7020 3240 7038
rect 3222 7038 3240 7056
rect 3222 7056 3240 7074
rect 3222 7074 3240 7092
rect 3222 7092 3240 7110
rect 3222 7110 3240 7128
rect 3222 7128 3240 7146
rect 3222 7146 3240 7164
rect 3222 7164 3240 7182
rect 3222 7182 3240 7200
rect 3222 7200 3240 7218
rect 3222 7218 3240 7236
rect 3222 7236 3240 7254
rect 3240 36 3258 54
rect 3240 54 3258 72
rect 3240 72 3258 90
rect 3240 90 3258 108
rect 3240 108 3258 126
rect 3240 126 3258 144
rect 3240 144 3258 162
rect 3240 162 3258 180
rect 3240 180 3258 198
rect 3240 198 3258 216
rect 3240 216 3258 234
rect 3240 234 3258 252
rect 3240 252 3258 270
rect 3240 270 3258 288
rect 3240 288 3258 306
rect 3240 306 3258 324
rect 3240 324 3258 342
rect 3240 342 3258 360
rect 3240 360 3258 378
rect 3240 378 3258 396
rect 3240 396 3258 414
rect 3240 414 3258 432
rect 3240 432 3258 450
rect 3240 450 3258 468
rect 3240 468 3258 486
rect 3240 486 3258 504
rect 3240 504 3258 522
rect 3240 522 3258 540
rect 3240 540 3258 558
rect 3240 558 3258 576
rect 3240 576 3258 594
rect 3240 720 3258 738
rect 3240 738 3258 756
rect 3240 756 3258 774
rect 3240 774 3258 792
rect 3240 792 3258 810
rect 3240 810 3258 828
rect 3240 828 3258 846
rect 3240 846 3258 864
rect 3240 864 3258 882
rect 3240 882 3258 900
rect 3240 900 3258 918
rect 3240 918 3258 936
rect 3240 936 3258 954
rect 3240 954 3258 972
rect 3240 972 3258 990
rect 3240 990 3258 1008
rect 3240 1008 3258 1026
rect 3240 1026 3258 1044
rect 3240 1224 3258 1242
rect 3240 1242 3258 1260
rect 3240 1260 3258 1278
rect 3240 1278 3258 1296
rect 3240 1296 3258 1314
rect 3240 1314 3258 1332
rect 3240 1332 3258 1350
rect 3240 1350 3258 1368
rect 3240 1368 3258 1386
rect 3240 1386 3258 1404
rect 3240 1404 3258 1422
rect 3240 1422 3258 1440
rect 3240 1440 3258 1458
rect 3240 1458 3258 1476
rect 3240 1476 3258 1494
rect 3240 1494 3258 1512
rect 3240 1512 3258 1530
rect 3240 1530 3258 1548
rect 3240 1548 3258 1566
rect 3240 1566 3258 1584
rect 3240 1584 3258 1602
rect 3240 1602 3258 1620
rect 3240 1620 3258 1638
rect 3240 1638 3258 1656
rect 3240 1656 3258 1674
rect 3240 1674 3258 1692
rect 3240 1692 3258 1710
rect 3240 1710 3258 1728
rect 3240 1728 3258 1746
rect 3240 1746 3258 1764
rect 3240 1764 3258 1782
rect 3240 1782 3258 1800
rect 3240 1800 3258 1818
rect 3240 1818 3258 1836
rect 3240 1836 3258 1854
rect 3240 1854 3258 1872
rect 3240 1872 3258 1890
rect 3240 1890 3258 1908
rect 3240 2196 3258 2214
rect 3240 2214 3258 2232
rect 3240 2232 3258 2250
rect 3240 2250 3258 2268
rect 3240 2268 3258 2286
rect 3240 2286 3258 2304
rect 3240 2304 3258 2322
rect 3240 2322 3258 2340
rect 3240 2340 3258 2358
rect 3240 2358 3258 2376
rect 3240 2376 3258 2394
rect 3240 2394 3258 2412
rect 3240 2412 3258 2430
rect 3240 2430 3258 2448
rect 3240 2448 3258 2466
rect 3240 2466 3258 2484
rect 3240 2484 3258 2502
rect 3240 2502 3258 2520
rect 3240 2520 3258 2538
rect 3240 2538 3258 2556
rect 3240 2556 3258 2574
rect 3240 2574 3258 2592
rect 3240 2592 3258 2610
rect 3240 2610 3258 2628
rect 3240 2628 3258 2646
rect 3240 2646 3258 2664
rect 3240 2664 3258 2682
rect 3240 2682 3258 2700
rect 3240 2700 3258 2718
rect 3240 2718 3258 2736
rect 3240 2736 3258 2754
rect 3240 2754 3258 2772
rect 3240 2772 3258 2790
rect 3240 2790 3258 2808
rect 3240 2808 3258 2826
rect 3240 2826 3258 2844
rect 3240 2844 3258 2862
rect 3240 2862 3258 2880
rect 3240 2880 3258 2898
rect 3240 2898 3258 2916
rect 3240 2916 3258 2934
rect 3240 2934 3258 2952
rect 3240 2952 3258 2970
rect 3240 2970 3258 2988
rect 3240 2988 3258 3006
rect 3240 3006 3258 3024
rect 3240 3024 3258 3042
rect 3240 3042 3258 3060
rect 3240 3060 3258 3078
rect 3240 3078 3258 3096
rect 3240 3096 3258 3114
rect 3240 3114 3258 3132
rect 3240 3132 3258 3150
rect 3240 3150 3258 3168
rect 3240 3168 3258 3186
rect 3240 3186 3258 3204
rect 3240 3204 3258 3222
rect 3240 3222 3258 3240
rect 3240 3240 3258 3258
rect 3240 3258 3258 3276
rect 3240 3276 3258 3294
rect 3240 3294 3258 3312
rect 3240 3312 3258 3330
rect 3240 3330 3258 3348
rect 3240 3348 3258 3366
rect 3240 3366 3258 3384
rect 3240 3384 3258 3402
rect 3240 3402 3258 3420
rect 3240 3420 3258 3438
rect 3240 3438 3258 3456
rect 3240 3456 3258 3474
rect 3240 3474 3258 3492
rect 3240 3492 3258 3510
rect 3240 3510 3258 3528
rect 3240 3528 3258 3546
rect 3240 3546 3258 3564
rect 3240 3564 3258 3582
rect 3240 3582 3258 3600
rect 3240 3600 3258 3618
rect 3240 3618 3258 3636
rect 3240 3636 3258 3654
rect 3240 3654 3258 3672
rect 3240 3672 3258 3690
rect 3240 3690 3258 3708
rect 3240 3708 3258 3726
rect 3240 3726 3258 3744
rect 3240 3744 3258 3762
rect 3240 3762 3258 3780
rect 3240 3780 3258 3798
rect 3240 3798 3258 3816
rect 3240 3816 3258 3834
rect 3240 3834 3258 3852
rect 3240 3852 3258 3870
rect 3240 3870 3258 3888
rect 3240 3888 3258 3906
rect 3240 3906 3258 3924
rect 3240 3924 3258 3942
rect 3240 3942 3258 3960
rect 3240 3960 3258 3978
rect 3240 3978 3258 3996
rect 3240 3996 3258 4014
rect 3240 4014 3258 4032
rect 3240 4032 3258 4050
rect 3240 4050 3258 4068
rect 3240 4068 3258 4086
rect 3240 4086 3258 4104
rect 3240 4104 3258 4122
rect 3240 4122 3258 4140
rect 3240 6624 3258 6642
rect 3240 6642 3258 6660
rect 3240 6660 3258 6678
rect 3240 6678 3258 6696
rect 3240 6696 3258 6714
rect 3240 6714 3258 6732
rect 3240 6732 3258 6750
rect 3240 6750 3258 6768
rect 3240 6768 3258 6786
rect 3240 6786 3258 6804
rect 3240 6804 3258 6822
rect 3240 6822 3258 6840
rect 3240 6840 3258 6858
rect 3240 6858 3258 6876
rect 3240 6876 3258 6894
rect 3240 6894 3258 6912
rect 3240 6912 3258 6930
rect 3240 6930 3258 6948
rect 3240 6948 3258 6966
rect 3240 6966 3258 6984
rect 3240 6984 3258 7002
rect 3240 7002 3258 7020
rect 3240 7020 3258 7038
rect 3240 7038 3258 7056
rect 3240 7056 3258 7074
rect 3240 7074 3258 7092
rect 3240 7092 3258 7110
rect 3240 7110 3258 7128
rect 3240 7128 3258 7146
rect 3240 7146 3258 7164
rect 3240 7164 3258 7182
rect 3240 7182 3258 7200
rect 3240 7200 3258 7218
rect 3240 7218 3258 7236
rect 3240 7236 3258 7254
rect 3258 36 3276 54
rect 3258 54 3276 72
rect 3258 72 3276 90
rect 3258 90 3276 108
rect 3258 108 3276 126
rect 3258 126 3276 144
rect 3258 144 3276 162
rect 3258 162 3276 180
rect 3258 180 3276 198
rect 3258 198 3276 216
rect 3258 216 3276 234
rect 3258 234 3276 252
rect 3258 252 3276 270
rect 3258 270 3276 288
rect 3258 288 3276 306
rect 3258 306 3276 324
rect 3258 324 3276 342
rect 3258 342 3276 360
rect 3258 360 3276 378
rect 3258 378 3276 396
rect 3258 396 3276 414
rect 3258 414 3276 432
rect 3258 432 3276 450
rect 3258 450 3276 468
rect 3258 468 3276 486
rect 3258 486 3276 504
rect 3258 504 3276 522
rect 3258 522 3276 540
rect 3258 540 3276 558
rect 3258 558 3276 576
rect 3258 576 3276 594
rect 3258 594 3276 612
rect 3258 720 3276 738
rect 3258 738 3276 756
rect 3258 756 3276 774
rect 3258 774 3276 792
rect 3258 792 3276 810
rect 3258 810 3276 828
rect 3258 828 3276 846
rect 3258 846 3276 864
rect 3258 864 3276 882
rect 3258 882 3276 900
rect 3258 900 3276 918
rect 3258 918 3276 936
rect 3258 936 3276 954
rect 3258 954 3276 972
rect 3258 972 3276 990
rect 3258 990 3276 1008
rect 3258 1008 3276 1026
rect 3258 1026 3276 1044
rect 3258 1242 3276 1260
rect 3258 1260 3276 1278
rect 3258 1278 3276 1296
rect 3258 1296 3276 1314
rect 3258 1314 3276 1332
rect 3258 1332 3276 1350
rect 3258 1350 3276 1368
rect 3258 1368 3276 1386
rect 3258 1386 3276 1404
rect 3258 1404 3276 1422
rect 3258 1422 3276 1440
rect 3258 1440 3276 1458
rect 3258 1458 3276 1476
rect 3258 1476 3276 1494
rect 3258 1494 3276 1512
rect 3258 1512 3276 1530
rect 3258 1530 3276 1548
rect 3258 1548 3276 1566
rect 3258 1566 3276 1584
rect 3258 1584 3276 1602
rect 3258 1602 3276 1620
rect 3258 1620 3276 1638
rect 3258 1638 3276 1656
rect 3258 1656 3276 1674
rect 3258 1674 3276 1692
rect 3258 1692 3276 1710
rect 3258 1710 3276 1728
rect 3258 1728 3276 1746
rect 3258 1746 3276 1764
rect 3258 1764 3276 1782
rect 3258 1782 3276 1800
rect 3258 1800 3276 1818
rect 3258 1818 3276 1836
rect 3258 1836 3276 1854
rect 3258 1854 3276 1872
rect 3258 1872 3276 1890
rect 3258 1890 3276 1908
rect 3258 1908 3276 1926
rect 3258 1926 3276 1944
rect 3258 2214 3276 2232
rect 3258 2232 3276 2250
rect 3258 2250 3276 2268
rect 3258 2268 3276 2286
rect 3258 2286 3276 2304
rect 3258 2304 3276 2322
rect 3258 2322 3276 2340
rect 3258 2340 3276 2358
rect 3258 2358 3276 2376
rect 3258 2376 3276 2394
rect 3258 2394 3276 2412
rect 3258 2412 3276 2430
rect 3258 2430 3276 2448
rect 3258 2448 3276 2466
rect 3258 2466 3276 2484
rect 3258 2484 3276 2502
rect 3258 2502 3276 2520
rect 3258 2520 3276 2538
rect 3258 2538 3276 2556
rect 3258 2556 3276 2574
rect 3258 2574 3276 2592
rect 3258 2592 3276 2610
rect 3258 2610 3276 2628
rect 3258 2628 3276 2646
rect 3258 2646 3276 2664
rect 3258 2664 3276 2682
rect 3258 2682 3276 2700
rect 3258 2700 3276 2718
rect 3258 2718 3276 2736
rect 3258 2736 3276 2754
rect 3258 2754 3276 2772
rect 3258 2772 3276 2790
rect 3258 2790 3276 2808
rect 3258 2808 3276 2826
rect 3258 2826 3276 2844
rect 3258 2844 3276 2862
rect 3258 2862 3276 2880
rect 3258 2880 3276 2898
rect 3258 2898 3276 2916
rect 3258 2916 3276 2934
rect 3258 2934 3276 2952
rect 3258 2952 3276 2970
rect 3258 2970 3276 2988
rect 3258 2988 3276 3006
rect 3258 3006 3276 3024
rect 3258 3024 3276 3042
rect 3258 3042 3276 3060
rect 3258 3060 3276 3078
rect 3258 3078 3276 3096
rect 3258 3096 3276 3114
rect 3258 3114 3276 3132
rect 3258 3132 3276 3150
rect 3258 3150 3276 3168
rect 3258 3168 3276 3186
rect 3258 3186 3276 3204
rect 3258 3204 3276 3222
rect 3258 3222 3276 3240
rect 3258 3240 3276 3258
rect 3258 3258 3276 3276
rect 3258 3276 3276 3294
rect 3258 3294 3276 3312
rect 3258 3312 3276 3330
rect 3258 3330 3276 3348
rect 3258 3348 3276 3366
rect 3258 3366 3276 3384
rect 3258 3384 3276 3402
rect 3258 3402 3276 3420
rect 3258 3420 3276 3438
rect 3258 3438 3276 3456
rect 3258 3456 3276 3474
rect 3258 3474 3276 3492
rect 3258 3492 3276 3510
rect 3258 3510 3276 3528
rect 3258 3528 3276 3546
rect 3258 3546 3276 3564
rect 3258 3564 3276 3582
rect 3258 3582 3276 3600
rect 3258 3600 3276 3618
rect 3258 3618 3276 3636
rect 3258 3636 3276 3654
rect 3258 3654 3276 3672
rect 3258 3672 3276 3690
rect 3258 3690 3276 3708
rect 3258 3708 3276 3726
rect 3258 3726 3276 3744
rect 3258 3744 3276 3762
rect 3258 3762 3276 3780
rect 3258 3780 3276 3798
rect 3258 3798 3276 3816
rect 3258 3816 3276 3834
rect 3258 3834 3276 3852
rect 3258 3852 3276 3870
rect 3258 3870 3276 3888
rect 3258 3888 3276 3906
rect 3258 3906 3276 3924
rect 3258 3924 3276 3942
rect 3258 3942 3276 3960
rect 3258 3960 3276 3978
rect 3258 3978 3276 3996
rect 3258 3996 3276 4014
rect 3258 4014 3276 4032
rect 3258 4032 3276 4050
rect 3258 4050 3276 4068
rect 3258 4068 3276 4086
rect 3258 4086 3276 4104
rect 3258 4104 3276 4122
rect 3258 4122 3276 4140
rect 3258 4140 3276 4158
rect 3258 4158 3276 4176
rect 3258 4176 3276 4194
rect 3258 6624 3276 6642
rect 3258 6642 3276 6660
rect 3258 6660 3276 6678
rect 3258 6678 3276 6696
rect 3258 6696 3276 6714
rect 3258 6714 3276 6732
rect 3258 6732 3276 6750
rect 3258 6750 3276 6768
rect 3258 6768 3276 6786
rect 3258 6786 3276 6804
rect 3258 6804 3276 6822
rect 3258 6822 3276 6840
rect 3258 6840 3276 6858
rect 3258 6858 3276 6876
rect 3258 6876 3276 6894
rect 3258 6894 3276 6912
rect 3258 6912 3276 6930
rect 3258 6930 3276 6948
rect 3258 6948 3276 6966
rect 3258 6966 3276 6984
rect 3258 6984 3276 7002
rect 3258 7002 3276 7020
rect 3258 7020 3276 7038
rect 3258 7038 3276 7056
rect 3258 7056 3276 7074
rect 3258 7074 3276 7092
rect 3258 7092 3276 7110
rect 3258 7110 3276 7128
rect 3258 7128 3276 7146
rect 3258 7146 3276 7164
rect 3258 7164 3276 7182
rect 3258 7182 3276 7200
rect 3258 7200 3276 7218
rect 3258 7218 3276 7236
rect 3258 7236 3276 7254
rect 3276 36 3294 54
rect 3276 54 3294 72
rect 3276 72 3294 90
rect 3276 90 3294 108
rect 3276 108 3294 126
rect 3276 126 3294 144
rect 3276 144 3294 162
rect 3276 162 3294 180
rect 3276 180 3294 198
rect 3276 198 3294 216
rect 3276 216 3294 234
rect 3276 234 3294 252
rect 3276 252 3294 270
rect 3276 270 3294 288
rect 3276 288 3294 306
rect 3276 306 3294 324
rect 3276 324 3294 342
rect 3276 342 3294 360
rect 3276 360 3294 378
rect 3276 378 3294 396
rect 3276 396 3294 414
rect 3276 414 3294 432
rect 3276 432 3294 450
rect 3276 450 3294 468
rect 3276 468 3294 486
rect 3276 486 3294 504
rect 3276 504 3294 522
rect 3276 522 3294 540
rect 3276 540 3294 558
rect 3276 558 3294 576
rect 3276 576 3294 594
rect 3276 594 3294 612
rect 3276 612 3294 630
rect 3276 720 3294 738
rect 3276 738 3294 756
rect 3276 756 3294 774
rect 3276 774 3294 792
rect 3276 792 3294 810
rect 3276 810 3294 828
rect 3276 828 3294 846
rect 3276 846 3294 864
rect 3276 864 3294 882
rect 3276 882 3294 900
rect 3276 900 3294 918
rect 3276 918 3294 936
rect 3276 936 3294 954
rect 3276 954 3294 972
rect 3276 972 3294 990
rect 3276 990 3294 1008
rect 3276 1008 3294 1026
rect 3276 1026 3294 1044
rect 3276 1044 3294 1062
rect 3276 1260 3294 1278
rect 3276 1278 3294 1296
rect 3276 1296 3294 1314
rect 3276 1314 3294 1332
rect 3276 1332 3294 1350
rect 3276 1350 3294 1368
rect 3276 1368 3294 1386
rect 3276 1386 3294 1404
rect 3276 1404 3294 1422
rect 3276 1422 3294 1440
rect 3276 1440 3294 1458
rect 3276 1458 3294 1476
rect 3276 1476 3294 1494
rect 3276 1494 3294 1512
rect 3276 1512 3294 1530
rect 3276 1530 3294 1548
rect 3276 1548 3294 1566
rect 3276 1566 3294 1584
rect 3276 1584 3294 1602
rect 3276 1602 3294 1620
rect 3276 1620 3294 1638
rect 3276 1638 3294 1656
rect 3276 1656 3294 1674
rect 3276 1674 3294 1692
rect 3276 1692 3294 1710
rect 3276 1710 3294 1728
rect 3276 1728 3294 1746
rect 3276 1746 3294 1764
rect 3276 1764 3294 1782
rect 3276 1782 3294 1800
rect 3276 1800 3294 1818
rect 3276 1818 3294 1836
rect 3276 1836 3294 1854
rect 3276 1854 3294 1872
rect 3276 1872 3294 1890
rect 3276 1890 3294 1908
rect 3276 1908 3294 1926
rect 3276 1926 3294 1944
rect 3276 1944 3294 1962
rect 3276 2250 3294 2268
rect 3276 2268 3294 2286
rect 3276 2286 3294 2304
rect 3276 2304 3294 2322
rect 3276 2322 3294 2340
rect 3276 2340 3294 2358
rect 3276 2358 3294 2376
rect 3276 2376 3294 2394
rect 3276 2394 3294 2412
rect 3276 2412 3294 2430
rect 3276 2430 3294 2448
rect 3276 2448 3294 2466
rect 3276 2466 3294 2484
rect 3276 2484 3294 2502
rect 3276 2502 3294 2520
rect 3276 2520 3294 2538
rect 3276 2538 3294 2556
rect 3276 2556 3294 2574
rect 3276 2574 3294 2592
rect 3276 2592 3294 2610
rect 3276 2610 3294 2628
rect 3276 2628 3294 2646
rect 3276 2646 3294 2664
rect 3276 2664 3294 2682
rect 3276 2682 3294 2700
rect 3276 2700 3294 2718
rect 3276 2718 3294 2736
rect 3276 2736 3294 2754
rect 3276 2754 3294 2772
rect 3276 2772 3294 2790
rect 3276 2790 3294 2808
rect 3276 2808 3294 2826
rect 3276 2826 3294 2844
rect 3276 2844 3294 2862
rect 3276 2862 3294 2880
rect 3276 2880 3294 2898
rect 3276 2898 3294 2916
rect 3276 2916 3294 2934
rect 3276 2934 3294 2952
rect 3276 2952 3294 2970
rect 3276 2970 3294 2988
rect 3276 2988 3294 3006
rect 3276 3006 3294 3024
rect 3276 3024 3294 3042
rect 3276 3042 3294 3060
rect 3276 3060 3294 3078
rect 3276 3078 3294 3096
rect 3276 3096 3294 3114
rect 3276 3114 3294 3132
rect 3276 3132 3294 3150
rect 3276 3150 3294 3168
rect 3276 3168 3294 3186
rect 3276 3186 3294 3204
rect 3276 3204 3294 3222
rect 3276 3222 3294 3240
rect 3276 3240 3294 3258
rect 3276 3258 3294 3276
rect 3276 3276 3294 3294
rect 3276 3294 3294 3312
rect 3276 3312 3294 3330
rect 3276 3330 3294 3348
rect 3276 3348 3294 3366
rect 3276 3366 3294 3384
rect 3276 3384 3294 3402
rect 3276 3402 3294 3420
rect 3276 3420 3294 3438
rect 3276 3438 3294 3456
rect 3276 3456 3294 3474
rect 3276 3474 3294 3492
rect 3276 3492 3294 3510
rect 3276 3510 3294 3528
rect 3276 3528 3294 3546
rect 3276 3546 3294 3564
rect 3276 3564 3294 3582
rect 3276 3582 3294 3600
rect 3276 3600 3294 3618
rect 3276 3618 3294 3636
rect 3276 3636 3294 3654
rect 3276 3654 3294 3672
rect 3276 3672 3294 3690
rect 3276 3690 3294 3708
rect 3276 3708 3294 3726
rect 3276 3726 3294 3744
rect 3276 3744 3294 3762
rect 3276 3762 3294 3780
rect 3276 3780 3294 3798
rect 3276 3798 3294 3816
rect 3276 3816 3294 3834
rect 3276 3834 3294 3852
rect 3276 3852 3294 3870
rect 3276 3870 3294 3888
rect 3276 3888 3294 3906
rect 3276 3906 3294 3924
rect 3276 3924 3294 3942
rect 3276 3942 3294 3960
rect 3276 3960 3294 3978
rect 3276 3978 3294 3996
rect 3276 3996 3294 4014
rect 3276 4014 3294 4032
rect 3276 4032 3294 4050
rect 3276 4050 3294 4068
rect 3276 4068 3294 4086
rect 3276 4086 3294 4104
rect 3276 4104 3294 4122
rect 3276 4122 3294 4140
rect 3276 4140 3294 4158
rect 3276 4158 3294 4176
rect 3276 4176 3294 4194
rect 3276 4194 3294 4212
rect 3276 4212 3294 4230
rect 3276 4230 3294 4248
rect 3276 6624 3294 6642
rect 3276 6642 3294 6660
rect 3276 6660 3294 6678
rect 3276 6678 3294 6696
rect 3276 6696 3294 6714
rect 3276 6714 3294 6732
rect 3276 6732 3294 6750
rect 3276 6750 3294 6768
rect 3276 6768 3294 6786
rect 3276 6786 3294 6804
rect 3276 6804 3294 6822
rect 3276 6822 3294 6840
rect 3276 6840 3294 6858
rect 3276 6858 3294 6876
rect 3276 6876 3294 6894
rect 3276 6894 3294 6912
rect 3276 6912 3294 6930
rect 3276 6930 3294 6948
rect 3276 6948 3294 6966
rect 3276 6966 3294 6984
rect 3276 6984 3294 7002
rect 3276 7002 3294 7020
rect 3276 7020 3294 7038
rect 3276 7038 3294 7056
rect 3276 7056 3294 7074
rect 3276 7074 3294 7092
rect 3276 7092 3294 7110
rect 3276 7110 3294 7128
rect 3276 7128 3294 7146
rect 3276 7146 3294 7164
rect 3276 7164 3294 7182
rect 3276 7182 3294 7200
rect 3276 7200 3294 7218
rect 3276 7218 3294 7236
rect 3276 7236 3294 7254
rect 3294 36 3312 54
rect 3294 54 3312 72
rect 3294 72 3312 90
rect 3294 90 3312 108
rect 3294 108 3312 126
rect 3294 126 3312 144
rect 3294 144 3312 162
rect 3294 162 3312 180
rect 3294 180 3312 198
rect 3294 198 3312 216
rect 3294 216 3312 234
rect 3294 234 3312 252
rect 3294 252 3312 270
rect 3294 270 3312 288
rect 3294 288 3312 306
rect 3294 306 3312 324
rect 3294 324 3312 342
rect 3294 342 3312 360
rect 3294 360 3312 378
rect 3294 378 3312 396
rect 3294 396 3312 414
rect 3294 414 3312 432
rect 3294 432 3312 450
rect 3294 450 3312 468
rect 3294 468 3312 486
rect 3294 486 3312 504
rect 3294 504 3312 522
rect 3294 522 3312 540
rect 3294 540 3312 558
rect 3294 558 3312 576
rect 3294 576 3312 594
rect 3294 594 3312 612
rect 3294 612 3312 630
rect 3294 738 3312 756
rect 3294 756 3312 774
rect 3294 774 3312 792
rect 3294 792 3312 810
rect 3294 810 3312 828
rect 3294 828 3312 846
rect 3294 846 3312 864
rect 3294 864 3312 882
rect 3294 882 3312 900
rect 3294 900 3312 918
rect 3294 918 3312 936
rect 3294 936 3312 954
rect 3294 954 3312 972
rect 3294 972 3312 990
rect 3294 990 3312 1008
rect 3294 1008 3312 1026
rect 3294 1026 3312 1044
rect 3294 1044 3312 1062
rect 3294 1062 3312 1080
rect 3294 1260 3312 1278
rect 3294 1278 3312 1296
rect 3294 1296 3312 1314
rect 3294 1314 3312 1332
rect 3294 1332 3312 1350
rect 3294 1350 3312 1368
rect 3294 1368 3312 1386
rect 3294 1386 3312 1404
rect 3294 1404 3312 1422
rect 3294 1422 3312 1440
rect 3294 1440 3312 1458
rect 3294 1458 3312 1476
rect 3294 1476 3312 1494
rect 3294 1494 3312 1512
rect 3294 1512 3312 1530
rect 3294 1530 3312 1548
rect 3294 1548 3312 1566
rect 3294 1566 3312 1584
rect 3294 1584 3312 1602
rect 3294 1602 3312 1620
rect 3294 1620 3312 1638
rect 3294 1638 3312 1656
rect 3294 1656 3312 1674
rect 3294 1674 3312 1692
rect 3294 1692 3312 1710
rect 3294 1710 3312 1728
rect 3294 1728 3312 1746
rect 3294 1746 3312 1764
rect 3294 1764 3312 1782
rect 3294 1782 3312 1800
rect 3294 1800 3312 1818
rect 3294 1818 3312 1836
rect 3294 1836 3312 1854
rect 3294 1854 3312 1872
rect 3294 1872 3312 1890
rect 3294 1890 3312 1908
rect 3294 1908 3312 1926
rect 3294 1926 3312 1944
rect 3294 1944 3312 1962
rect 3294 1962 3312 1980
rect 3294 1980 3312 1998
rect 3294 2268 3312 2286
rect 3294 2286 3312 2304
rect 3294 2304 3312 2322
rect 3294 2322 3312 2340
rect 3294 2340 3312 2358
rect 3294 2358 3312 2376
rect 3294 2376 3312 2394
rect 3294 2394 3312 2412
rect 3294 2412 3312 2430
rect 3294 2430 3312 2448
rect 3294 2448 3312 2466
rect 3294 2466 3312 2484
rect 3294 2484 3312 2502
rect 3294 2502 3312 2520
rect 3294 2520 3312 2538
rect 3294 2538 3312 2556
rect 3294 2556 3312 2574
rect 3294 2574 3312 2592
rect 3294 2592 3312 2610
rect 3294 2610 3312 2628
rect 3294 2628 3312 2646
rect 3294 2646 3312 2664
rect 3294 2664 3312 2682
rect 3294 2682 3312 2700
rect 3294 2700 3312 2718
rect 3294 2718 3312 2736
rect 3294 2736 3312 2754
rect 3294 2754 3312 2772
rect 3294 2772 3312 2790
rect 3294 2790 3312 2808
rect 3294 2808 3312 2826
rect 3294 2826 3312 2844
rect 3294 2844 3312 2862
rect 3294 2862 3312 2880
rect 3294 2880 3312 2898
rect 3294 2898 3312 2916
rect 3294 2916 3312 2934
rect 3294 2934 3312 2952
rect 3294 2952 3312 2970
rect 3294 2970 3312 2988
rect 3294 2988 3312 3006
rect 3294 3006 3312 3024
rect 3294 3024 3312 3042
rect 3294 3042 3312 3060
rect 3294 3060 3312 3078
rect 3294 3078 3312 3096
rect 3294 3096 3312 3114
rect 3294 3114 3312 3132
rect 3294 3132 3312 3150
rect 3294 3150 3312 3168
rect 3294 3168 3312 3186
rect 3294 3186 3312 3204
rect 3294 3204 3312 3222
rect 3294 3222 3312 3240
rect 3294 3240 3312 3258
rect 3294 3258 3312 3276
rect 3294 3276 3312 3294
rect 3294 3294 3312 3312
rect 3294 3312 3312 3330
rect 3294 3330 3312 3348
rect 3294 3348 3312 3366
rect 3294 3366 3312 3384
rect 3294 3384 3312 3402
rect 3294 3402 3312 3420
rect 3294 3420 3312 3438
rect 3294 3438 3312 3456
rect 3294 3456 3312 3474
rect 3294 3474 3312 3492
rect 3294 3492 3312 3510
rect 3294 3510 3312 3528
rect 3294 3528 3312 3546
rect 3294 3546 3312 3564
rect 3294 3564 3312 3582
rect 3294 3582 3312 3600
rect 3294 3600 3312 3618
rect 3294 3618 3312 3636
rect 3294 3636 3312 3654
rect 3294 3654 3312 3672
rect 3294 3672 3312 3690
rect 3294 3690 3312 3708
rect 3294 3708 3312 3726
rect 3294 3726 3312 3744
rect 3294 3744 3312 3762
rect 3294 3762 3312 3780
rect 3294 3780 3312 3798
rect 3294 3798 3312 3816
rect 3294 3816 3312 3834
rect 3294 3834 3312 3852
rect 3294 3852 3312 3870
rect 3294 3870 3312 3888
rect 3294 3888 3312 3906
rect 3294 3906 3312 3924
rect 3294 3924 3312 3942
rect 3294 3942 3312 3960
rect 3294 3960 3312 3978
rect 3294 3978 3312 3996
rect 3294 3996 3312 4014
rect 3294 4014 3312 4032
rect 3294 4032 3312 4050
rect 3294 4050 3312 4068
rect 3294 4068 3312 4086
rect 3294 4086 3312 4104
rect 3294 4104 3312 4122
rect 3294 4122 3312 4140
rect 3294 4140 3312 4158
rect 3294 4158 3312 4176
rect 3294 4176 3312 4194
rect 3294 4194 3312 4212
rect 3294 4212 3312 4230
rect 3294 4230 3312 4248
rect 3294 4248 3312 4266
rect 3294 4266 3312 4284
rect 3294 4284 3312 4302
rect 3294 6624 3312 6642
rect 3294 6642 3312 6660
rect 3294 6660 3312 6678
rect 3294 6678 3312 6696
rect 3294 6696 3312 6714
rect 3294 6714 3312 6732
rect 3294 6732 3312 6750
rect 3294 6750 3312 6768
rect 3294 6768 3312 6786
rect 3294 6786 3312 6804
rect 3294 6804 3312 6822
rect 3294 6822 3312 6840
rect 3294 6840 3312 6858
rect 3294 6858 3312 6876
rect 3294 6876 3312 6894
rect 3294 6894 3312 6912
rect 3294 6912 3312 6930
rect 3294 6930 3312 6948
rect 3294 6948 3312 6966
rect 3294 6966 3312 6984
rect 3294 6984 3312 7002
rect 3294 7002 3312 7020
rect 3294 7020 3312 7038
rect 3294 7038 3312 7056
rect 3294 7056 3312 7074
rect 3294 7074 3312 7092
rect 3294 7092 3312 7110
rect 3294 7110 3312 7128
rect 3294 7128 3312 7146
rect 3294 7146 3312 7164
rect 3294 7164 3312 7182
rect 3294 7182 3312 7200
rect 3294 7200 3312 7218
rect 3294 7218 3312 7236
rect 3294 7236 3312 7254
rect 3312 36 3330 54
rect 3312 54 3330 72
rect 3312 72 3330 90
rect 3312 90 3330 108
rect 3312 108 3330 126
rect 3312 126 3330 144
rect 3312 144 3330 162
rect 3312 162 3330 180
rect 3312 180 3330 198
rect 3312 198 3330 216
rect 3312 216 3330 234
rect 3312 234 3330 252
rect 3312 252 3330 270
rect 3312 270 3330 288
rect 3312 288 3330 306
rect 3312 306 3330 324
rect 3312 324 3330 342
rect 3312 342 3330 360
rect 3312 360 3330 378
rect 3312 378 3330 396
rect 3312 396 3330 414
rect 3312 414 3330 432
rect 3312 432 3330 450
rect 3312 450 3330 468
rect 3312 468 3330 486
rect 3312 486 3330 504
rect 3312 504 3330 522
rect 3312 522 3330 540
rect 3312 540 3330 558
rect 3312 558 3330 576
rect 3312 576 3330 594
rect 3312 594 3330 612
rect 3312 612 3330 630
rect 3312 738 3330 756
rect 3312 756 3330 774
rect 3312 774 3330 792
rect 3312 792 3330 810
rect 3312 810 3330 828
rect 3312 828 3330 846
rect 3312 846 3330 864
rect 3312 864 3330 882
rect 3312 882 3330 900
rect 3312 900 3330 918
rect 3312 918 3330 936
rect 3312 936 3330 954
rect 3312 954 3330 972
rect 3312 972 3330 990
rect 3312 990 3330 1008
rect 3312 1008 3330 1026
rect 3312 1026 3330 1044
rect 3312 1044 3330 1062
rect 3312 1062 3330 1080
rect 3312 1278 3330 1296
rect 3312 1296 3330 1314
rect 3312 1314 3330 1332
rect 3312 1332 3330 1350
rect 3312 1350 3330 1368
rect 3312 1368 3330 1386
rect 3312 1386 3330 1404
rect 3312 1404 3330 1422
rect 3312 1422 3330 1440
rect 3312 1440 3330 1458
rect 3312 1458 3330 1476
rect 3312 1476 3330 1494
rect 3312 1494 3330 1512
rect 3312 1512 3330 1530
rect 3312 1530 3330 1548
rect 3312 1548 3330 1566
rect 3312 1566 3330 1584
rect 3312 1584 3330 1602
rect 3312 1602 3330 1620
rect 3312 1620 3330 1638
rect 3312 1638 3330 1656
rect 3312 1656 3330 1674
rect 3312 1674 3330 1692
rect 3312 1692 3330 1710
rect 3312 1710 3330 1728
rect 3312 1728 3330 1746
rect 3312 1746 3330 1764
rect 3312 1764 3330 1782
rect 3312 1782 3330 1800
rect 3312 1800 3330 1818
rect 3312 1818 3330 1836
rect 3312 1836 3330 1854
rect 3312 1854 3330 1872
rect 3312 1872 3330 1890
rect 3312 1890 3330 1908
rect 3312 1908 3330 1926
rect 3312 1926 3330 1944
rect 3312 1944 3330 1962
rect 3312 1962 3330 1980
rect 3312 1980 3330 1998
rect 3312 1998 3330 2016
rect 3312 2016 3330 2034
rect 3312 2304 3330 2322
rect 3312 2322 3330 2340
rect 3312 2340 3330 2358
rect 3312 2358 3330 2376
rect 3312 2376 3330 2394
rect 3312 2394 3330 2412
rect 3312 2412 3330 2430
rect 3312 2430 3330 2448
rect 3312 2448 3330 2466
rect 3312 2466 3330 2484
rect 3312 2484 3330 2502
rect 3312 2502 3330 2520
rect 3312 2520 3330 2538
rect 3312 2538 3330 2556
rect 3312 2556 3330 2574
rect 3312 2574 3330 2592
rect 3312 2592 3330 2610
rect 3312 2610 3330 2628
rect 3312 2628 3330 2646
rect 3312 2646 3330 2664
rect 3312 2664 3330 2682
rect 3312 2682 3330 2700
rect 3312 2700 3330 2718
rect 3312 2718 3330 2736
rect 3312 2736 3330 2754
rect 3312 2754 3330 2772
rect 3312 2772 3330 2790
rect 3312 2790 3330 2808
rect 3312 2808 3330 2826
rect 3312 2826 3330 2844
rect 3312 2844 3330 2862
rect 3312 2862 3330 2880
rect 3312 2880 3330 2898
rect 3312 2898 3330 2916
rect 3312 2916 3330 2934
rect 3312 2934 3330 2952
rect 3312 2952 3330 2970
rect 3312 2970 3330 2988
rect 3312 2988 3330 3006
rect 3312 3006 3330 3024
rect 3312 3024 3330 3042
rect 3312 3042 3330 3060
rect 3312 3060 3330 3078
rect 3312 3078 3330 3096
rect 3312 3096 3330 3114
rect 3312 3114 3330 3132
rect 3312 3132 3330 3150
rect 3312 3150 3330 3168
rect 3312 3168 3330 3186
rect 3312 3186 3330 3204
rect 3312 3204 3330 3222
rect 3312 3222 3330 3240
rect 3312 3240 3330 3258
rect 3312 3258 3330 3276
rect 3312 3276 3330 3294
rect 3312 3294 3330 3312
rect 3312 3312 3330 3330
rect 3312 3330 3330 3348
rect 3312 3348 3330 3366
rect 3312 3366 3330 3384
rect 3312 3384 3330 3402
rect 3312 3402 3330 3420
rect 3312 3420 3330 3438
rect 3312 3438 3330 3456
rect 3312 3456 3330 3474
rect 3312 3474 3330 3492
rect 3312 3492 3330 3510
rect 3312 3510 3330 3528
rect 3312 3528 3330 3546
rect 3312 3546 3330 3564
rect 3312 3564 3330 3582
rect 3312 3582 3330 3600
rect 3312 3600 3330 3618
rect 3312 3618 3330 3636
rect 3312 3636 3330 3654
rect 3312 3654 3330 3672
rect 3312 3672 3330 3690
rect 3312 3690 3330 3708
rect 3312 3708 3330 3726
rect 3312 3726 3330 3744
rect 3312 3744 3330 3762
rect 3312 3762 3330 3780
rect 3312 3780 3330 3798
rect 3312 3798 3330 3816
rect 3312 3816 3330 3834
rect 3312 3834 3330 3852
rect 3312 3852 3330 3870
rect 3312 3870 3330 3888
rect 3312 3888 3330 3906
rect 3312 3906 3330 3924
rect 3312 3924 3330 3942
rect 3312 3942 3330 3960
rect 3312 3960 3330 3978
rect 3312 3978 3330 3996
rect 3312 3996 3330 4014
rect 3312 4014 3330 4032
rect 3312 4032 3330 4050
rect 3312 4050 3330 4068
rect 3312 4068 3330 4086
rect 3312 4086 3330 4104
rect 3312 4104 3330 4122
rect 3312 4122 3330 4140
rect 3312 4140 3330 4158
rect 3312 4158 3330 4176
rect 3312 4176 3330 4194
rect 3312 4194 3330 4212
rect 3312 4212 3330 4230
rect 3312 4230 3330 4248
rect 3312 4248 3330 4266
rect 3312 4266 3330 4284
rect 3312 4284 3330 4302
rect 3312 4302 3330 4320
rect 3312 4320 3330 4338
rect 3312 4338 3330 4356
rect 3312 6624 3330 6642
rect 3312 6642 3330 6660
rect 3312 6660 3330 6678
rect 3312 6678 3330 6696
rect 3312 6696 3330 6714
rect 3312 6714 3330 6732
rect 3312 6732 3330 6750
rect 3312 6750 3330 6768
rect 3312 6768 3330 6786
rect 3312 6786 3330 6804
rect 3312 6804 3330 6822
rect 3312 6822 3330 6840
rect 3312 6840 3330 6858
rect 3312 6858 3330 6876
rect 3312 6876 3330 6894
rect 3312 6894 3330 6912
rect 3312 6912 3330 6930
rect 3312 6930 3330 6948
rect 3312 6948 3330 6966
rect 3312 6966 3330 6984
rect 3312 6984 3330 7002
rect 3312 7002 3330 7020
rect 3312 7020 3330 7038
rect 3312 7038 3330 7056
rect 3312 7056 3330 7074
rect 3312 7074 3330 7092
rect 3312 7092 3330 7110
rect 3312 7110 3330 7128
rect 3312 7128 3330 7146
rect 3312 7146 3330 7164
rect 3312 7164 3330 7182
rect 3312 7182 3330 7200
rect 3312 7200 3330 7218
rect 3312 7218 3330 7236
rect 3312 7236 3330 7254
rect 3330 36 3348 54
rect 3330 54 3348 72
rect 3330 72 3348 90
rect 3330 90 3348 108
rect 3330 108 3348 126
rect 3330 126 3348 144
rect 3330 144 3348 162
rect 3330 162 3348 180
rect 3330 180 3348 198
rect 3330 198 3348 216
rect 3330 216 3348 234
rect 3330 234 3348 252
rect 3330 252 3348 270
rect 3330 270 3348 288
rect 3330 288 3348 306
rect 3330 306 3348 324
rect 3330 324 3348 342
rect 3330 342 3348 360
rect 3330 360 3348 378
rect 3330 378 3348 396
rect 3330 396 3348 414
rect 3330 414 3348 432
rect 3330 432 3348 450
rect 3330 450 3348 468
rect 3330 468 3348 486
rect 3330 486 3348 504
rect 3330 504 3348 522
rect 3330 522 3348 540
rect 3330 540 3348 558
rect 3330 558 3348 576
rect 3330 576 3348 594
rect 3330 594 3348 612
rect 3330 612 3348 630
rect 3330 756 3348 774
rect 3330 774 3348 792
rect 3330 792 3348 810
rect 3330 810 3348 828
rect 3330 828 3348 846
rect 3330 846 3348 864
rect 3330 864 3348 882
rect 3330 882 3348 900
rect 3330 900 3348 918
rect 3330 918 3348 936
rect 3330 936 3348 954
rect 3330 954 3348 972
rect 3330 972 3348 990
rect 3330 990 3348 1008
rect 3330 1008 3348 1026
rect 3330 1026 3348 1044
rect 3330 1044 3348 1062
rect 3330 1062 3348 1080
rect 3330 1080 3348 1098
rect 3330 1296 3348 1314
rect 3330 1314 3348 1332
rect 3330 1332 3348 1350
rect 3330 1350 3348 1368
rect 3330 1368 3348 1386
rect 3330 1386 3348 1404
rect 3330 1404 3348 1422
rect 3330 1422 3348 1440
rect 3330 1440 3348 1458
rect 3330 1458 3348 1476
rect 3330 1476 3348 1494
rect 3330 1494 3348 1512
rect 3330 1512 3348 1530
rect 3330 1530 3348 1548
rect 3330 1548 3348 1566
rect 3330 1566 3348 1584
rect 3330 1584 3348 1602
rect 3330 1602 3348 1620
rect 3330 1620 3348 1638
rect 3330 1638 3348 1656
rect 3330 1656 3348 1674
rect 3330 1674 3348 1692
rect 3330 1692 3348 1710
rect 3330 1710 3348 1728
rect 3330 1728 3348 1746
rect 3330 1746 3348 1764
rect 3330 1764 3348 1782
rect 3330 1782 3348 1800
rect 3330 1800 3348 1818
rect 3330 1818 3348 1836
rect 3330 1836 3348 1854
rect 3330 1854 3348 1872
rect 3330 1872 3348 1890
rect 3330 1890 3348 1908
rect 3330 1908 3348 1926
rect 3330 1926 3348 1944
rect 3330 1944 3348 1962
rect 3330 1962 3348 1980
rect 3330 1980 3348 1998
rect 3330 1998 3348 2016
rect 3330 2016 3348 2034
rect 3330 2034 3348 2052
rect 3330 2340 3348 2358
rect 3330 2358 3348 2376
rect 3330 2376 3348 2394
rect 3330 2394 3348 2412
rect 3330 2412 3348 2430
rect 3330 2430 3348 2448
rect 3330 2448 3348 2466
rect 3330 2466 3348 2484
rect 3330 2484 3348 2502
rect 3330 2502 3348 2520
rect 3330 2520 3348 2538
rect 3330 2538 3348 2556
rect 3330 2556 3348 2574
rect 3330 2574 3348 2592
rect 3330 2592 3348 2610
rect 3330 2610 3348 2628
rect 3330 2628 3348 2646
rect 3330 2646 3348 2664
rect 3330 2664 3348 2682
rect 3330 2682 3348 2700
rect 3330 2700 3348 2718
rect 3330 2718 3348 2736
rect 3330 2736 3348 2754
rect 3330 2754 3348 2772
rect 3330 2772 3348 2790
rect 3330 2790 3348 2808
rect 3330 2808 3348 2826
rect 3330 2826 3348 2844
rect 3330 2844 3348 2862
rect 3330 2862 3348 2880
rect 3330 2880 3348 2898
rect 3330 2898 3348 2916
rect 3330 2916 3348 2934
rect 3330 2934 3348 2952
rect 3330 2952 3348 2970
rect 3330 2970 3348 2988
rect 3330 2988 3348 3006
rect 3330 3006 3348 3024
rect 3330 3024 3348 3042
rect 3330 3042 3348 3060
rect 3330 3060 3348 3078
rect 3330 3078 3348 3096
rect 3330 3096 3348 3114
rect 3330 3114 3348 3132
rect 3330 3132 3348 3150
rect 3330 3150 3348 3168
rect 3330 3168 3348 3186
rect 3330 3186 3348 3204
rect 3330 3204 3348 3222
rect 3330 3222 3348 3240
rect 3330 3240 3348 3258
rect 3330 3258 3348 3276
rect 3330 3276 3348 3294
rect 3330 3294 3348 3312
rect 3330 3312 3348 3330
rect 3330 3330 3348 3348
rect 3330 3348 3348 3366
rect 3330 3366 3348 3384
rect 3330 3384 3348 3402
rect 3330 3402 3348 3420
rect 3330 3420 3348 3438
rect 3330 3438 3348 3456
rect 3330 3456 3348 3474
rect 3330 3474 3348 3492
rect 3330 3492 3348 3510
rect 3330 3510 3348 3528
rect 3330 3528 3348 3546
rect 3330 3546 3348 3564
rect 3330 3564 3348 3582
rect 3330 3582 3348 3600
rect 3330 3600 3348 3618
rect 3330 3618 3348 3636
rect 3330 3636 3348 3654
rect 3330 3654 3348 3672
rect 3330 3672 3348 3690
rect 3330 3690 3348 3708
rect 3330 3708 3348 3726
rect 3330 3726 3348 3744
rect 3330 3744 3348 3762
rect 3330 3762 3348 3780
rect 3330 3780 3348 3798
rect 3330 3798 3348 3816
rect 3330 3816 3348 3834
rect 3330 3834 3348 3852
rect 3330 3852 3348 3870
rect 3330 3870 3348 3888
rect 3330 3888 3348 3906
rect 3330 3906 3348 3924
rect 3330 3924 3348 3942
rect 3330 3942 3348 3960
rect 3330 3960 3348 3978
rect 3330 3978 3348 3996
rect 3330 3996 3348 4014
rect 3330 4014 3348 4032
rect 3330 4032 3348 4050
rect 3330 4050 3348 4068
rect 3330 4068 3348 4086
rect 3330 4086 3348 4104
rect 3330 4104 3348 4122
rect 3330 4122 3348 4140
rect 3330 4140 3348 4158
rect 3330 4158 3348 4176
rect 3330 4176 3348 4194
rect 3330 4194 3348 4212
rect 3330 4212 3348 4230
rect 3330 4230 3348 4248
rect 3330 4248 3348 4266
rect 3330 4266 3348 4284
rect 3330 4284 3348 4302
rect 3330 4302 3348 4320
rect 3330 4320 3348 4338
rect 3330 4338 3348 4356
rect 3330 4356 3348 4374
rect 3330 4374 3348 4392
rect 3330 4392 3348 4410
rect 3330 6624 3348 6642
rect 3330 6642 3348 6660
rect 3330 6660 3348 6678
rect 3330 6678 3348 6696
rect 3330 6696 3348 6714
rect 3330 6714 3348 6732
rect 3330 6732 3348 6750
rect 3330 6750 3348 6768
rect 3330 6768 3348 6786
rect 3330 6786 3348 6804
rect 3330 6804 3348 6822
rect 3330 6822 3348 6840
rect 3330 6840 3348 6858
rect 3330 6858 3348 6876
rect 3330 6876 3348 6894
rect 3330 6894 3348 6912
rect 3330 6912 3348 6930
rect 3330 6930 3348 6948
rect 3330 6948 3348 6966
rect 3330 6966 3348 6984
rect 3330 6984 3348 7002
rect 3330 7002 3348 7020
rect 3330 7020 3348 7038
rect 3330 7038 3348 7056
rect 3330 7056 3348 7074
rect 3330 7074 3348 7092
rect 3330 7092 3348 7110
rect 3330 7110 3348 7128
rect 3330 7128 3348 7146
rect 3330 7146 3348 7164
rect 3330 7164 3348 7182
rect 3330 7182 3348 7200
rect 3330 7200 3348 7218
rect 3330 7218 3348 7236
rect 3330 7236 3348 7254
rect 3348 36 3366 54
rect 3348 54 3366 72
rect 3348 72 3366 90
rect 3348 90 3366 108
rect 3348 108 3366 126
rect 3348 126 3366 144
rect 3348 144 3366 162
rect 3348 162 3366 180
rect 3348 180 3366 198
rect 3348 198 3366 216
rect 3348 216 3366 234
rect 3348 234 3366 252
rect 3348 252 3366 270
rect 3348 270 3366 288
rect 3348 288 3366 306
rect 3348 306 3366 324
rect 3348 324 3366 342
rect 3348 342 3366 360
rect 3348 360 3366 378
rect 3348 378 3366 396
rect 3348 396 3366 414
rect 3348 414 3366 432
rect 3348 432 3366 450
rect 3348 450 3366 468
rect 3348 468 3366 486
rect 3348 486 3366 504
rect 3348 504 3366 522
rect 3348 522 3366 540
rect 3348 540 3366 558
rect 3348 558 3366 576
rect 3348 576 3366 594
rect 3348 594 3366 612
rect 3348 612 3366 630
rect 3348 756 3366 774
rect 3348 774 3366 792
rect 3348 792 3366 810
rect 3348 810 3366 828
rect 3348 828 3366 846
rect 3348 846 3366 864
rect 3348 864 3366 882
rect 3348 882 3366 900
rect 3348 900 3366 918
rect 3348 918 3366 936
rect 3348 936 3366 954
rect 3348 954 3366 972
rect 3348 972 3366 990
rect 3348 990 3366 1008
rect 3348 1008 3366 1026
rect 3348 1026 3366 1044
rect 3348 1044 3366 1062
rect 3348 1062 3366 1080
rect 3348 1080 3366 1098
rect 3348 1098 3366 1116
rect 3348 1314 3366 1332
rect 3348 1332 3366 1350
rect 3348 1350 3366 1368
rect 3348 1368 3366 1386
rect 3348 1386 3366 1404
rect 3348 1404 3366 1422
rect 3348 1422 3366 1440
rect 3348 1440 3366 1458
rect 3348 1458 3366 1476
rect 3348 1476 3366 1494
rect 3348 1494 3366 1512
rect 3348 1512 3366 1530
rect 3348 1530 3366 1548
rect 3348 1548 3366 1566
rect 3348 1566 3366 1584
rect 3348 1584 3366 1602
rect 3348 1602 3366 1620
rect 3348 1620 3366 1638
rect 3348 1638 3366 1656
rect 3348 1656 3366 1674
rect 3348 1674 3366 1692
rect 3348 1692 3366 1710
rect 3348 1710 3366 1728
rect 3348 1728 3366 1746
rect 3348 1746 3366 1764
rect 3348 1764 3366 1782
rect 3348 1782 3366 1800
rect 3348 1800 3366 1818
rect 3348 1818 3366 1836
rect 3348 1836 3366 1854
rect 3348 1854 3366 1872
rect 3348 1872 3366 1890
rect 3348 1890 3366 1908
rect 3348 1908 3366 1926
rect 3348 1926 3366 1944
rect 3348 1944 3366 1962
rect 3348 1962 3366 1980
rect 3348 1980 3366 1998
rect 3348 1998 3366 2016
rect 3348 2016 3366 2034
rect 3348 2034 3366 2052
rect 3348 2052 3366 2070
rect 3348 2070 3366 2088
rect 3348 2358 3366 2376
rect 3348 2376 3366 2394
rect 3348 2394 3366 2412
rect 3348 2412 3366 2430
rect 3348 2430 3366 2448
rect 3348 2448 3366 2466
rect 3348 2466 3366 2484
rect 3348 2484 3366 2502
rect 3348 2502 3366 2520
rect 3348 2520 3366 2538
rect 3348 2538 3366 2556
rect 3348 2556 3366 2574
rect 3348 2574 3366 2592
rect 3348 2592 3366 2610
rect 3348 2610 3366 2628
rect 3348 2628 3366 2646
rect 3348 2646 3366 2664
rect 3348 2664 3366 2682
rect 3348 2682 3366 2700
rect 3348 2700 3366 2718
rect 3348 2718 3366 2736
rect 3348 2736 3366 2754
rect 3348 2754 3366 2772
rect 3348 2772 3366 2790
rect 3348 2790 3366 2808
rect 3348 2808 3366 2826
rect 3348 2826 3366 2844
rect 3348 2844 3366 2862
rect 3348 2862 3366 2880
rect 3348 2880 3366 2898
rect 3348 2898 3366 2916
rect 3348 2916 3366 2934
rect 3348 2934 3366 2952
rect 3348 2952 3366 2970
rect 3348 2970 3366 2988
rect 3348 2988 3366 3006
rect 3348 3006 3366 3024
rect 3348 3024 3366 3042
rect 3348 3042 3366 3060
rect 3348 3060 3366 3078
rect 3348 3078 3366 3096
rect 3348 3096 3366 3114
rect 3348 3114 3366 3132
rect 3348 3132 3366 3150
rect 3348 3150 3366 3168
rect 3348 3168 3366 3186
rect 3348 3186 3366 3204
rect 3348 3204 3366 3222
rect 3348 3222 3366 3240
rect 3348 3240 3366 3258
rect 3348 3258 3366 3276
rect 3348 3276 3366 3294
rect 3348 3294 3366 3312
rect 3348 3312 3366 3330
rect 3348 3330 3366 3348
rect 3348 3348 3366 3366
rect 3348 3366 3366 3384
rect 3348 3384 3366 3402
rect 3348 3402 3366 3420
rect 3348 3420 3366 3438
rect 3348 3438 3366 3456
rect 3348 3456 3366 3474
rect 3348 3474 3366 3492
rect 3348 3492 3366 3510
rect 3348 3510 3366 3528
rect 3348 3528 3366 3546
rect 3348 3546 3366 3564
rect 3348 3564 3366 3582
rect 3348 3582 3366 3600
rect 3348 3600 3366 3618
rect 3348 3618 3366 3636
rect 3348 3636 3366 3654
rect 3348 3654 3366 3672
rect 3348 3672 3366 3690
rect 3348 3690 3366 3708
rect 3348 3708 3366 3726
rect 3348 3726 3366 3744
rect 3348 3744 3366 3762
rect 3348 3762 3366 3780
rect 3348 3780 3366 3798
rect 3348 3798 3366 3816
rect 3348 3816 3366 3834
rect 3348 3834 3366 3852
rect 3348 3852 3366 3870
rect 3348 3870 3366 3888
rect 3348 3888 3366 3906
rect 3348 3906 3366 3924
rect 3348 3924 3366 3942
rect 3348 3942 3366 3960
rect 3348 3960 3366 3978
rect 3348 3978 3366 3996
rect 3348 3996 3366 4014
rect 3348 4014 3366 4032
rect 3348 4032 3366 4050
rect 3348 4050 3366 4068
rect 3348 4068 3366 4086
rect 3348 4086 3366 4104
rect 3348 4104 3366 4122
rect 3348 4122 3366 4140
rect 3348 4140 3366 4158
rect 3348 4158 3366 4176
rect 3348 4176 3366 4194
rect 3348 4194 3366 4212
rect 3348 4212 3366 4230
rect 3348 4230 3366 4248
rect 3348 4248 3366 4266
rect 3348 4266 3366 4284
rect 3348 4284 3366 4302
rect 3348 4302 3366 4320
rect 3348 4320 3366 4338
rect 3348 4338 3366 4356
rect 3348 4356 3366 4374
rect 3348 4374 3366 4392
rect 3348 4392 3366 4410
rect 3348 4410 3366 4428
rect 3348 4428 3366 4446
rect 3348 4446 3366 4464
rect 3348 6642 3366 6660
rect 3348 6660 3366 6678
rect 3348 6678 3366 6696
rect 3348 6696 3366 6714
rect 3348 6714 3366 6732
rect 3348 6732 3366 6750
rect 3348 6750 3366 6768
rect 3348 6768 3366 6786
rect 3348 6786 3366 6804
rect 3348 6804 3366 6822
rect 3348 6822 3366 6840
rect 3348 6840 3366 6858
rect 3348 6858 3366 6876
rect 3348 6876 3366 6894
rect 3348 6894 3366 6912
rect 3348 6912 3366 6930
rect 3348 6930 3366 6948
rect 3348 6948 3366 6966
rect 3348 6966 3366 6984
rect 3348 6984 3366 7002
rect 3348 7002 3366 7020
rect 3348 7020 3366 7038
rect 3348 7038 3366 7056
rect 3348 7056 3366 7074
rect 3348 7074 3366 7092
rect 3348 7092 3366 7110
rect 3348 7110 3366 7128
rect 3348 7128 3366 7146
rect 3348 7146 3366 7164
rect 3348 7164 3366 7182
rect 3348 7182 3366 7200
rect 3348 7200 3366 7218
rect 3348 7218 3366 7236
rect 3348 7236 3366 7254
rect 3366 36 3384 54
rect 3366 54 3384 72
rect 3366 72 3384 90
rect 3366 90 3384 108
rect 3366 108 3384 126
rect 3366 126 3384 144
rect 3366 144 3384 162
rect 3366 162 3384 180
rect 3366 180 3384 198
rect 3366 198 3384 216
rect 3366 216 3384 234
rect 3366 234 3384 252
rect 3366 252 3384 270
rect 3366 270 3384 288
rect 3366 288 3384 306
rect 3366 306 3384 324
rect 3366 324 3384 342
rect 3366 342 3384 360
rect 3366 360 3384 378
rect 3366 378 3384 396
rect 3366 396 3384 414
rect 3366 414 3384 432
rect 3366 432 3384 450
rect 3366 450 3384 468
rect 3366 468 3384 486
rect 3366 486 3384 504
rect 3366 504 3384 522
rect 3366 522 3384 540
rect 3366 540 3384 558
rect 3366 558 3384 576
rect 3366 576 3384 594
rect 3366 594 3384 612
rect 3366 612 3384 630
rect 3366 774 3384 792
rect 3366 792 3384 810
rect 3366 810 3384 828
rect 3366 828 3384 846
rect 3366 846 3384 864
rect 3366 864 3384 882
rect 3366 882 3384 900
rect 3366 900 3384 918
rect 3366 918 3384 936
rect 3366 936 3384 954
rect 3366 954 3384 972
rect 3366 972 3384 990
rect 3366 990 3384 1008
rect 3366 1008 3384 1026
rect 3366 1026 3384 1044
rect 3366 1044 3384 1062
rect 3366 1062 3384 1080
rect 3366 1080 3384 1098
rect 3366 1098 3384 1116
rect 3366 1116 3384 1134
rect 3366 1332 3384 1350
rect 3366 1350 3384 1368
rect 3366 1368 3384 1386
rect 3366 1386 3384 1404
rect 3366 1404 3384 1422
rect 3366 1422 3384 1440
rect 3366 1440 3384 1458
rect 3366 1458 3384 1476
rect 3366 1476 3384 1494
rect 3366 1494 3384 1512
rect 3366 1512 3384 1530
rect 3366 1530 3384 1548
rect 3366 1548 3384 1566
rect 3366 1566 3384 1584
rect 3366 1584 3384 1602
rect 3366 1602 3384 1620
rect 3366 1620 3384 1638
rect 3366 1638 3384 1656
rect 3366 1656 3384 1674
rect 3366 1674 3384 1692
rect 3366 1692 3384 1710
rect 3366 1710 3384 1728
rect 3366 1728 3384 1746
rect 3366 1746 3384 1764
rect 3366 1764 3384 1782
rect 3366 1782 3384 1800
rect 3366 1800 3384 1818
rect 3366 1818 3384 1836
rect 3366 1836 3384 1854
rect 3366 1854 3384 1872
rect 3366 1872 3384 1890
rect 3366 1890 3384 1908
rect 3366 1908 3384 1926
rect 3366 1926 3384 1944
rect 3366 1944 3384 1962
rect 3366 1962 3384 1980
rect 3366 1980 3384 1998
rect 3366 1998 3384 2016
rect 3366 2016 3384 2034
rect 3366 2034 3384 2052
rect 3366 2052 3384 2070
rect 3366 2070 3384 2088
rect 3366 2088 3384 2106
rect 3366 2394 3384 2412
rect 3366 2412 3384 2430
rect 3366 2430 3384 2448
rect 3366 2448 3384 2466
rect 3366 2466 3384 2484
rect 3366 2484 3384 2502
rect 3366 2502 3384 2520
rect 3366 2520 3384 2538
rect 3366 2538 3384 2556
rect 3366 2556 3384 2574
rect 3366 2574 3384 2592
rect 3366 2592 3384 2610
rect 3366 2610 3384 2628
rect 3366 2628 3384 2646
rect 3366 2646 3384 2664
rect 3366 2664 3384 2682
rect 3366 2682 3384 2700
rect 3366 2700 3384 2718
rect 3366 2718 3384 2736
rect 3366 2736 3384 2754
rect 3366 2754 3384 2772
rect 3366 2772 3384 2790
rect 3366 2790 3384 2808
rect 3366 2808 3384 2826
rect 3366 2826 3384 2844
rect 3366 2844 3384 2862
rect 3366 2862 3384 2880
rect 3366 2880 3384 2898
rect 3366 2898 3384 2916
rect 3366 2916 3384 2934
rect 3366 2934 3384 2952
rect 3366 2952 3384 2970
rect 3366 2970 3384 2988
rect 3366 2988 3384 3006
rect 3366 3006 3384 3024
rect 3366 3024 3384 3042
rect 3366 3042 3384 3060
rect 3366 3060 3384 3078
rect 3366 3078 3384 3096
rect 3366 3096 3384 3114
rect 3366 3114 3384 3132
rect 3366 3132 3384 3150
rect 3366 3150 3384 3168
rect 3366 3168 3384 3186
rect 3366 3186 3384 3204
rect 3366 3204 3384 3222
rect 3366 3222 3384 3240
rect 3366 3240 3384 3258
rect 3366 3258 3384 3276
rect 3366 3276 3384 3294
rect 3366 3294 3384 3312
rect 3366 3312 3384 3330
rect 3366 3330 3384 3348
rect 3366 3348 3384 3366
rect 3366 3366 3384 3384
rect 3366 3384 3384 3402
rect 3366 3402 3384 3420
rect 3366 3420 3384 3438
rect 3366 3438 3384 3456
rect 3366 3456 3384 3474
rect 3366 3474 3384 3492
rect 3366 3492 3384 3510
rect 3366 3510 3384 3528
rect 3366 3528 3384 3546
rect 3366 3546 3384 3564
rect 3366 3564 3384 3582
rect 3366 3582 3384 3600
rect 3366 3600 3384 3618
rect 3366 3618 3384 3636
rect 3366 3636 3384 3654
rect 3366 3654 3384 3672
rect 3366 3672 3384 3690
rect 3366 3690 3384 3708
rect 3366 3708 3384 3726
rect 3366 3726 3384 3744
rect 3366 3744 3384 3762
rect 3366 3762 3384 3780
rect 3366 3780 3384 3798
rect 3366 3798 3384 3816
rect 3366 3816 3384 3834
rect 3366 3834 3384 3852
rect 3366 3852 3384 3870
rect 3366 3870 3384 3888
rect 3366 3888 3384 3906
rect 3366 3906 3384 3924
rect 3366 3924 3384 3942
rect 3366 3942 3384 3960
rect 3366 3960 3384 3978
rect 3366 3978 3384 3996
rect 3366 3996 3384 4014
rect 3366 4014 3384 4032
rect 3366 4032 3384 4050
rect 3366 4050 3384 4068
rect 3366 4068 3384 4086
rect 3366 4086 3384 4104
rect 3366 4104 3384 4122
rect 3366 4122 3384 4140
rect 3366 4140 3384 4158
rect 3366 4158 3384 4176
rect 3366 4176 3384 4194
rect 3366 4194 3384 4212
rect 3366 4212 3384 4230
rect 3366 4230 3384 4248
rect 3366 4248 3384 4266
rect 3366 4266 3384 4284
rect 3366 4284 3384 4302
rect 3366 4302 3384 4320
rect 3366 4320 3384 4338
rect 3366 4338 3384 4356
rect 3366 4356 3384 4374
rect 3366 4374 3384 4392
rect 3366 4392 3384 4410
rect 3366 4410 3384 4428
rect 3366 4428 3384 4446
rect 3366 4446 3384 4464
rect 3366 4464 3384 4482
rect 3366 4482 3384 4500
rect 3366 4500 3384 4518
rect 3366 6642 3384 6660
rect 3366 6660 3384 6678
rect 3366 6678 3384 6696
rect 3366 6696 3384 6714
rect 3366 6714 3384 6732
rect 3366 6732 3384 6750
rect 3366 6750 3384 6768
rect 3366 6768 3384 6786
rect 3366 6786 3384 6804
rect 3366 6804 3384 6822
rect 3366 6822 3384 6840
rect 3366 6840 3384 6858
rect 3366 6858 3384 6876
rect 3366 6876 3384 6894
rect 3366 6894 3384 6912
rect 3366 6912 3384 6930
rect 3366 6930 3384 6948
rect 3366 6948 3384 6966
rect 3366 6966 3384 6984
rect 3366 6984 3384 7002
rect 3366 7002 3384 7020
rect 3366 7020 3384 7038
rect 3366 7038 3384 7056
rect 3366 7056 3384 7074
rect 3366 7074 3384 7092
rect 3366 7092 3384 7110
rect 3366 7110 3384 7128
rect 3366 7128 3384 7146
rect 3366 7146 3384 7164
rect 3366 7164 3384 7182
rect 3366 7182 3384 7200
rect 3366 7200 3384 7218
rect 3366 7218 3384 7236
rect 3366 7236 3384 7254
rect 3384 18 3402 36
rect 3384 36 3402 54
rect 3384 54 3402 72
rect 3384 72 3402 90
rect 3384 90 3402 108
rect 3384 108 3402 126
rect 3384 126 3402 144
rect 3384 144 3402 162
rect 3384 162 3402 180
rect 3384 180 3402 198
rect 3384 198 3402 216
rect 3384 216 3402 234
rect 3384 234 3402 252
rect 3384 252 3402 270
rect 3384 270 3402 288
rect 3384 288 3402 306
rect 3384 306 3402 324
rect 3384 324 3402 342
rect 3384 342 3402 360
rect 3384 360 3402 378
rect 3384 378 3402 396
rect 3384 396 3402 414
rect 3384 414 3402 432
rect 3384 432 3402 450
rect 3384 450 3402 468
rect 3384 468 3402 486
rect 3384 486 3402 504
rect 3384 504 3402 522
rect 3384 522 3402 540
rect 3384 540 3402 558
rect 3384 558 3402 576
rect 3384 576 3402 594
rect 3384 594 3402 612
rect 3384 612 3402 630
rect 3384 774 3402 792
rect 3384 792 3402 810
rect 3384 810 3402 828
rect 3384 828 3402 846
rect 3384 846 3402 864
rect 3384 864 3402 882
rect 3384 882 3402 900
rect 3384 900 3402 918
rect 3384 918 3402 936
rect 3384 936 3402 954
rect 3384 954 3402 972
rect 3384 972 3402 990
rect 3384 990 3402 1008
rect 3384 1008 3402 1026
rect 3384 1026 3402 1044
rect 3384 1044 3402 1062
rect 3384 1062 3402 1080
rect 3384 1080 3402 1098
rect 3384 1098 3402 1116
rect 3384 1116 3402 1134
rect 3384 1332 3402 1350
rect 3384 1350 3402 1368
rect 3384 1368 3402 1386
rect 3384 1386 3402 1404
rect 3384 1404 3402 1422
rect 3384 1422 3402 1440
rect 3384 1440 3402 1458
rect 3384 1458 3402 1476
rect 3384 1476 3402 1494
rect 3384 1494 3402 1512
rect 3384 1512 3402 1530
rect 3384 1530 3402 1548
rect 3384 1548 3402 1566
rect 3384 1566 3402 1584
rect 3384 1584 3402 1602
rect 3384 1602 3402 1620
rect 3384 1620 3402 1638
rect 3384 1638 3402 1656
rect 3384 1656 3402 1674
rect 3384 1674 3402 1692
rect 3384 1692 3402 1710
rect 3384 1710 3402 1728
rect 3384 1728 3402 1746
rect 3384 1746 3402 1764
rect 3384 1764 3402 1782
rect 3384 1782 3402 1800
rect 3384 1800 3402 1818
rect 3384 1818 3402 1836
rect 3384 1836 3402 1854
rect 3384 1854 3402 1872
rect 3384 1872 3402 1890
rect 3384 1890 3402 1908
rect 3384 1908 3402 1926
rect 3384 1926 3402 1944
rect 3384 1944 3402 1962
rect 3384 1962 3402 1980
rect 3384 1980 3402 1998
rect 3384 1998 3402 2016
rect 3384 2016 3402 2034
rect 3384 2034 3402 2052
rect 3384 2052 3402 2070
rect 3384 2070 3402 2088
rect 3384 2088 3402 2106
rect 3384 2106 3402 2124
rect 3384 2124 3402 2142
rect 3384 2430 3402 2448
rect 3384 2448 3402 2466
rect 3384 2466 3402 2484
rect 3384 2484 3402 2502
rect 3384 2502 3402 2520
rect 3384 2520 3402 2538
rect 3384 2538 3402 2556
rect 3384 2556 3402 2574
rect 3384 2574 3402 2592
rect 3384 2592 3402 2610
rect 3384 2610 3402 2628
rect 3384 2628 3402 2646
rect 3384 2646 3402 2664
rect 3384 2664 3402 2682
rect 3384 2682 3402 2700
rect 3384 2700 3402 2718
rect 3384 2718 3402 2736
rect 3384 2736 3402 2754
rect 3384 2754 3402 2772
rect 3384 2772 3402 2790
rect 3384 2790 3402 2808
rect 3384 2808 3402 2826
rect 3384 2826 3402 2844
rect 3384 2844 3402 2862
rect 3384 2862 3402 2880
rect 3384 2880 3402 2898
rect 3384 2898 3402 2916
rect 3384 2916 3402 2934
rect 3384 2934 3402 2952
rect 3384 2952 3402 2970
rect 3384 2970 3402 2988
rect 3384 2988 3402 3006
rect 3384 3006 3402 3024
rect 3384 3024 3402 3042
rect 3384 3042 3402 3060
rect 3384 3060 3402 3078
rect 3384 3078 3402 3096
rect 3384 3096 3402 3114
rect 3384 3114 3402 3132
rect 3384 3132 3402 3150
rect 3384 3150 3402 3168
rect 3384 3168 3402 3186
rect 3384 3186 3402 3204
rect 3384 3204 3402 3222
rect 3384 3222 3402 3240
rect 3384 3240 3402 3258
rect 3384 3258 3402 3276
rect 3384 3276 3402 3294
rect 3384 3294 3402 3312
rect 3384 3312 3402 3330
rect 3384 3330 3402 3348
rect 3384 3348 3402 3366
rect 3384 3366 3402 3384
rect 3384 3384 3402 3402
rect 3384 3402 3402 3420
rect 3384 3420 3402 3438
rect 3384 3438 3402 3456
rect 3384 3456 3402 3474
rect 3384 3474 3402 3492
rect 3384 3492 3402 3510
rect 3384 3510 3402 3528
rect 3384 3528 3402 3546
rect 3384 3546 3402 3564
rect 3384 3564 3402 3582
rect 3384 3582 3402 3600
rect 3384 3600 3402 3618
rect 3384 3618 3402 3636
rect 3384 3636 3402 3654
rect 3384 3654 3402 3672
rect 3384 3672 3402 3690
rect 3384 3690 3402 3708
rect 3384 3708 3402 3726
rect 3384 3726 3402 3744
rect 3384 3744 3402 3762
rect 3384 3762 3402 3780
rect 3384 3780 3402 3798
rect 3384 3798 3402 3816
rect 3384 3816 3402 3834
rect 3384 3834 3402 3852
rect 3384 3852 3402 3870
rect 3384 3870 3402 3888
rect 3384 3888 3402 3906
rect 3384 3906 3402 3924
rect 3384 3924 3402 3942
rect 3384 3942 3402 3960
rect 3384 3960 3402 3978
rect 3384 3978 3402 3996
rect 3384 3996 3402 4014
rect 3384 4014 3402 4032
rect 3384 4032 3402 4050
rect 3384 4050 3402 4068
rect 3384 4068 3402 4086
rect 3384 4086 3402 4104
rect 3384 4104 3402 4122
rect 3384 4122 3402 4140
rect 3384 4140 3402 4158
rect 3384 4158 3402 4176
rect 3384 4176 3402 4194
rect 3384 4194 3402 4212
rect 3384 4212 3402 4230
rect 3384 4230 3402 4248
rect 3384 4248 3402 4266
rect 3384 4266 3402 4284
rect 3384 4284 3402 4302
rect 3384 4302 3402 4320
rect 3384 4320 3402 4338
rect 3384 4338 3402 4356
rect 3384 4356 3402 4374
rect 3384 4374 3402 4392
rect 3384 4392 3402 4410
rect 3384 4410 3402 4428
rect 3384 4428 3402 4446
rect 3384 4446 3402 4464
rect 3384 4464 3402 4482
rect 3384 4482 3402 4500
rect 3384 4500 3402 4518
rect 3384 4518 3402 4536
rect 3384 4536 3402 4554
rect 3384 4554 3402 4572
rect 3384 6642 3402 6660
rect 3384 6660 3402 6678
rect 3384 6678 3402 6696
rect 3384 6696 3402 6714
rect 3384 6714 3402 6732
rect 3384 6732 3402 6750
rect 3384 6750 3402 6768
rect 3384 6768 3402 6786
rect 3384 6786 3402 6804
rect 3384 6804 3402 6822
rect 3384 6822 3402 6840
rect 3384 6840 3402 6858
rect 3384 6858 3402 6876
rect 3384 6876 3402 6894
rect 3384 6894 3402 6912
rect 3384 6912 3402 6930
rect 3384 6930 3402 6948
rect 3384 6948 3402 6966
rect 3384 6966 3402 6984
rect 3384 6984 3402 7002
rect 3384 7002 3402 7020
rect 3384 7020 3402 7038
rect 3384 7038 3402 7056
rect 3384 7056 3402 7074
rect 3384 7074 3402 7092
rect 3384 7092 3402 7110
rect 3384 7110 3402 7128
rect 3384 7128 3402 7146
rect 3384 7146 3402 7164
rect 3384 7164 3402 7182
rect 3384 7182 3402 7200
rect 3384 7200 3402 7218
rect 3384 7218 3402 7236
rect 3384 7236 3402 7254
rect 3384 7254 3402 7272
rect 3402 18 3420 36
rect 3402 36 3420 54
rect 3402 54 3420 72
rect 3402 72 3420 90
rect 3402 90 3420 108
rect 3402 108 3420 126
rect 3402 126 3420 144
rect 3402 144 3420 162
rect 3402 162 3420 180
rect 3402 180 3420 198
rect 3402 198 3420 216
rect 3402 216 3420 234
rect 3402 234 3420 252
rect 3402 252 3420 270
rect 3402 270 3420 288
rect 3402 288 3420 306
rect 3402 306 3420 324
rect 3402 324 3420 342
rect 3402 342 3420 360
rect 3402 360 3420 378
rect 3402 378 3420 396
rect 3402 396 3420 414
rect 3402 414 3420 432
rect 3402 432 3420 450
rect 3402 450 3420 468
rect 3402 468 3420 486
rect 3402 486 3420 504
rect 3402 504 3420 522
rect 3402 522 3420 540
rect 3402 540 3420 558
rect 3402 558 3420 576
rect 3402 576 3420 594
rect 3402 594 3420 612
rect 3402 612 3420 630
rect 3402 774 3420 792
rect 3402 792 3420 810
rect 3402 810 3420 828
rect 3402 828 3420 846
rect 3402 846 3420 864
rect 3402 864 3420 882
rect 3402 882 3420 900
rect 3402 900 3420 918
rect 3402 918 3420 936
rect 3402 936 3420 954
rect 3402 954 3420 972
rect 3402 972 3420 990
rect 3402 990 3420 1008
rect 3402 1008 3420 1026
rect 3402 1026 3420 1044
rect 3402 1044 3420 1062
rect 3402 1062 3420 1080
rect 3402 1080 3420 1098
rect 3402 1098 3420 1116
rect 3402 1116 3420 1134
rect 3402 1134 3420 1152
rect 3402 1350 3420 1368
rect 3402 1368 3420 1386
rect 3402 1386 3420 1404
rect 3402 1404 3420 1422
rect 3402 1422 3420 1440
rect 3402 1440 3420 1458
rect 3402 1458 3420 1476
rect 3402 1476 3420 1494
rect 3402 1494 3420 1512
rect 3402 1512 3420 1530
rect 3402 1530 3420 1548
rect 3402 1548 3420 1566
rect 3402 1566 3420 1584
rect 3402 1584 3420 1602
rect 3402 1602 3420 1620
rect 3402 1620 3420 1638
rect 3402 1638 3420 1656
rect 3402 1656 3420 1674
rect 3402 1674 3420 1692
rect 3402 1692 3420 1710
rect 3402 1710 3420 1728
rect 3402 1728 3420 1746
rect 3402 1746 3420 1764
rect 3402 1764 3420 1782
rect 3402 1782 3420 1800
rect 3402 1800 3420 1818
rect 3402 1818 3420 1836
rect 3402 1836 3420 1854
rect 3402 1854 3420 1872
rect 3402 1872 3420 1890
rect 3402 1890 3420 1908
rect 3402 1908 3420 1926
rect 3402 1926 3420 1944
rect 3402 1944 3420 1962
rect 3402 1962 3420 1980
rect 3402 1980 3420 1998
rect 3402 1998 3420 2016
rect 3402 2016 3420 2034
rect 3402 2034 3420 2052
rect 3402 2052 3420 2070
rect 3402 2070 3420 2088
rect 3402 2088 3420 2106
rect 3402 2106 3420 2124
rect 3402 2124 3420 2142
rect 3402 2142 3420 2160
rect 3402 2160 3420 2178
rect 3402 2448 3420 2466
rect 3402 2466 3420 2484
rect 3402 2484 3420 2502
rect 3402 2502 3420 2520
rect 3402 2520 3420 2538
rect 3402 2538 3420 2556
rect 3402 2556 3420 2574
rect 3402 2574 3420 2592
rect 3402 2592 3420 2610
rect 3402 2610 3420 2628
rect 3402 2628 3420 2646
rect 3402 2646 3420 2664
rect 3402 2664 3420 2682
rect 3402 2682 3420 2700
rect 3402 2700 3420 2718
rect 3402 2718 3420 2736
rect 3402 2736 3420 2754
rect 3402 2754 3420 2772
rect 3402 2772 3420 2790
rect 3402 2790 3420 2808
rect 3402 2808 3420 2826
rect 3402 2826 3420 2844
rect 3402 2844 3420 2862
rect 3402 2862 3420 2880
rect 3402 2880 3420 2898
rect 3402 2898 3420 2916
rect 3402 2916 3420 2934
rect 3402 2934 3420 2952
rect 3402 2952 3420 2970
rect 3402 2970 3420 2988
rect 3402 2988 3420 3006
rect 3402 3006 3420 3024
rect 3402 3024 3420 3042
rect 3402 3042 3420 3060
rect 3402 3060 3420 3078
rect 3402 3078 3420 3096
rect 3402 3096 3420 3114
rect 3402 3114 3420 3132
rect 3402 3132 3420 3150
rect 3402 3150 3420 3168
rect 3402 3168 3420 3186
rect 3402 3186 3420 3204
rect 3402 3204 3420 3222
rect 3402 3222 3420 3240
rect 3402 3240 3420 3258
rect 3402 3258 3420 3276
rect 3402 3276 3420 3294
rect 3402 3294 3420 3312
rect 3402 3312 3420 3330
rect 3402 3330 3420 3348
rect 3402 3348 3420 3366
rect 3402 3366 3420 3384
rect 3402 3384 3420 3402
rect 3402 3402 3420 3420
rect 3402 3420 3420 3438
rect 3402 3438 3420 3456
rect 3402 3456 3420 3474
rect 3402 3474 3420 3492
rect 3402 3492 3420 3510
rect 3402 3510 3420 3528
rect 3402 3528 3420 3546
rect 3402 3546 3420 3564
rect 3402 3564 3420 3582
rect 3402 3582 3420 3600
rect 3402 3600 3420 3618
rect 3402 3618 3420 3636
rect 3402 3636 3420 3654
rect 3402 3654 3420 3672
rect 3402 3672 3420 3690
rect 3402 3690 3420 3708
rect 3402 3708 3420 3726
rect 3402 3726 3420 3744
rect 3402 3744 3420 3762
rect 3402 3762 3420 3780
rect 3402 3780 3420 3798
rect 3402 3798 3420 3816
rect 3402 3816 3420 3834
rect 3402 3834 3420 3852
rect 3402 3852 3420 3870
rect 3402 3870 3420 3888
rect 3402 3888 3420 3906
rect 3402 3906 3420 3924
rect 3402 3924 3420 3942
rect 3402 3942 3420 3960
rect 3402 3960 3420 3978
rect 3402 3978 3420 3996
rect 3402 3996 3420 4014
rect 3402 4014 3420 4032
rect 3402 4032 3420 4050
rect 3402 4050 3420 4068
rect 3402 4068 3420 4086
rect 3402 4086 3420 4104
rect 3402 4104 3420 4122
rect 3402 4122 3420 4140
rect 3402 4140 3420 4158
rect 3402 4158 3420 4176
rect 3402 4176 3420 4194
rect 3402 4194 3420 4212
rect 3402 4212 3420 4230
rect 3402 4230 3420 4248
rect 3402 4248 3420 4266
rect 3402 4266 3420 4284
rect 3402 4284 3420 4302
rect 3402 4302 3420 4320
rect 3402 4320 3420 4338
rect 3402 4338 3420 4356
rect 3402 4356 3420 4374
rect 3402 4374 3420 4392
rect 3402 4392 3420 4410
rect 3402 4410 3420 4428
rect 3402 4428 3420 4446
rect 3402 4446 3420 4464
rect 3402 4464 3420 4482
rect 3402 4482 3420 4500
rect 3402 4500 3420 4518
rect 3402 4518 3420 4536
rect 3402 4536 3420 4554
rect 3402 4554 3420 4572
rect 3402 4572 3420 4590
rect 3402 4590 3420 4608
rect 3402 4608 3420 4626
rect 3402 6642 3420 6660
rect 3402 6660 3420 6678
rect 3402 6678 3420 6696
rect 3402 6696 3420 6714
rect 3402 6714 3420 6732
rect 3402 6732 3420 6750
rect 3402 6750 3420 6768
rect 3402 6768 3420 6786
rect 3402 6786 3420 6804
rect 3402 6804 3420 6822
rect 3402 6822 3420 6840
rect 3402 6840 3420 6858
rect 3402 6858 3420 6876
rect 3402 6876 3420 6894
rect 3402 6894 3420 6912
rect 3402 6912 3420 6930
rect 3402 6930 3420 6948
rect 3402 6948 3420 6966
rect 3402 6966 3420 6984
rect 3402 6984 3420 7002
rect 3402 7002 3420 7020
rect 3402 7020 3420 7038
rect 3402 7038 3420 7056
rect 3402 7056 3420 7074
rect 3402 7074 3420 7092
rect 3402 7092 3420 7110
rect 3402 7110 3420 7128
rect 3402 7128 3420 7146
rect 3402 7146 3420 7164
rect 3402 7164 3420 7182
rect 3402 7182 3420 7200
rect 3402 7200 3420 7218
rect 3402 7218 3420 7236
rect 3402 7236 3420 7254
rect 3402 7254 3420 7272
rect 3420 18 3438 36
rect 3420 36 3438 54
rect 3420 54 3438 72
rect 3420 72 3438 90
rect 3420 90 3438 108
rect 3420 108 3438 126
rect 3420 126 3438 144
rect 3420 144 3438 162
rect 3420 162 3438 180
rect 3420 180 3438 198
rect 3420 198 3438 216
rect 3420 216 3438 234
rect 3420 234 3438 252
rect 3420 252 3438 270
rect 3420 270 3438 288
rect 3420 288 3438 306
rect 3420 306 3438 324
rect 3420 324 3438 342
rect 3420 342 3438 360
rect 3420 360 3438 378
rect 3420 378 3438 396
rect 3420 396 3438 414
rect 3420 414 3438 432
rect 3420 432 3438 450
rect 3420 450 3438 468
rect 3420 468 3438 486
rect 3420 486 3438 504
rect 3420 504 3438 522
rect 3420 522 3438 540
rect 3420 540 3438 558
rect 3420 558 3438 576
rect 3420 576 3438 594
rect 3420 594 3438 612
rect 3420 612 3438 630
rect 3420 792 3438 810
rect 3420 810 3438 828
rect 3420 828 3438 846
rect 3420 846 3438 864
rect 3420 864 3438 882
rect 3420 882 3438 900
rect 3420 900 3438 918
rect 3420 918 3438 936
rect 3420 936 3438 954
rect 3420 954 3438 972
rect 3420 972 3438 990
rect 3420 990 3438 1008
rect 3420 1008 3438 1026
rect 3420 1026 3438 1044
rect 3420 1044 3438 1062
rect 3420 1062 3438 1080
rect 3420 1080 3438 1098
rect 3420 1098 3438 1116
rect 3420 1116 3438 1134
rect 3420 1134 3438 1152
rect 3420 1152 3438 1170
rect 3420 1368 3438 1386
rect 3420 1386 3438 1404
rect 3420 1404 3438 1422
rect 3420 1422 3438 1440
rect 3420 1440 3438 1458
rect 3420 1458 3438 1476
rect 3420 1476 3438 1494
rect 3420 1494 3438 1512
rect 3420 1512 3438 1530
rect 3420 1530 3438 1548
rect 3420 1548 3438 1566
rect 3420 1566 3438 1584
rect 3420 1584 3438 1602
rect 3420 1602 3438 1620
rect 3420 1620 3438 1638
rect 3420 1638 3438 1656
rect 3420 1656 3438 1674
rect 3420 1674 3438 1692
rect 3420 1692 3438 1710
rect 3420 1710 3438 1728
rect 3420 1728 3438 1746
rect 3420 1746 3438 1764
rect 3420 1764 3438 1782
rect 3420 1782 3438 1800
rect 3420 1800 3438 1818
rect 3420 1818 3438 1836
rect 3420 1836 3438 1854
rect 3420 1854 3438 1872
rect 3420 1872 3438 1890
rect 3420 1890 3438 1908
rect 3420 1908 3438 1926
rect 3420 1926 3438 1944
rect 3420 1944 3438 1962
rect 3420 1962 3438 1980
rect 3420 1980 3438 1998
rect 3420 1998 3438 2016
rect 3420 2016 3438 2034
rect 3420 2034 3438 2052
rect 3420 2052 3438 2070
rect 3420 2070 3438 2088
rect 3420 2088 3438 2106
rect 3420 2106 3438 2124
rect 3420 2124 3438 2142
rect 3420 2142 3438 2160
rect 3420 2160 3438 2178
rect 3420 2178 3438 2196
rect 3420 2484 3438 2502
rect 3420 2502 3438 2520
rect 3420 2520 3438 2538
rect 3420 2538 3438 2556
rect 3420 2556 3438 2574
rect 3420 2574 3438 2592
rect 3420 2592 3438 2610
rect 3420 2610 3438 2628
rect 3420 2628 3438 2646
rect 3420 2646 3438 2664
rect 3420 2664 3438 2682
rect 3420 2682 3438 2700
rect 3420 2700 3438 2718
rect 3420 2718 3438 2736
rect 3420 2736 3438 2754
rect 3420 2754 3438 2772
rect 3420 2772 3438 2790
rect 3420 2790 3438 2808
rect 3420 2808 3438 2826
rect 3420 2826 3438 2844
rect 3420 2844 3438 2862
rect 3420 2862 3438 2880
rect 3420 2880 3438 2898
rect 3420 2898 3438 2916
rect 3420 2916 3438 2934
rect 3420 2934 3438 2952
rect 3420 2952 3438 2970
rect 3420 2970 3438 2988
rect 3420 2988 3438 3006
rect 3420 3006 3438 3024
rect 3420 3024 3438 3042
rect 3420 3042 3438 3060
rect 3420 3060 3438 3078
rect 3420 3078 3438 3096
rect 3420 3096 3438 3114
rect 3420 3114 3438 3132
rect 3420 3132 3438 3150
rect 3420 3150 3438 3168
rect 3420 3168 3438 3186
rect 3420 3186 3438 3204
rect 3420 3204 3438 3222
rect 3420 3222 3438 3240
rect 3420 3240 3438 3258
rect 3420 3258 3438 3276
rect 3420 3276 3438 3294
rect 3420 3294 3438 3312
rect 3420 3312 3438 3330
rect 3420 3330 3438 3348
rect 3420 3348 3438 3366
rect 3420 3366 3438 3384
rect 3420 3384 3438 3402
rect 3420 3402 3438 3420
rect 3420 3420 3438 3438
rect 3420 3438 3438 3456
rect 3420 3456 3438 3474
rect 3420 3474 3438 3492
rect 3420 3492 3438 3510
rect 3420 3510 3438 3528
rect 3420 3528 3438 3546
rect 3420 3546 3438 3564
rect 3420 3564 3438 3582
rect 3420 3582 3438 3600
rect 3420 3600 3438 3618
rect 3420 3618 3438 3636
rect 3420 3636 3438 3654
rect 3420 3654 3438 3672
rect 3420 3672 3438 3690
rect 3420 3690 3438 3708
rect 3420 3708 3438 3726
rect 3420 3726 3438 3744
rect 3420 3744 3438 3762
rect 3420 3762 3438 3780
rect 3420 3780 3438 3798
rect 3420 3798 3438 3816
rect 3420 3816 3438 3834
rect 3420 3834 3438 3852
rect 3420 3852 3438 3870
rect 3420 3870 3438 3888
rect 3420 3888 3438 3906
rect 3420 3906 3438 3924
rect 3420 3924 3438 3942
rect 3420 3942 3438 3960
rect 3420 3960 3438 3978
rect 3420 3978 3438 3996
rect 3420 3996 3438 4014
rect 3420 4014 3438 4032
rect 3420 4032 3438 4050
rect 3420 4050 3438 4068
rect 3420 4068 3438 4086
rect 3420 4086 3438 4104
rect 3420 4104 3438 4122
rect 3420 4122 3438 4140
rect 3420 4140 3438 4158
rect 3420 4158 3438 4176
rect 3420 4176 3438 4194
rect 3420 4194 3438 4212
rect 3420 4212 3438 4230
rect 3420 4230 3438 4248
rect 3420 4248 3438 4266
rect 3420 4266 3438 4284
rect 3420 4284 3438 4302
rect 3420 4302 3438 4320
rect 3420 4320 3438 4338
rect 3420 4338 3438 4356
rect 3420 4356 3438 4374
rect 3420 4374 3438 4392
rect 3420 4392 3438 4410
rect 3420 4410 3438 4428
rect 3420 4428 3438 4446
rect 3420 4446 3438 4464
rect 3420 4464 3438 4482
rect 3420 4482 3438 4500
rect 3420 4500 3438 4518
rect 3420 4518 3438 4536
rect 3420 4536 3438 4554
rect 3420 4554 3438 4572
rect 3420 4572 3438 4590
rect 3420 4590 3438 4608
rect 3420 4608 3438 4626
rect 3420 4626 3438 4644
rect 3420 4644 3438 4662
rect 3420 6642 3438 6660
rect 3420 6660 3438 6678
rect 3420 6678 3438 6696
rect 3420 6696 3438 6714
rect 3420 6714 3438 6732
rect 3420 6732 3438 6750
rect 3420 6750 3438 6768
rect 3420 6768 3438 6786
rect 3420 6786 3438 6804
rect 3420 6804 3438 6822
rect 3420 6822 3438 6840
rect 3420 6840 3438 6858
rect 3420 6858 3438 6876
rect 3420 6876 3438 6894
rect 3420 6894 3438 6912
rect 3420 6912 3438 6930
rect 3420 6930 3438 6948
rect 3420 6948 3438 6966
rect 3420 6966 3438 6984
rect 3420 6984 3438 7002
rect 3420 7002 3438 7020
rect 3420 7020 3438 7038
rect 3420 7038 3438 7056
rect 3420 7056 3438 7074
rect 3420 7074 3438 7092
rect 3420 7092 3438 7110
rect 3420 7110 3438 7128
rect 3420 7128 3438 7146
rect 3420 7146 3438 7164
rect 3420 7164 3438 7182
rect 3420 7182 3438 7200
rect 3420 7200 3438 7218
rect 3420 7218 3438 7236
rect 3420 7236 3438 7254
rect 3420 7254 3438 7272
rect 3438 18 3456 36
rect 3438 36 3456 54
rect 3438 54 3456 72
rect 3438 72 3456 90
rect 3438 90 3456 108
rect 3438 108 3456 126
rect 3438 126 3456 144
rect 3438 144 3456 162
rect 3438 162 3456 180
rect 3438 180 3456 198
rect 3438 198 3456 216
rect 3438 216 3456 234
rect 3438 234 3456 252
rect 3438 252 3456 270
rect 3438 270 3456 288
rect 3438 288 3456 306
rect 3438 306 3456 324
rect 3438 324 3456 342
rect 3438 342 3456 360
rect 3438 360 3456 378
rect 3438 378 3456 396
rect 3438 396 3456 414
rect 3438 414 3456 432
rect 3438 432 3456 450
rect 3438 450 3456 468
rect 3438 468 3456 486
rect 3438 486 3456 504
rect 3438 504 3456 522
rect 3438 522 3456 540
rect 3438 540 3456 558
rect 3438 558 3456 576
rect 3438 576 3456 594
rect 3438 594 3456 612
rect 3438 612 3456 630
rect 3438 792 3456 810
rect 3438 810 3456 828
rect 3438 828 3456 846
rect 3438 846 3456 864
rect 3438 864 3456 882
rect 3438 882 3456 900
rect 3438 900 3456 918
rect 3438 918 3456 936
rect 3438 936 3456 954
rect 3438 954 3456 972
rect 3438 972 3456 990
rect 3438 990 3456 1008
rect 3438 1008 3456 1026
rect 3438 1026 3456 1044
rect 3438 1044 3456 1062
rect 3438 1062 3456 1080
rect 3438 1080 3456 1098
rect 3438 1098 3456 1116
rect 3438 1116 3456 1134
rect 3438 1134 3456 1152
rect 3438 1152 3456 1170
rect 3438 1170 3456 1188
rect 3438 1386 3456 1404
rect 3438 1404 3456 1422
rect 3438 1422 3456 1440
rect 3438 1440 3456 1458
rect 3438 1458 3456 1476
rect 3438 1476 3456 1494
rect 3438 1494 3456 1512
rect 3438 1512 3456 1530
rect 3438 1530 3456 1548
rect 3438 1548 3456 1566
rect 3438 1566 3456 1584
rect 3438 1584 3456 1602
rect 3438 1602 3456 1620
rect 3438 1620 3456 1638
rect 3438 1638 3456 1656
rect 3438 1656 3456 1674
rect 3438 1674 3456 1692
rect 3438 1692 3456 1710
rect 3438 1710 3456 1728
rect 3438 1728 3456 1746
rect 3438 1746 3456 1764
rect 3438 1764 3456 1782
rect 3438 1782 3456 1800
rect 3438 1800 3456 1818
rect 3438 1818 3456 1836
rect 3438 1836 3456 1854
rect 3438 1854 3456 1872
rect 3438 1872 3456 1890
rect 3438 1890 3456 1908
rect 3438 1908 3456 1926
rect 3438 1926 3456 1944
rect 3438 1944 3456 1962
rect 3438 1962 3456 1980
rect 3438 1980 3456 1998
rect 3438 1998 3456 2016
rect 3438 2016 3456 2034
rect 3438 2034 3456 2052
rect 3438 2052 3456 2070
rect 3438 2070 3456 2088
rect 3438 2088 3456 2106
rect 3438 2106 3456 2124
rect 3438 2124 3456 2142
rect 3438 2142 3456 2160
rect 3438 2160 3456 2178
rect 3438 2178 3456 2196
rect 3438 2196 3456 2214
rect 3438 2214 3456 2232
rect 3438 2502 3456 2520
rect 3438 2520 3456 2538
rect 3438 2538 3456 2556
rect 3438 2556 3456 2574
rect 3438 2574 3456 2592
rect 3438 2592 3456 2610
rect 3438 2610 3456 2628
rect 3438 2628 3456 2646
rect 3438 2646 3456 2664
rect 3438 2664 3456 2682
rect 3438 2682 3456 2700
rect 3438 2700 3456 2718
rect 3438 2718 3456 2736
rect 3438 2736 3456 2754
rect 3438 2754 3456 2772
rect 3438 2772 3456 2790
rect 3438 2790 3456 2808
rect 3438 2808 3456 2826
rect 3438 2826 3456 2844
rect 3438 2844 3456 2862
rect 3438 2862 3456 2880
rect 3438 2880 3456 2898
rect 3438 2898 3456 2916
rect 3438 2916 3456 2934
rect 3438 2934 3456 2952
rect 3438 2952 3456 2970
rect 3438 2970 3456 2988
rect 3438 2988 3456 3006
rect 3438 3006 3456 3024
rect 3438 3024 3456 3042
rect 3438 3042 3456 3060
rect 3438 3060 3456 3078
rect 3438 3078 3456 3096
rect 3438 3096 3456 3114
rect 3438 3114 3456 3132
rect 3438 3132 3456 3150
rect 3438 3150 3456 3168
rect 3438 3168 3456 3186
rect 3438 3186 3456 3204
rect 3438 3204 3456 3222
rect 3438 3222 3456 3240
rect 3438 3240 3456 3258
rect 3438 3258 3456 3276
rect 3438 3276 3456 3294
rect 3438 3294 3456 3312
rect 3438 3312 3456 3330
rect 3438 3330 3456 3348
rect 3438 3348 3456 3366
rect 3438 3366 3456 3384
rect 3438 3384 3456 3402
rect 3438 3402 3456 3420
rect 3438 3420 3456 3438
rect 3438 3438 3456 3456
rect 3438 3456 3456 3474
rect 3438 3474 3456 3492
rect 3438 3492 3456 3510
rect 3438 3510 3456 3528
rect 3438 3528 3456 3546
rect 3438 3546 3456 3564
rect 3438 3564 3456 3582
rect 3438 3582 3456 3600
rect 3438 3600 3456 3618
rect 3438 3618 3456 3636
rect 3438 3636 3456 3654
rect 3438 3654 3456 3672
rect 3438 3672 3456 3690
rect 3438 3690 3456 3708
rect 3438 3708 3456 3726
rect 3438 3726 3456 3744
rect 3438 3744 3456 3762
rect 3438 3762 3456 3780
rect 3438 3780 3456 3798
rect 3438 3798 3456 3816
rect 3438 3816 3456 3834
rect 3438 3834 3456 3852
rect 3438 3852 3456 3870
rect 3438 3870 3456 3888
rect 3438 3888 3456 3906
rect 3438 3906 3456 3924
rect 3438 3924 3456 3942
rect 3438 3942 3456 3960
rect 3438 3960 3456 3978
rect 3438 3978 3456 3996
rect 3438 3996 3456 4014
rect 3438 4014 3456 4032
rect 3438 4032 3456 4050
rect 3438 4050 3456 4068
rect 3438 4068 3456 4086
rect 3438 4086 3456 4104
rect 3438 4104 3456 4122
rect 3438 4122 3456 4140
rect 3438 4140 3456 4158
rect 3438 4158 3456 4176
rect 3438 4176 3456 4194
rect 3438 4194 3456 4212
rect 3438 4212 3456 4230
rect 3438 4230 3456 4248
rect 3438 4248 3456 4266
rect 3438 4266 3456 4284
rect 3438 4284 3456 4302
rect 3438 4302 3456 4320
rect 3438 4320 3456 4338
rect 3438 4338 3456 4356
rect 3438 4356 3456 4374
rect 3438 4374 3456 4392
rect 3438 4392 3456 4410
rect 3438 4410 3456 4428
rect 3438 4428 3456 4446
rect 3438 4446 3456 4464
rect 3438 4464 3456 4482
rect 3438 4482 3456 4500
rect 3438 4500 3456 4518
rect 3438 4518 3456 4536
rect 3438 4536 3456 4554
rect 3438 4554 3456 4572
rect 3438 4572 3456 4590
rect 3438 4590 3456 4608
rect 3438 4608 3456 4626
rect 3438 4626 3456 4644
rect 3438 4644 3456 4662
rect 3438 4662 3456 4680
rect 3438 4680 3456 4698
rect 3438 4698 3456 4716
rect 3438 6642 3456 6660
rect 3438 6660 3456 6678
rect 3438 6678 3456 6696
rect 3438 6696 3456 6714
rect 3438 6714 3456 6732
rect 3438 6732 3456 6750
rect 3438 6750 3456 6768
rect 3438 6768 3456 6786
rect 3438 6786 3456 6804
rect 3438 6804 3456 6822
rect 3438 6822 3456 6840
rect 3438 6840 3456 6858
rect 3438 6858 3456 6876
rect 3438 6876 3456 6894
rect 3438 6894 3456 6912
rect 3438 6912 3456 6930
rect 3438 6930 3456 6948
rect 3438 6948 3456 6966
rect 3438 6966 3456 6984
rect 3438 6984 3456 7002
rect 3438 7002 3456 7020
rect 3438 7020 3456 7038
rect 3438 7038 3456 7056
rect 3438 7056 3456 7074
rect 3438 7074 3456 7092
rect 3438 7092 3456 7110
rect 3438 7110 3456 7128
rect 3438 7128 3456 7146
rect 3438 7146 3456 7164
rect 3438 7164 3456 7182
rect 3438 7182 3456 7200
rect 3438 7200 3456 7218
rect 3438 7218 3456 7236
rect 3438 7236 3456 7254
rect 3438 7254 3456 7272
rect 3456 18 3474 36
rect 3456 36 3474 54
rect 3456 54 3474 72
rect 3456 72 3474 90
rect 3456 90 3474 108
rect 3456 108 3474 126
rect 3456 126 3474 144
rect 3456 144 3474 162
rect 3456 162 3474 180
rect 3456 180 3474 198
rect 3456 198 3474 216
rect 3456 216 3474 234
rect 3456 234 3474 252
rect 3456 252 3474 270
rect 3456 270 3474 288
rect 3456 288 3474 306
rect 3456 306 3474 324
rect 3456 324 3474 342
rect 3456 342 3474 360
rect 3456 360 3474 378
rect 3456 378 3474 396
rect 3456 396 3474 414
rect 3456 414 3474 432
rect 3456 432 3474 450
rect 3456 450 3474 468
rect 3456 468 3474 486
rect 3456 486 3474 504
rect 3456 504 3474 522
rect 3456 522 3474 540
rect 3456 540 3474 558
rect 3456 558 3474 576
rect 3456 576 3474 594
rect 3456 594 3474 612
rect 3456 612 3474 630
rect 3456 810 3474 828
rect 3456 828 3474 846
rect 3456 846 3474 864
rect 3456 864 3474 882
rect 3456 882 3474 900
rect 3456 900 3474 918
rect 3456 918 3474 936
rect 3456 936 3474 954
rect 3456 954 3474 972
rect 3456 972 3474 990
rect 3456 990 3474 1008
rect 3456 1008 3474 1026
rect 3456 1026 3474 1044
rect 3456 1044 3474 1062
rect 3456 1062 3474 1080
rect 3456 1080 3474 1098
rect 3456 1098 3474 1116
rect 3456 1116 3474 1134
rect 3456 1134 3474 1152
rect 3456 1152 3474 1170
rect 3456 1170 3474 1188
rect 3456 1404 3474 1422
rect 3456 1422 3474 1440
rect 3456 1440 3474 1458
rect 3456 1458 3474 1476
rect 3456 1476 3474 1494
rect 3456 1494 3474 1512
rect 3456 1512 3474 1530
rect 3456 1530 3474 1548
rect 3456 1548 3474 1566
rect 3456 1566 3474 1584
rect 3456 1584 3474 1602
rect 3456 1602 3474 1620
rect 3456 1620 3474 1638
rect 3456 1638 3474 1656
rect 3456 1656 3474 1674
rect 3456 1674 3474 1692
rect 3456 1692 3474 1710
rect 3456 1710 3474 1728
rect 3456 1728 3474 1746
rect 3456 1746 3474 1764
rect 3456 1764 3474 1782
rect 3456 1782 3474 1800
rect 3456 1800 3474 1818
rect 3456 1818 3474 1836
rect 3456 1836 3474 1854
rect 3456 1854 3474 1872
rect 3456 1872 3474 1890
rect 3456 1890 3474 1908
rect 3456 1908 3474 1926
rect 3456 1926 3474 1944
rect 3456 1944 3474 1962
rect 3456 1962 3474 1980
rect 3456 1980 3474 1998
rect 3456 1998 3474 2016
rect 3456 2016 3474 2034
rect 3456 2034 3474 2052
rect 3456 2052 3474 2070
rect 3456 2070 3474 2088
rect 3456 2088 3474 2106
rect 3456 2106 3474 2124
rect 3456 2124 3474 2142
rect 3456 2142 3474 2160
rect 3456 2160 3474 2178
rect 3456 2178 3474 2196
rect 3456 2196 3474 2214
rect 3456 2214 3474 2232
rect 3456 2232 3474 2250
rect 3456 2250 3474 2268
rect 3456 2538 3474 2556
rect 3456 2556 3474 2574
rect 3456 2574 3474 2592
rect 3456 2592 3474 2610
rect 3456 2610 3474 2628
rect 3456 2628 3474 2646
rect 3456 2646 3474 2664
rect 3456 2664 3474 2682
rect 3456 2682 3474 2700
rect 3456 2700 3474 2718
rect 3456 2718 3474 2736
rect 3456 2736 3474 2754
rect 3456 2754 3474 2772
rect 3456 2772 3474 2790
rect 3456 2790 3474 2808
rect 3456 2808 3474 2826
rect 3456 2826 3474 2844
rect 3456 2844 3474 2862
rect 3456 2862 3474 2880
rect 3456 2880 3474 2898
rect 3456 2898 3474 2916
rect 3456 2916 3474 2934
rect 3456 2934 3474 2952
rect 3456 2952 3474 2970
rect 3456 2970 3474 2988
rect 3456 2988 3474 3006
rect 3456 3006 3474 3024
rect 3456 3024 3474 3042
rect 3456 3042 3474 3060
rect 3456 3060 3474 3078
rect 3456 3078 3474 3096
rect 3456 3096 3474 3114
rect 3456 3114 3474 3132
rect 3456 3132 3474 3150
rect 3456 3150 3474 3168
rect 3456 3168 3474 3186
rect 3456 3186 3474 3204
rect 3456 3204 3474 3222
rect 3456 3222 3474 3240
rect 3456 3240 3474 3258
rect 3456 3258 3474 3276
rect 3456 3276 3474 3294
rect 3456 3294 3474 3312
rect 3456 3312 3474 3330
rect 3456 3330 3474 3348
rect 3456 3348 3474 3366
rect 3456 3366 3474 3384
rect 3456 3384 3474 3402
rect 3456 3402 3474 3420
rect 3456 3420 3474 3438
rect 3456 3438 3474 3456
rect 3456 3456 3474 3474
rect 3456 3474 3474 3492
rect 3456 3492 3474 3510
rect 3456 3510 3474 3528
rect 3456 3528 3474 3546
rect 3456 3546 3474 3564
rect 3456 3564 3474 3582
rect 3456 3582 3474 3600
rect 3456 3600 3474 3618
rect 3456 3618 3474 3636
rect 3456 3636 3474 3654
rect 3456 3654 3474 3672
rect 3456 3672 3474 3690
rect 3456 3690 3474 3708
rect 3456 3708 3474 3726
rect 3456 3726 3474 3744
rect 3456 3744 3474 3762
rect 3456 3762 3474 3780
rect 3456 3780 3474 3798
rect 3456 3798 3474 3816
rect 3456 3816 3474 3834
rect 3456 3834 3474 3852
rect 3456 3852 3474 3870
rect 3456 3870 3474 3888
rect 3456 3888 3474 3906
rect 3456 3906 3474 3924
rect 3456 3924 3474 3942
rect 3456 3942 3474 3960
rect 3456 3960 3474 3978
rect 3456 3978 3474 3996
rect 3456 3996 3474 4014
rect 3456 4014 3474 4032
rect 3456 4032 3474 4050
rect 3456 4050 3474 4068
rect 3456 4068 3474 4086
rect 3456 4086 3474 4104
rect 3456 4104 3474 4122
rect 3456 4122 3474 4140
rect 3456 4140 3474 4158
rect 3456 4158 3474 4176
rect 3456 4176 3474 4194
rect 3456 4194 3474 4212
rect 3456 4212 3474 4230
rect 3456 4230 3474 4248
rect 3456 4248 3474 4266
rect 3456 4266 3474 4284
rect 3456 4284 3474 4302
rect 3456 4302 3474 4320
rect 3456 4320 3474 4338
rect 3456 4338 3474 4356
rect 3456 4356 3474 4374
rect 3456 4374 3474 4392
rect 3456 4392 3474 4410
rect 3456 4410 3474 4428
rect 3456 4428 3474 4446
rect 3456 4446 3474 4464
rect 3456 4464 3474 4482
rect 3456 4482 3474 4500
rect 3456 4500 3474 4518
rect 3456 4518 3474 4536
rect 3456 4536 3474 4554
rect 3456 4554 3474 4572
rect 3456 4572 3474 4590
rect 3456 4590 3474 4608
rect 3456 4608 3474 4626
rect 3456 4626 3474 4644
rect 3456 4644 3474 4662
rect 3456 4662 3474 4680
rect 3456 4680 3474 4698
rect 3456 4698 3474 4716
rect 3456 4716 3474 4734
rect 3456 4734 3474 4752
rect 3456 4752 3474 4770
rect 3456 6642 3474 6660
rect 3456 6660 3474 6678
rect 3456 6678 3474 6696
rect 3456 6696 3474 6714
rect 3456 6714 3474 6732
rect 3456 6732 3474 6750
rect 3456 6750 3474 6768
rect 3456 6768 3474 6786
rect 3456 6786 3474 6804
rect 3456 6804 3474 6822
rect 3456 6822 3474 6840
rect 3456 6840 3474 6858
rect 3456 6858 3474 6876
rect 3456 6876 3474 6894
rect 3456 6894 3474 6912
rect 3456 6912 3474 6930
rect 3456 6930 3474 6948
rect 3456 6948 3474 6966
rect 3456 6966 3474 6984
rect 3456 6984 3474 7002
rect 3456 7002 3474 7020
rect 3456 7020 3474 7038
rect 3456 7038 3474 7056
rect 3456 7056 3474 7074
rect 3456 7074 3474 7092
rect 3456 7092 3474 7110
rect 3456 7110 3474 7128
rect 3456 7128 3474 7146
rect 3456 7146 3474 7164
rect 3456 7164 3474 7182
rect 3456 7182 3474 7200
rect 3456 7200 3474 7218
rect 3456 7218 3474 7236
rect 3456 7236 3474 7254
rect 3456 7254 3474 7272
rect 3474 18 3492 36
rect 3474 36 3492 54
rect 3474 54 3492 72
rect 3474 72 3492 90
rect 3474 90 3492 108
rect 3474 108 3492 126
rect 3474 126 3492 144
rect 3474 144 3492 162
rect 3474 162 3492 180
rect 3474 180 3492 198
rect 3474 198 3492 216
rect 3474 216 3492 234
rect 3474 234 3492 252
rect 3474 252 3492 270
rect 3474 270 3492 288
rect 3474 288 3492 306
rect 3474 306 3492 324
rect 3474 324 3492 342
rect 3474 342 3492 360
rect 3474 360 3492 378
rect 3474 378 3492 396
rect 3474 396 3492 414
rect 3474 414 3492 432
rect 3474 432 3492 450
rect 3474 450 3492 468
rect 3474 468 3492 486
rect 3474 486 3492 504
rect 3474 504 3492 522
rect 3474 522 3492 540
rect 3474 540 3492 558
rect 3474 558 3492 576
rect 3474 576 3492 594
rect 3474 594 3492 612
rect 3474 612 3492 630
rect 3474 810 3492 828
rect 3474 828 3492 846
rect 3474 846 3492 864
rect 3474 864 3492 882
rect 3474 882 3492 900
rect 3474 900 3492 918
rect 3474 918 3492 936
rect 3474 936 3492 954
rect 3474 954 3492 972
rect 3474 972 3492 990
rect 3474 990 3492 1008
rect 3474 1008 3492 1026
rect 3474 1026 3492 1044
rect 3474 1044 3492 1062
rect 3474 1062 3492 1080
rect 3474 1080 3492 1098
rect 3474 1098 3492 1116
rect 3474 1116 3492 1134
rect 3474 1134 3492 1152
rect 3474 1152 3492 1170
rect 3474 1170 3492 1188
rect 3474 1188 3492 1206
rect 3474 1404 3492 1422
rect 3474 1422 3492 1440
rect 3474 1440 3492 1458
rect 3474 1458 3492 1476
rect 3474 1476 3492 1494
rect 3474 1494 3492 1512
rect 3474 1512 3492 1530
rect 3474 1530 3492 1548
rect 3474 1548 3492 1566
rect 3474 1566 3492 1584
rect 3474 1584 3492 1602
rect 3474 1602 3492 1620
rect 3474 1620 3492 1638
rect 3474 1638 3492 1656
rect 3474 1656 3492 1674
rect 3474 1674 3492 1692
rect 3474 1692 3492 1710
rect 3474 1710 3492 1728
rect 3474 1728 3492 1746
rect 3474 1746 3492 1764
rect 3474 1764 3492 1782
rect 3474 1782 3492 1800
rect 3474 1800 3492 1818
rect 3474 1818 3492 1836
rect 3474 1836 3492 1854
rect 3474 1854 3492 1872
rect 3474 1872 3492 1890
rect 3474 1890 3492 1908
rect 3474 1908 3492 1926
rect 3474 1926 3492 1944
rect 3474 1944 3492 1962
rect 3474 1962 3492 1980
rect 3474 1980 3492 1998
rect 3474 1998 3492 2016
rect 3474 2016 3492 2034
rect 3474 2034 3492 2052
rect 3474 2052 3492 2070
rect 3474 2070 3492 2088
rect 3474 2088 3492 2106
rect 3474 2106 3492 2124
rect 3474 2124 3492 2142
rect 3474 2142 3492 2160
rect 3474 2160 3492 2178
rect 3474 2178 3492 2196
rect 3474 2196 3492 2214
rect 3474 2214 3492 2232
rect 3474 2232 3492 2250
rect 3474 2250 3492 2268
rect 3474 2268 3492 2286
rect 3474 2556 3492 2574
rect 3474 2574 3492 2592
rect 3474 2592 3492 2610
rect 3474 2610 3492 2628
rect 3474 2628 3492 2646
rect 3474 2646 3492 2664
rect 3474 2664 3492 2682
rect 3474 2682 3492 2700
rect 3474 2700 3492 2718
rect 3474 2718 3492 2736
rect 3474 2736 3492 2754
rect 3474 2754 3492 2772
rect 3474 2772 3492 2790
rect 3474 2790 3492 2808
rect 3474 2808 3492 2826
rect 3474 2826 3492 2844
rect 3474 2844 3492 2862
rect 3474 2862 3492 2880
rect 3474 2880 3492 2898
rect 3474 2898 3492 2916
rect 3474 2916 3492 2934
rect 3474 2934 3492 2952
rect 3474 2952 3492 2970
rect 3474 2970 3492 2988
rect 3474 2988 3492 3006
rect 3474 3006 3492 3024
rect 3474 3024 3492 3042
rect 3474 3042 3492 3060
rect 3474 3060 3492 3078
rect 3474 3078 3492 3096
rect 3474 3096 3492 3114
rect 3474 3114 3492 3132
rect 3474 3132 3492 3150
rect 3474 3150 3492 3168
rect 3474 3168 3492 3186
rect 3474 3186 3492 3204
rect 3474 3204 3492 3222
rect 3474 3222 3492 3240
rect 3474 3240 3492 3258
rect 3474 3258 3492 3276
rect 3474 3276 3492 3294
rect 3474 3294 3492 3312
rect 3474 3312 3492 3330
rect 3474 3330 3492 3348
rect 3474 3348 3492 3366
rect 3474 3366 3492 3384
rect 3474 3384 3492 3402
rect 3474 3402 3492 3420
rect 3474 3420 3492 3438
rect 3474 3438 3492 3456
rect 3474 3456 3492 3474
rect 3474 3474 3492 3492
rect 3474 3492 3492 3510
rect 3474 3510 3492 3528
rect 3474 3528 3492 3546
rect 3474 3546 3492 3564
rect 3474 3564 3492 3582
rect 3474 3582 3492 3600
rect 3474 3600 3492 3618
rect 3474 3618 3492 3636
rect 3474 3636 3492 3654
rect 3474 3654 3492 3672
rect 3474 3672 3492 3690
rect 3474 3690 3492 3708
rect 3474 3708 3492 3726
rect 3474 3726 3492 3744
rect 3474 3744 3492 3762
rect 3474 3762 3492 3780
rect 3474 3780 3492 3798
rect 3474 3798 3492 3816
rect 3474 3816 3492 3834
rect 3474 3834 3492 3852
rect 3474 3852 3492 3870
rect 3474 3870 3492 3888
rect 3474 3888 3492 3906
rect 3474 3906 3492 3924
rect 3474 3924 3492 3942
rect 3474 3942 3492 3960
rect 3474 3960 3492 3978
rect 3474 3978 3492 3996
rect 3474 3996 3492 4014
rect 3474 4014 3492 4032
rect 3474 4032 3492 4050
rect 3474 4050 3492 4068
rect 3474 4068 3492 4086
rect 3474 4086 3492 4104
rect 3474 4104 3492 4122
rect 3474 4122 3492 4140
rect 3474 4140 3492 4158
rect 3474 4158 3492 4176
rect 3474 4176 3492 4194
rect 3474 4194 3492 4212
rect 3474 4212 3492 4230
rect 3474 4230 3492 4248
rect 3474 4248 3492 4266
rect 3474 4266 3492 4284
rect 3474 4284 3492 4302
rect 3474 4302 3492 4320
rect 3474 4320 3492 4338
rect 3474 4338 3492 4356
rect 3474 4356 3492 4374
rect 3474 4374 3492 4392
rect 3474 4392 3492 4410
rect 3474 4410 3492 4428
rect 3474 4428 3492 4446
rect 3474 4446 3492 4464
rect 3474 4464 3492 4482
rect 3474 4482 3492 4500
rect 3474 4500 3492 4518
rect 3474 4518 3492 4536
rect 3474 4536 3492 4554
rect 3474 4554 3492 4572
rect 3474 4572 3492 4590
rect 3474 4590 3492 4608
rect 3474 4608 3492 4626
rect 3474 4626 3492 4644
rect 3474 4644 3492 4662
rect 3474 4662 3492 4680
rect 3474 4680 3492 4698
rect 3474 4698 3492 4716
rect 3474 4716 3492 4734
rect 3474 4734 3492 4752
rect 3474 4752 3492 4770
rect 3474 4770 3492 4788
rect 3474 4788 3492 4806
rect 3474 4806 3492 4824
rect 3474 6642 3492 6660
rect 3474 6660 3492 6678
rect 3474 6678 3492 6696
rect 3474 6696 3492 6714
rect 3474 6714 3492 6732
rect 3474 6732 3492 6750
rect 3474 6750 3492 6768
rect 3474 6768 3492 6786
rect 3474 6786 3492 6804
rect 3474 6804 3492 6822
rect 3474 6822 3492 6840
rect 3474 6840 3492 6858
rect 3474 6858 3492 6876
rect 3474 6876 3492 6894
rect 3474 6894 3492 6912
rect 3474 6912 3492 6930
rect 3474 6930 3492 6948
rect 3474 6948 3492 6966
rect 3474 6966 3492 6984
rect 3474 6984 3492 7002
rect 3474 7002 3492 7020
rect 3474 7020 3492 7038
rect 3474 7038 3492 7056
rect 3474 7056 3492 7074
rect 3474 7074 3492 7092
rect 3474 7092 3492 7110
rect 3474 7110 3492 7128
rect 3474 7128 3492 7146
rect 3474 7146 3492 7164
rect 3474 7164 3492 7182
rect 3474 7182 3492 7200
rect 3474 7200 3492 7218
rect 3474 7218 3492 7236
rect 3474 7236 3492 7254
rect 3474 7254 3492 7272
rect 3492 18 3510 36
rect 3492 36 3510 54
rect 3492 54 3510 72
rect 3492 72 3510 90
rect 3492 90 3510 108
rect 3492 108 3510 126
rect 3492 126 3510 144
rect 3492 144 3510 162
rect 3492 162 3510 180
rect 3492 180 3510 198
rect 3492 198 3510 216
rect 3492 216 3510 234
rect 3492 234 3510 252
rect 3492 252 3510 270
rect 3492 270 3510 288
rect 3492 288 3510 306
rect 3492 306 3510 324
rect 3492 324 3510 342
rect 3492 342 3510 360
rect 3492 360 3510 378
rect 3492 378 3510 396
rect 3492 396 3510 414
rect 3492 414 3510 432
rect 3492 432 3510 450
rect 3492 450 3510 468
rect 3492 468 3510 486
rect 3492 486 3510 504
rect 3492 504 3510 522
rect 3492 522 3510 540
rect 3492 540 3510 558
rect 3492 558 3510 576
rect 3492 576 3510 594
rect 3492 594 3510 612
rect 3492 612 3510 630
rect 3492 810 3510 828
rect 3492 828 3510 846
rect 3492 846 3510 864
rect 3492 864 3510 882
rect 3492 882 3510 900
rect 3492 900 3510 918
rect 3492 918 3510 936
rect 3492 936 3510 954
rect 3492 954 3510 972
rect 3492 972 3510 990
rect 3492 990 3510 1008
rect 3492 1008 3510 1026
rect 3492 1026 3510 1044
rect 3492 1044 3510 1062
rect 3492 1062 3510 1080
rect 3492 1080 3510 1098
rect 3492 1098 3510 1116
rect 3492 1116 3510 1134
rect 3492 1134 3510 1152
rect 3492 1152 3510 1170
rect 3492 1170 3510 1188
rect 3492 1188 3510 1206
rect 3492 1206 3510 1224
rect 3492 1422 3510 1440
rect 3492 1440 3510 1458
rect 3492 1458 3510 1476
rect 3492 1476 3510 1494
rect 3492 1494 3510 1512
rect 3492 1512 3510 1530
rect 3492 1530 3510 1548
rect 3492 1548 3510 1566
rect 3492 1566 3510 1584
rect 3492 1584 3510 1602
rect 3492 1602 3510 1620
rect 3492 1620 3510 1638
rect 3492 1638 3510 1656
rect 3492 1656 3510 1674
rect 3492 1674 3510 1692
rect 3492 1692 3510 1710
rect 3492 1710 3510 1728
rect 3492 1728 3510 1746
rect 3492 1746 3510 1764
rect 3492 1764 3510 1782
rect 3492 1782 3510 1800
rect 3492 1800 3510 1818
rect 3492 1818 3510 1836
rect 3492 1836 3510 1854
rect 3492 1854 3510 1872
rect 3492 1872 3510 1890
rect 3492 1890 3510 1908
rect 3492 1908 3510 1926
rect 3492 1926 3510 1944
rect 3492 1944 3510 1962
rect 3492 1962 3510 1980
rect 3492 1980 3510 1998
rect 3492 1998 3510 2016
rect 3492 2016 3510 2034
rect 3492 2034 3510 2052
rect 3492 2052 3510 2070
rect 3492 2070 3510 2088
rect 3492 2088 3510 2106
rect 3492 2106 3510 2124
rect 3492 2124 3510 2142
rect 3492 2142 3510 2160
rect 3492 2160 3510 2178
rect 3492 2178 3510 2196
rect 3492 2196 3510 2214
rect 3492 2214 3510 2232
rect 3492 2232 3510 2250
rect 3492 2250 3510 2268
rect 3492 2268 3510 2286
rect 3492 2286 3510 2304
rect 3492 2304 3510 2322
rect 3492 2592 3510 2610
rect 3492 2610 3510 2628
rect 3492 2628 3510 2646
rect 3492 2646 3510 2664
rect 3492 2664 3510 2682
rect 3492 2682 3510 2700
rect 3492 2700 3510 2718
rect 3492 2718 3510 2736
rect 3492 2736 3510 2754
rect 3492 2754 3510 2772
rect 3492 2772 3510 2790
rect 3492 2790 3510 2808
rect 3492 2808 3510 2826
rect 3492 2826 3510 2844
rect 3492 2844 3510 2862
rect 3492 2862 3510 2880
rect 3492 2880 3510 2898
rect 3492 2898 3510 2916
rect 3492 2916 3510 2934
rect 3492 2934 3510 2952
rect 3492 2952 3510 2970
rect 3492 2970 3510 2988
rect 3492 2988 3510 3006
rect 3492 3006 3510 3024
rect 3492 3024 3510 3042
rect 3492 3042 3510 3060
rect 3492 3060 3510 3078
rect 3492 3078 3510 3096
rect 3492 3096 3510 3114
rect 3492 3114 3510 3132
rect 3492 3132 3510 3150
rect 3492 3150 3510 3168
rect 3492 3168 3510 3186
rect 3492 3186 3510 3204
rect 3492 3204 3510 3222
rect 3492 3222 3510 3240
rect 3492 3240 3510 3258
rect 3492 3258 3510 3276
rect 3492 3276 3510 3294
rect 3492 3294 3510 3312
rect 3492 3312 3510 3330
rect 3492 3330 3510 3348
rect 3492 3348 3510 3366
rect 3492 3366 3510 3384
rect 3492 3384 3510 3402
rect 3492 3402 3510 3420
rect 3492 3420 3510 3438
rect 3492 3438 3510 3456
rect 3492 3456 3510 3474
rect 3492 3474 3510 3492
rect 3492 3492 3510 3510
rect 3492 3510 3510 3528
rect 3492 3528 3510 3546
rect 3492 3546 3510 3564
rect 3492 3564 3510 3582
rect 3492 3582 3510 3600
rect 3492 3600 3510 3618
rect 3492 3618 3510 3636
rect 3492 3636 3510 3654
rect 3492 3654 3510 3672
rect 3492 3672 3510 3690
rect 3492 3690 3510 3708
rect 3492 3708 3510 3726
rect 3492 3726 3510 3744
rect 3492 3744 3510 3762
rect 3492 3762 3510 3780
rect 3492 3780 3510 3798
rect 3492 3798 3510 3816
rect 3492 3816 3510 3834
rect 3492 3834 3510 3852
rect 3492 3852 3510 3870
rect 3492 3870 3510 3888
rect 3492 3888 3510 3906
rect 3492 3906 3510 3924
rect 3492 3924 3510 3942
rect 3492 3942 3510 3960
rect 3492 3960 3510 3978
rect 3492 3978 3510 3996
rect 3492 3996 3510 4014
rect 3492 4014 3510 4032
rect 3492 4032 3510 4050
rect 3492 4050 3510 4068
rect 3492 4068 3510 4086
rect 3492 4086 3510 4104
rect 3492 4104 3510 4122
rect 3492 4122 3510 4140
rect 3492 4140 3510 4158
rect 3492 4158 3510 4176
rect 3492 4176 3510 4194
rect 3492 4194 3510 4212
rect 3492 4212 3510 4230
rect 3492 4230 3510 4248
rect 3492 4248 3510 4266
rect 3492 4266 3510 4284
rect 3492 4284 3510 4302
rect 3492 4302 3510 4320
rect 3492 4320 3510 4338
rect 3492 4338 3510 4356
rect 3492 4356 3510 4374
rect 3492 4374 3510 4392
rect 3492 4392 3510 4410
rect 3492 4410 3510 4428
rect 3492 4428 3510 4446
rect 3492 4446 3510 4464
rect 3492 4464 3510 4482
rect 3492 4482 3510 4500
rect 3492 4500 3510 4518
rect 3492 4518 3510 4536
rect 3492 4536 3510 4554
rect 3492 4554 3510 4572
rect 3492 4572 3510 4590
rect 3492 4590 3510 4608
rect 3492 4608 3510 4626
rect 3492 4626 3510 4644
rect 3492 4644 3510 4662
rect 3492 4662 3510 4680
rect 3492 4680 3510 4698
rect 3492 4698 3510 4716
rect 3492 4716 3510 4734
rect 3492 4734 3510 4752
rect 3492 4752 3510 4770
rect 3492 4770 3510 4788
rect 3492 4788 3510 4806
rect 3492 4806 3510 4824
rect 3492 4824 3510 4842
rect 3492 4842 3510 4860
rect 3492 6642 3510 6660
rect 3492 6660 3510 6678
rect 3492 6678 3510 6696
rect 3492 6696 3510 6714
rect 3492 6714 3510 6732
rect 3492 6732 3510 6750
rect 3492 6750 3510 6768
rect 3492 6768 3510 6786
rect 3492 6786 3510 6804
rect 3492 6804 3510 6822
rect 3492 6822 3510 6840
rect 3492 6840 3510 6858
rect 3492 6858 3510 6876
rect 3492 6876 3510 6894
rect 3492 6894 3510 6912
rect 3492 6912 3510 6930
rect 3492 6930 3510 6948
rect 3492 6948 3510 6966
rect 3492 6966 3510 6984
rect 3492 6984 3510 7002
rect 3492 7002 3510 7020
rect 3492 7020 3510 7038
rect 3492 7038 3510 7056
rect 3492 7056 3510 7074
rect 3492 7074 3510 7092
rect 3492 7092 3510 7110
rect 3492 7110 3510 7128
rect 3492 7128 3510 7146
rect 3492 7146 3510 7164
rect 3492 7164 3510 7182
rect 3492 7182 3510 7200
rect 3492 7200 3510 7218
rect 3492 7218 3510 7236
rect 3492 7236 3510 7254
rect 3492 7254 3510 7272
rect 3510 18 3528 36
rect 3510 36 3528 54
rect 3510 54 3528 72
rect 3510 72 3528 90
rect 3510 90 3528 108
rect 3510 108 3528 126
rect 3510 126 3528 144
rect 3510 144 3528 162
rect 3510 162 3528 180
rect 3510 180 3528 198
rect 3510 198 3528 216
rect 3510 216 3528 234
rect 3510 234 3528 252
rect 3510 252 3528 270
rect 3510 270 3528 288
rect 3510 288 3528 306
rect 3510 306 3528 324
rect 3510 324 3528 342
rect 3510 342 3528 360
rect 3510 360 3528 378
rect 3510 378 3528 396
rect 3510 396 3528 414
rect 3510 414 3528 432
rect 3510 432 3528 450
rect 3510 450 3528 468
rect 3510 468 3528 486
rect 3510 486 3528 504
rect 3510 504 3528 522
rect 3510 522 3528 540
rect 3510 540 3528 558
rect 3510 558 3528 576
rect 3510 576 3528 594
rect 3510 594 3528 612
rect 3510 810 3528 828
rect 3510 828 3528 846
rect 3510 846 3528 864
rect 3510 864 3528 882
rect 3510 882 3528 900
rect 3510 900 3528 918
rect 3510 918 3528 936
rect 3510 936 3528 954
rect 3510 954 3528 972
rect 3510 972 3528 990
rect 3510 990 3528 1008
rect 3510 1008 3528 1026
rect 3510 1026 3528 1044
rect 3510 1044 3528 1062
rect 3510 1062 3528 1080
rect 3510 1080 3528 1098
rect 3510 1098 3528 1116
rect 3510 1116 3528 1134
rect 3510 1134 3528 1152
rect 3510 1152 3528 1170
rect 3510 1170 3528 1188
rect 3510 1188 3528 1206
rect 3510 1206 3528 1224
rect 3510 1440 3528 1458
rect 3510 1458 3528 1476
rect 3510 1476 3528 1494
rect 3510 1494 3528 1512
rect 3510 1512 3528 1530
rect 3510 1530 3528 1548
rect 3510 1548 3528 1566
rect 3510 1566 3528 1584
rect 3510 1584 3528 1602
rect 3510 1602 3528 1620
rect 3510 1620 3528 1638
rect 3510 1638 3528 1656
rect 3510 1656 3528 1674
rect 3510 1674 3528 1692
rect 3510 1692 3528 1710
rect 3510 1710 3528 1728
rect 3510 1728 3528 1746
rect 3510 1746 3528 1764
rect 3510 1764 3528 1782
rect 3510 1782 3528 1800
rect 3510 1800 3528 1818
rect 3510 1818 3528 1836
rect 3510 1836 3528 1854
rect 3510 1854 3528 1872
rect 3510 1872 3528 1890
rect 3510 1890 3528 1908
rect 3510 1908 3528 1926
rect 3510 1926 3528 1944
rect 3510 1944 3528 1962
rect 3510 1962 3528 1980
rect 3510 1980 3528 1998
rect 3510 1998 3528 2016
rect 3510 2016 3528 2034
rect 3510 2034 3528 2052
rect 3510 2052 3528 2070
rect 3510 2070 3528 2088
rect 3510 2088 3528 2106
rect 3510 2106 3528 2124
rect 3510 2124 3528 2142
rect 3510 2142 3528 2160
rect 3510 2160 3528 2178
rect 3510 2178 3528 2196
rect 3510 2196 3528 2214
rect 3510 2214 3528 2232
rect 3510 2232 3528 2250
rect 3510 2250 3528 2268
rect 3510 2268 3528 2286
rect 3510 2286 3528 2304
rect 3510 2304 3528 2322
rect 3510 2322 3528 2340
rect 3510 2610 3528 2628
rect 3510 2628 3528 2646
rect 3510 2646 3528 2664
rect 3510 2664 3528 2682
rect 3510 2682 3528 2700
rect 3510 2700 3528 2718
rect 3510 2718 3528 2736
rect 3510 2736 3528 2754
rect 3510 2754 3528 2772
rect 3510 2772 3528 2790
rect 3510 2790 3528 2808
rect 3510 2808 3528 2826
rect 3510 2826 3528 2844
rect 3510 2844 3528 2862
rect 3510 2862 3528 2880
rect 3510 2880 3528 2898
rect 3510 2898 3528 2916
rect 3510 2916 3528 2934
rect 3510 2934 3528 2952
rect 3510 2952 3528 2970
rect 3510 2970 3528 2988
rect 3510 2988 3528 3006
rect 3510 3006 3528 3024
rect 3510 3024 3528 3042
rect 3510 3042 3528 3060
rect 3510 3060 3528 3078
rect 3510 3078 3528 3096
rect 3510 3096 3528 3114
rect 3510 3114 3528 3132
rect 3510 3132 3528 3150
rect 3510 3150 3528 3168
rect 3510 3168 3528 3186
rect 3510 3186 3528 3204
rect 3510 3204 3528 3222
rect 3510 3222 3528 3240
rect 3510 3240 3528 3258
rect 3510 3258 3528 3276
rect 3510 3276 3528 3294
rect 3510 3294 3528 3312
rect 3510 3312 3528 3330
rect 3510 3330 3528 3348
rect 3510 3348 3528 3366
rect 3510 3366 3528 3384
rect 3510 3384 3528 3402
rect 3510 3402 3528 3420
rect 3510 3420 3528 3438
rect 3510 3438 3528 3456
rect 3510 3456 3528 3474
rect 3510 3474 3528 3492
rect 3510 3492 3528 3510
rect 3510 3510 3528 3528
rect 3510 3528 3528 3546
rect 3510 3546 3528 3564
rect 3510 3564 3528 3582
rect 3510 3582 3528 3600
rect 3510 3600 3528 3618
rect 3510 3618 3528 3636
rect 3510 3636 3528 3654
rect 3510 3654 3528 3672
rect 3510 3672 3528 3690
rect 3510 3690 3528 3708
rect 3510 3708 3528 3726
rect 3510 3726 3528 3744
rect 3510 3744 3528 3762
rect 3510 3762 3528 3780
rect 3510 3780 3528 3798
rect 3510 3798 3528 3816
rect 3510 3816 3528 3834
rect 3510 3834 3528 3852
rect 3510 3852 3528 3870
rect 3510 3870 3528 3888
rect 3510 3888 3528 3906
rect 3510 3906 3528 3924
rect 3510 3924 3528 3942
rect 3510 3942 3528 3960
rect 3510 3960 3528 3978
rect 3510 3978 3528 3996
rect 3510 3996 3528 4014
rect 3510 4014 3528 4032
rect 3510 4032 3528 4050
rect 3510 4050 3528 4068
rect 3510 4068 3528 4086
rect 3510 4086 3528 4104
rect 3510 4104 3528 4122
rect 3510 4122 3528 4140
rect 3510 4140 3528 4158
rect 3510 4158 3528 4176
rect 3510 4176 3528 4194
rect 3510 4194 3528 4212
rect 3510 4212 3528 4230
rect 3510 4230 3528 4248
rect 3510 4248 3528 4266
rect 3510 4266 3528 4284
rect 3510 4284 3528 4302
rect 3510 4302 3528 4320
rect 3510 4320 3528 4338
rect 3510 4338 3528 4356
rect 3510 4356 3528 4374
rect 3510 4374 3528 4392
rect 3510 4392 3528 4410
rect 3510 4410 3528 4428
rect 3510 4428 3528 4446
rect 3510 4446 3528 4464
rect 3510 4464 3528 4482
rect 3510 4482 3528 4500
rect 3510 4500 3528 4518
rect 3510 4518 3528 4536
rect 3510 4536 3528 4554
rect 3510 4554 3528 4572
rect 3510 4572 3528 4590
rect 3510 4590 3528 4608
rect 3510 4608 3528 4626
rect 3510 4626 3528 4644
rect 3510 4644 3528 4662
rect 3510 4662 3528 4680
rect 3510 4680 3528 4698
rect 3510 4698 3528 4716
rect 3510 4716 3528 4734
rect 3510 4734 3528 4752
rect 3510 4752 3528 4770
rect 3510 4770 3528 4788
rect 3510 4788 3528 4806
rect 3510 4806 3528 4824
rect 3510 4824 3528 4842
rect 3510 4842 3528 4860
rect 3510 4860 3528 4878
rect 3510 4878 3528 4896
rect 3510 4896 3528 4914
rect 3510 6642 3528 6660
rect 3510 6660 3528 6678
rect 3510 6678 3528 6696
rect 3510 6696 3528 6714
rect 3510 6714 3528 6732
rect 3510 6732 3528 6750
rect 3510 6750 3528 6768
rect 3510 6768 3528 6786
rect 3510 6786 3528 6804
rect 3510 6804 3528 6822
rect 3510 6822 3528 6840
rect 3510 6840 3528 6858
rect 3510 6858 3528 6876
rect 3510 6876 3528 6894
rect 3510 6894 3528 6912
rect 3510 6912 3528 6930
rect 3510 6930 3528 6948
rect 3510 6948 3528 6966
rect 3510 6966 3528 6984
rect 3510 6984 3528 7002
rect 3510 7002 3528 7020
rect 3510 7020 3528 7038
rect 3510 7038 3528 7056
rect 3510 7056 3528 7074
rect 3510 7074 3528 7092
rect 3510 7092 3528 7110
rect 3510 7110 3528 7128
rect 3510 7128 3528 7146
rect 3510 7146 3528 7164
rect 3510 7164 3528 7182
rect 3510 7182 3528 7200
rect 3510 7200 3528 7218
rect 3510 7218 3528 7236
rect 3510 7236 3528 7254
rect 3510 7254 3528 7272
rect 3528 18 3546 36
rect 3528 36 3546 54
rect 3528 54 3546 72
rect 3528 72 3546 90
rect 3528 90 3546 108
rect 3528 108 3546 126
rect 3528 126 3546 144
rect 3528 144 3546 162
rect 3528 162 3546 180
rect 3528 180 3546 198
rect 3528 198 3546 216
rect 3528 216 3546 234
rect 3528 234 3546 252
rect 3528 252 3546 270
rect 3528 270 3546 288
rect 3528 288 3546 306
rect 3528 306 3546 324
rect 3528 324 3546 342
rect 3528 342 3546 360
rect 3528 360 3546 378
rect 3528 378 3546 396
rect 3528 396 3546 414
rect 3528 414 3546 432
rect 3528 432 3546 450
rect 3528 450 3546 468
rect 3528 468 3546 486
rect 3528 486 3546 504
rect 3528 504 3546 522
rect 3528 522 3546 540
rect 3528 540 3546 558
rect 3528 558 3546 576
rect 3528 576 3546 594
rect 3528 594 3546 612
rect 3528 828 3546 846
rect 3528 846 3546 864
rect 3528 864 3546 882
rect 3528 882 3546 900
rect 3528 900 3546 918
rect 3528 918 3546 936
rect 3528 936 3546 954
rect 3528 954 3546 972
rect 3528 972 3546 990
rect 3528 990 3546 1008
rect 3528 1008 3546 1026
rect 3528 1026 3546 1044
rect 3528 1044 3546 1062
rect 3528 1062 3546 1080
rect 3528 1080 3546 1098
rect 3528 1098 3546 1116
rect 3528 1116 3546 1134
rect 3528 1134 3546 1152
rect 3528 1152 3546 1170
rect 3528 1170 3546 1188
rect 3528 1188 3546 1206
rect 3528 1206 3546 1224
rect 3528 1224 3546 1242
rect 3528 1458 3546 1476
rect 3528 1476 3546 1494
rect 3528 1494 3546 1512
rect 3528 1512 3546 1530
rect 3528 1530 3546 1548
rect 3528 1548 3546 1566
rect 3528 1566 3546 1584
rect 3528 1584 3546 1602
rect 3528 1602 3546 1620
rect 3528 1620 3546 1638
rect 3528 1638 3546 1656
rect 3528 1656 3546 1674
rect 3528 1674 3546 1692
rect 3528 1692 3546 1710
rect 3528 1710 3546 1728
rect 3528 1728 3546 1746
rect 3528 1746 3546 1764
rect 3528 1764 3546 1782
rect 3528 1782 3546 1800
rect 3528 1800 3546 1818
rect 3528 1818 3546 1836
rect 3528 1836 3546 1854
rect 3528 1854 3546 1872
rect 3528 1872 3546 1890
rect 3528 1890 3546 1908
rect 3528 1908 3546 1926
rect 3528 1926 3546 1944
rect 3528 1944 3546 1962
rect 3528 1962 3546 1980
rect 3528 1980 3546 1998
rect 3528 1998 3546 2016
rect 3528 2016 3546 2034
rect 3528 2034 3546 2052
rect 3528 2052 3546 2070
rect 3528 2070 3546 2088
rect 3528 2088 3546 2106
rect 3528 2106 3546 2124
rect 3528 2124 3546 2142
rect 3528 2142 3546 2160
rect 3528 2160 3546 2178
rect 3528 2178 3546 2196
rect 3528 2196 3546 2214
rect 3528 2214 3546 2232
rect 3528 2232 3546 2250
rect 3528 2250 3546 2268
rect 3528 2268 3546 2286
rect 3528 2286 3546 2304
rect 3528 2304 3546 2322
rect 3528 2322 3546 2340
rect 3528 2340 3546 2358
rect 3528 2358 3546 2376
rect 3528 2646 3546 2664
rect 3528 2664 3546 2682
rect 3528 2682 3546 2700
rect 3528 2700 3546 2718
rect 3528 2718 3546 2736
rect 3528 2736 3546 2754
rect 3528 2754 3546 2772
rect 3528 2772 3546 2790
rect 3528 2790 3546 2808
rect 3528 2808 3546 2826
rect 3528 2826 3546 2844
rect 3528 2844 3546 2862
rect 3528 2862 3546 2880
rect 3528 2880 3546 2898
rect 3528 2898 3546 2916
rect 3528 2916 3546 2934
rect 3528 2934 3546 2952
rect 3528 2952 3546 2970
rect 3528 2970 3546 2988
rect 3528 2988 3546 3006
rect 3528 3006 3546 3024
rect 3528 3024 3546 3042
rect 3528 3042 3546 3060
rect 3528 3060 3546 3078
rect 3528 3078 3546 3096
rect 3528 3096 3546 3114
rect 3528 3114 3546 3132
rect 3528 3132 3546 3150
rect 3528 3150 3546 3168
rect 3528 3168 3546 3186
rect 3528 3186 3546 3204
rect 3528 3204 3546 3222
rect 3528 3222 3546 3240
rect 3528 3240 3546 3258
rect 3528 3258 3546 3276
rect 3528 3276 3546 3294
rect 3528 3294 3546 3312
rect 3528 3312 3546 3330
rect 3528 3330 3546 3348
rect 3528 3348 3546 3366
rect 3528 3366 3546 3384
rect 3528 3384 3546 3402
rect 3528 3402 3546 3420
rect 3528 3420 3546 3438
rect 3528 3438 3546 3456
rect 3528 3456 3546 3474
rect 3528 3474 3546 3492
rect 3528 3492 3546 3510
rect 3528 3510 3546 3528
rect 3528 3528 3546 3546
rect 3528 3546 3546 3564
rect 3528 3564 3546 3582
rect 3528 3582 3546 3600
rect 3528 3600 3546 3618
rect 3528 3618 3546 3636
rect 3528 3636 3546 3654
rect 3528 3654 3546 3672
rect 3528 3672 3546 3690
rect 3528 3690 3546 3708
rect 3528 3708 3546 3726
rect 3528 3726 3546 3744
rect 3528 3744 3546 3762
rect 3528 3762 3546 3780
rect 3528 3780 3546 3798
rect 3528 3798 3546 3816
rect 3528 3816 3546 3834
rect 3528 3834 3546 3852
rect 3528 3852 3546 3870
rect 3528 3870 3546 3888
rect 3528 3888 3546 3906
rect 3528 3906 3546 3924
rect 3528 3924 3546 3942
rect 3528 3942 3546 3960
rect 3528 3960 3546 3978
rect 3528 3978 3546 3996
rect 3528 3996 3546 4014
rect 3528 4014 3546 4032
rect 3528 4032 3546 4050
rect 3528 4050 3546 4068
rect 3528 4068 3546 4086
rect 3528 4086 3546 4104
rect 3528 4104 3546 4122
rect 3528 4122 3546 4140
rect 3528 4140 3546 4158
rect 3528 4158 3546 4176
rect 3528 4176 3546 4194
rect 3528 4194 3546 4212
rect 3528 4212 3546 4230
rect 3528 4230 3546 4248
rect 3528 4248 3546 4266
rect 3528 4266 3546 4284
rect 3528 4284 3546 4302
rect 3528 4302 3546 4320
rect 3528 4320 3546 4338
rect 3528 4338 3546 4356
rect 3528 4356 3546 4374
rect 3528 4374 3546 4392
rect 3528 4392 3546 4410
rect 3528 4410 3546 4428
rect 3528 4428 3546 4446
rect 3528 4446 3546 4464
rect 3528 4464 3546 4482
rect 3528 4482 3546 4500
rect 3528 4500 3546 4518
rect 3528 4518 3546 4536
rect 3528 4536 3546 4554
rect 3528 4554 3546 4572
rect 3528 4572 3546 4590
rect 3528 4590 3546 4608
rect 3528 4608 3546 4626
rect 3528 4626 3546 4644
rect 3528 4644 3546 4662
rect 3528 4662 3546 4680
rect 3528 4680 3546 4698
rect 3528 4698 3546 4716
rect 3528 4716 3546 4734
rect 3528 4734 3546 4752
rect 3528 4752 3546 4770
rect 3528 4770 3546 4788
rect 3528 4788 3546 4806
rect 3528 4806 3546 4824
rect 3528 4824 3546 4842
rect 3528 4842 3546 4860
rect 3528 4860 3546 4878
rect 3528 4878 3546 4896
rect 3528 4896 3546 4914
rect 3528 4914 3546 4932
rect 3528 4932 3546 4950
rect 3528 4950 3546 4968
rect 3528 6642 3546 6660
rect 3528 6660 3546 6678
rect 3528 6678 3546 6696
rect 3528 6696 3546 6714
rect 3528 6714 3546 6732
rect 3528 6732 3546 6750
rect 3528 6750 3546 6768
rect 3528 6768 3546 6786
rect 3528 6786 3546 6804
rect 3528 6804 3546 6822
rect 3528 6822 3546 6840
rect 3528 6840 3546 6858
rect 3528 6858 3546 6876
rect 3528 6876 3546 6894
rect 3528 6894 3546 6912
rect 3528 6912 3546 6930
rect 3528 6930 3546 6948
rect 3528 6948 3546 6966
rect 3528 6966 3546 6984
rect 3528 6984 3546 7002
rect 3528 7002 3546 7020
rect 3528 7020 3546 7038
rect 3528 7038 3546 7056
rect 3528 7056 3546 7074
rect 3528 7074 3546 7092
rect 3528 7092 3546 7110
rect 3528 7110 3546 7128
rect 3528 7128 3546 7146
rect 3528 7146 3546 7164
rect 3528 7164 3546 7182
rect 3528 7182 3546 7200
rect 3528 7200 3546 7218
rect 3528 7218 3546 7236
rect 3528 7236 3546 7254
rect 3528 7254 3546 7272
rect 3546 18 3564 36
rect 3546 36 3564 54
rect 3546 54 3564 72
rect 3546 72 3564 90
rect 3546 90 3564 108
rect 3546 108 3564 126
rect 3546 126 3564 144
rect 3546 144 3564 162
rect 3546 162 3564 180
rect 3546 180 3564 198
rect 3546 198 3564 216
rect 3546 216 3564 234
rect 3546 234 3564 252
rect 3546 252 3564 270
rect 3546 270 3564 288
rect 3546 288 3564 306
rect 3546 306 3564 324
rect 3546 324 3564 342
rect 3546 342 3564 360
rect 3546 360 3564 378
rect 3546 378 3564 396
rect 3546 396 3564 414
rect 3546 414 3564 432
rect 3546 432 3564 450
rect 3546 450 3564 468
rect 3546 468 3564 486
rect 3546 486 3564 504
rect 3546 504 3564 522
rect 3546 522 3564 540
rect 3546 540 3564 558
rect 3546 558 3564 576
rect 3546 576 3564 594
rect 3546 594 3564 612
rect 3546 828 3564 846
rect 3546 846 3564 864
rect 3546 864 3564 882
rect 3546 882 3564 900
rect 3546 900 3564 918
rect 3546 918 3564 936
rect 3546 936 3564 954
rect 3546 954 3564 972
rect 3546 972 3564 990
rect 3546 990 3564 1008
rect 3546 1008 3564 1026
rect 3546 1026 3564 1044
rect 3546 1044 3564 1062
rect 3546 1062 3564 1080
rect 3546 1080 3564 1098
rect 3546 1098 3564 1116
rect 3546 1116 3564 1134
rect 3546 1134 3564 1152
rect 3546 1152 3564 1170
rect 3546 1170 3564 1188
rect 3546 1188 3564 1206
rect 3546 1206 3564 1224
rect 3546 1224 3564 1242
rect 3546 1242 3564 1260
rect 3546 1458 3564 1476
rect 3546 1476 3564 1494
rect 3546 1494 3564 1512
rect 3546 1512 3564 1530
rect 3546 1530 3564 1548
rect 3546 1548 3564 1566
rect 3546 1566 3564 1584
rect 3546 1584 3564 1602
rect 3546 1602 3564 1620
rect 3546 1620 3564 1638
rect 3546 1638 3564 1656
rect 3546 1656 3564 1674
rect 3546 1674 3564 1692
rect 3546 1692 3564 1710
rect 3546 1710 3564 1728
rect 3546 1728 3564 1746
rect 3546 1746 3564 1764
rect 3546 1764 3564 1782
rect 3546 1782 3564 1800
rect 3546 1800 3564 1818
rect 3546 1818 3564 1836
rect 3546 1836 3564 1854
rect 3546 1854 3564 1872
rect 3546 1872 3564 1890
rect 3546 1890 3564 1908
rect 3546 1908 3564 1926
rect 3546 1926 3564 1944
rect 3546 1944 3564 1962
rect 3546 1962 3564 1980
rect 3546 1980 3564 1998
rect 3546 1998 3564 2016
rect 3546 2016 3564 2034
rect 3546 2034 3564 2052
rect 3546 2052 3564 2070
rect 3546 2070 3564 2088
rect 3546 2088 3564 2106
rect 3546 2106 3564 2124
rect 3546 2124 3564 2142
rect 3546 2142 3564 2160
rect 3546 2160 3564 2178
rect 3546 2178 3564 2196
rect 3546 2196 3564 2214
rect 3546 2214 3564 2232
rect 3546 2232 3564 2250
rect 3546 2250 3564 2268
rect 3546 2268 3564 2286
rect 3546 2286 3564 2304
rect 3546 2304 3564 2322
rect 3546 2322 3564 2340
rect 3546 2340 3564 2358
rect 3546 2358 3564 2376
rect 3546 2376 3564 2394
rect 3546 2394 3564 2412
rect 3546 2664 3564 2682
rect 3546 2682 3564 2700
rect 3546 2700 3564 2718
rect 3546 2718 3564 2736
rect 3546 2736 3564 2754
rect 3546 2754 3564 2772
rect 3546 2772 3564 2790
rect 3546 2790 3564 2808
rect 3546 2808 3564 2826
rect 3546 2826 3564 2844
rect 3546 2844 3564 2862
rect 3546 2862 3564 2880
rect 3546 2880 3564 2898
rect 3546 2898 3564 2916
rect 3546 2916 3564 2934
rect 3546 2934 3564 2952
rect 3546 2952 3564 2970
rect 3546 2970 3564 2988
rect 3546 2988 3564 3006
rect 3546 3006 3564 3024
rect 3546 3024 3564 3042
rect 3546 3042 3564 3060
rect 3546 3060 3564 3078
rect 3546 3078 3564 3096
rect 3546 3096 3564 3114
rect 3546 3114 3564 3132
rect 3546 3132 3564 3150
rect 3546 3150 3564 3168
rect 3546 3168 3564 3186
rect 3546 3186 3564 3204
rect 3546 3204 3564 3222
rect 3546 3222 3564 3240
rect 3546 3240 3564 3258
rect 3546 3258 3564 3276
rect 3546 3276 3564 3294
rect 3546 3294 3564 3312
rect 3546 3312 3564 3330
rect 3546 3330 3564 3348
rect 3546 3348 3564 3366
rect 3546 3366 3564 3384
rect 3546 3384 3564 3402
rect 3546 3402 3564 3420
rect 3546 3420 3564 3438
rect 3546 3438 3564 3456
rect 3546 3456 3564 3474
rect 3546 3474 3564 3492
rect 3546 3492 3564 3510
rect 3546 3510 3564 3528
rect 3546 3528 3564 3546
rect 3546 3546 3564 3564
rect 3546 3564 3564 3582
rect 3546 3582 3564 3600
rect 3546 3600 3564 3618
rect 3546 3618 3564 3636
rect 3546 3636 3564 3654
rect 3546 3654 3564 3672
rect 3546 3672 3564 3690
rect 3546 3690 3564 3708
rect 3546 3708 3564 3726
rect 3546 3726 3564 3744
rect 3546 3744 3564 3762
rect 3546 3762 3564 3780
rect 3546 3780 3564 3798
rect 3546 3798 3564 3816
rect 3546 3816 3564 3834
rect 3546 3834 3564 3852
rect 3546 3852 3564 3870
rect 3546 3870 3564 3888
rect 3546 3888 3564 3906
rect 3546 3906 3564 3924
rect 3546 3924 3564 3942
rect 3546 3942 3564 3960
rect 3546 3960 3564 3978
rect 3546 3978 3564 3996
rect 3546 3996 3564 4014
rect 3546 4014 3564 4032
rect 3546 4032 3564 4050
rect 3546 4050 3564 4068
rect 3546 4068 3564 4086
rect 3546 4086 3564 4104
rect 3546 4104 3564 4122
rect 3546 4122 3564 4140
rect 3546 4140 3564 4158
rect 3546 4158 3564 4176
rect 3546 4176 3564 4194
rect 3546 4194 3564 4212
rect 3546 4212 3564 4230
rect 3546 4230 3564 4248
rect 3546 4248 3564 4266
rect 3546 4266 3564 4284
rect 3546 4284 3564 4302
rect 3546 4302 3564 4320
rect 3546 4320 3564 4338
rect 3546 4338 3564 4356
rect 3546 4356 3564 4374
rect 3546 4374 3564 4392
rect 3546 4392 3564 4410
rect 3546 4410 3564 4428
rect 3546 4428 3564 4446
rect 3546 4446 3564 4464
rect 3546 4464 3564 4482
rect 3546 4482 3564 4500
rect 3546 4500 3564 4518
rect 3546 4518 3564 4536
rect 3546 4536 3564 4554
rect 3546 4554 3564 4572
rect 3546 4572 3564 4590
rect 3546 4590 3564 4608
rect 3546 4608 3564 4626
rect 3546 4626 3564 4644
rect 3546 4644 3564 4662
rect 3546 4662 3564 4680
rect 3546 4680 3564 4698
rect 3546 4698 3564 4716
rect 3546 4716 3564 4734
rect 3546 4734 3564 4752
rect 3546 4752 3564 4770
rect 3546 4770 3564 4788
rect 3546 4788 3564 4806
rect 3546 4806 3564 4824
rect 3546 4824 3564 4842
rect 3546 4842 3564 4860
rect 3546 4860 3564 4878
rect 3546 4878 3564 4896
rect 3546 4896 3564 4914
rect 3546 4914 3564 4932
rect 3546 4932 3564 4950
rect 3546 4950 3564 4968
rect 3546 4968 3564 4986
rect 3546 4986 3564 5004
rect 3546 6642 3564 6660
rect 3546 6660 3564 6678
rect 3546 6678 3564 6696
rect 3546 6696 3564 6714
rect 3546 6714 3564 6732
rect 3546 6732 3564 6750
rect 3546 6750 3564 6768
rect 3546 6768 3564 6786
rect 3546 6786 3564 6804
rect 3546 6804 3564 6822
rect 3546 6822 3564 6840
rect 3546 6840 3564 6858
rect 3546 6858 3564 6876
rect 3546 6876 3564 6894
rect 3546 6894 3564 6912
rect 3546 6912 3564 6930
rect 3546 6930 3564 6948
rect 3546 6948 3564 6966
rect 3546 6966 3564 6984
rect 3546 6984 3564 7002
rect 3546 7002 3564 7020
rect 3546 7020 3564 7038
rect 3546 7038 3564 7056
rect 3546 7056 3564 7074
rect 3546 7074 3564 7092
rect 3546 7092 3564 7110
rect 3546 7110 3564 7128
rect 3546 7128 3564 7146
rect 3546 7146 3564 7164
rect 3546 7164 3564 7182
rect 3546 7182 3564 7200
rect 3546 7200 3564 7218
rect 3546 7218 3564 7236
rect 3546 7236 3564 7254
rect 3546 7254 3564 7272
rect 3564 18 3582 36
rect 3564 36 3582 54
rect 3564 54 3582 72
rect 3564 72 3582 90
rect 3564 90 3582 108
rect 3564 108 3582 126
rect 3564 126 3582 144
rect 3564 144 3582 162
rect 3564 162 3582 180
rect 3564 180 3582 198
rect 3564 198 3582 216
rect 3564 216 3582 234
rect 3564 234 3582 252
rect 3564 252 3582 270
rect 3564 270 3582 288
rect 3564 288 3582 306
rect 3564 306 3582 324
rect 3564 324 3582 342
rect 3564 342 3582 360
rect 3564 360 3582 378
rect 3564 378 3582 396
rect 3564 396 3582 414
rect 3564 414 3582 432
rect 3564 432 3582 450
rect 3564 450 3582 468
rect 3564 468 3582 486
rect 3564 486 3582 504
rect 3564 504 3582 522
rect 3564 522 3582 540
rect 3564 540 3582 558
rect 3564 558 3582 576
rect 3564 576 3582 594
rect 3564 594 3582 612
rect 3564 828 3582 846
rect 3564 846 3582 864
rect 3564 864 3582 882
rect 3564 882 3582 900
rect 3564 900 3582 918
rect 3564 918 3582 936
rect 3564 936 3582 954
rect 3564 954 3582 972
rect 3564 972 3582 990
rect 3564 990 3582 1008
rect 3564 1008 3582 1026
rect 3564 1026 3582 1044
rect 3564 1044 3582 1062
rect 3564 1062 3582 1080
rect 3564 1080 3582 1098
rect 3564 1098 3582 1116
rect 3564 1116 3582 1134
rect 3564 1134 3582 1152
rect 3564 1152 3582 1170
rect 3564 1170 3582 1188
rect 3564 1188 3582 1206
rect 3564 1206 3582 1224
rect 3564 1224 3582 1242
rect 3564 1242 3582 1260
rect 3564 1476 3582 1494
rect 3564 1494 3582 1512
rect 3564 1512 3582 1530
rect 3564 1530 3582 1548
rect 3564 1548 3582 1566
rect 3564 1566 3582 1584
rect 3564 1584 3582 1602
rect 3564 1602 3582 1620
rect 3564 1620 3582 1638
rect 3564 1638 3582 1656
rect 3564 1656 3582 1674
rect 3564 1674 3582 1692
rect 3564 1692 3582 1710
rect 3564 1710 3582 1728
rect 3564 1728 3582 1746
rect 3564 1746 3582 1764
rect 3564 1764 3582 1782
rect 3564 1782 3582 1800
rect 3564 1800 3582 1818
rect 3564 1818 3582 1836
rect 3564 1836 3582 1854
rect 3564 1854 3582 1872
rect 3564 1872 3582 1890
rect 3564 1890 3582 1908
rect 3564 1908 3582 1926
rect 3564 1926 3582 1944
rect 3564 1944 3582 1962
rect 3564 1962 3582 1980
rect 3564 1980 3582 1998
rect 3564 1998 3582 2016
rect 3564 2016 3582 2034
rect 3564 2034 3582 2052
rect 3564 2052 3582 2070
rect 3564 2070 3582 2088
rect 3564 2088 3582 2106
rect 3564 2106 3582 2124
rect 3564 2124 3582 2142
rect 3564 2142 3582 2160
rect 3564 2160 3582 2178
rect 3564 2178 3582 2196
rect 3564 2196 3582 2214
rect 3564 2214 3582 2232
rect 3564 2232 3582 2250
rect 3564 2250 3582 2268
rect 3564 2268 3582 2286
rect 3564 2286 3582 2304
rect 3564 2304 3582 2322
rect 3564 2322 3582 2340
rect 3564 2340 3582 2358
rect 3564 2358 3582 2376
rect 3564 2376 3582 2394
rect 3564 2394 3582 2412
rect 3564 2412 3582 2430
rect 3564 2700 3582 2718
rect 3564 2718 3582 2736
rect 3564 2736 3582 2754
rect 3564 2754 3582 2772
rect 3564 2772 3582 2790
rect 3564 2790 3582 2808
rect 3564 2808 3582 2826
rect 3564 2826 3582 2844
rect 3564 2844 3582 2862
rect 3564 2862 3582 2880
rect 3564 2880 3582 2898
rect 3564 2898 3582 2916
rect 3564 2916 3582 2934
rect 3564 2934 3582 2952
rect 3564 2952 3582 2970
rect 3564 2970 3582 2988
rect 3564 2988 3582 3006
rect 3564 3006 3582 3024
rect 3564 3024 3582 3042
rect 3564 3042 3582 3060
rect 3564 3060 3582 3078
rect 3564 3078 3582 3096
rect 3564 3096 3582 3114
rect 3564 3114 3582 3132
rect 3564 3132 3582 3150
rect 3564 3150 3582 3168
rect 3564 3168 3582 3186
rect 3564 3186 3582 3204
rect 3564 3204 3582 3222
rect 3564 3222 3582 3240
rect 3564 3240 3582 3258
rect 3564 3258 3582 3276
rect 3564 3276 3582 3294
rect 3564 3294 3582 3312
rect 3564 3312 3582 3330
rect 3564 3330 3582 3348
rect 3564 3348 3582 3366
rect 3564 3366 3582 3384
rect 3564 3384 3582 3402
rect 3564 3402 3582 3420
rect 3564 3420 3582 3438
rect 3564 3438 3582 3456
rect 3564 3456 3582 3474
rect 3564 3474 3582 3492
rect 3564 3492 3582 3510
rect 3564 3510 3582 3528
rect 3564 3528 3582 3546
rect 3564 3546 3582 3564
rect 3564 3564 3582 3582
rect 3564 3582 3582 3600
rect 3564 3600 3582 3618
rect 3564 3618 3582 3636
rect 3564 3636 3582 3654
rect 3564 3654 3582 3672
rect 3564 3672 3582 3690
rect 3564 3690 3582 3708
rect 3564 3708 3582 3726
rect 3564 3726 3582 3744
rect 3564 3744 3582 3762
rect 3564 3762 3582 3780
rect 3564 3780 3582 3798
rect 3564 3798 3582 3816
rect 3564 3816 3582 3834
rect 3564 3834 3582 3852
rect 3564 3852 3582 3870
rect 3564 3870 3582 3888
rect 3564 3888 3582 3906
rect 3564 3906 3582 3924
rect 3564 3924 3582 3942
rect 3564 3942 3582 3960
rect 3564 3960 3582 3978
rect 3564 3978 3582 3996
rect 3564 3996 3582 4014
rect 3564 4014 3582 4032
rect 3564 4032 3582 4050
rect 3564 4050 3582 4068
rect 3564 4068 3582 4086
rect 3564 4086 3582 4104
rect 3564 4104 3582 4122
rect 3564 4122 3582 4140
rect 3564 4140 3582 4158
rect 3564 4158 3582 4176
rect 3564 4176 3582 4194
rect 3564 4194 3582 4212
rect 3564 4212 3582 4230
rect 3564 4230 3582 4248
rect 3564 4248 3582 4266
rect 3564 4266 3582 4284
rect 3564 4284 3582 4302
rect 3564 4302 3582 4320
rect 3564 4320 3582 4338
rect 3564 4338 3582 4356
rect 3564 4356 3582 4374
rect 3564 4374 3582 4392
rect 3564 4392 3582 4410
rect 3564 4410 3582 4428
rect 3564 4428 3582 4446
rect 3564 4446 3582 4464
rect 3564 4464 3582 4482
rect 3564 4482 3582 4500
rect 3564 4500 3582 4518
rect 3564 4518 3582 4536
rect 3564 4536 3582 4554
rect 3564 4554 3582 4572
rect 3564 4572 3582 4590
rect 3564 4590 3582 4608
rect 3564 4608 3582 4626
rect 3564 4626 3582 4644
rect 3564 4644 3582 4662
rect 3564 4662 3582 4680
rect 3564 4680 3582 4698
rect 3564 4698 3582 4716
rect 3564 4716 3582 4734
rect 3564 4734 3582 4752
rect 3564 4752 3582 4770
rect 3564 4770 3582 4788
rect 3564 4788 3582 4806
rect 3564 4806 3582 4824
rect 3564 4824 3582 4842
rect 3564 4842 3582 4860
rect 3564 4860 3582 4878
rect 3564 4878 3582 4896
rect 3564 4896 3582 4914
rect 3564 4914 3582 4932
rect 3564 4932 3582 4950
rect 3564 4950 3582 4968
rect 3564 4968 3582 4986
rect 3564 4986 3582 5004
rect 3564 5004 3582 5022
rect 3564 5022 3582 5040
rect 3564 5040 3582 5058
rect 3564 6642 3582 6660
rect 3564 6660 3582 6678
rect 3564 6678 3582 6696
rect 3564 6696 3582 6714
rect 3564 6714 3582 6732
rect 3564 6732 3582 6750
rect 3564 6750 3582 6768
rect 3564 6768 3582 6786
rect 3564 6786 3582 6804
rect 3564 6804 3582 6822
rect 3564 6822 3582 6840
rect 3564 6840 3582 6858
rect 3564 6858 3582 6876
rect 3564 6876 3582 6894
rect 3564 6894 3582 6912
rect 3564 6912 3582 6930
rect 3564 6930 3582 6948
rect 3564 6948 3582 6966
rect 3564 6966 3582 6984
rect 3564 6984 3582 7002
rect 3564 7002 3582 7020
rect 3564 7020 3582 7038
rect 3564 7038 3582 7056
rect 3564 7056 3582 7074
rect 3564 7074 3582 7092
rect 3564 7092 3582 7110
rect 3564 7110 3582 7128
rect 3564 7128 3582 7146
rect 3564 7146 3582 7164
rect 3564 7164 3582 7182
rect 3564 7182 3582 7200
rect 3564 7200 3582 7218
rect 3564 7218 3582 7236
rect 3564 7236 3582 7254
rect 3564 7254 3582 7272
rect 3582 18 3600 36
rect 3582 36 3600 54
rect 3582 54 3600 72
rect 3582 72 3600 90
rect 3582 90 3600 108
rect 3582 108 3600 126
rect 3582 126 3600 144
rect 3582 144 3600 162
rect 3582 162 3600 180
rect 3582 180 3600 198
rect 3582 198 3600 216
rect 3582 216 3600 234
rect 3582 234 3600 252
rect 3582 252 3600 270
rect 3582 270 3600 288
rect 3582 288 3600 306
rect 3582 306 3600 324
rect 3582 324 3600 342
rect 3582 342 3600 360
rect 3582 360 3600 378
rect 3582 378 3600 396
rect 3582 396 3600 414
rect 3582 414 3600 432
rect 3582 432 3600 450
rect 3582 450 3600 468
rect 3582 468 3600 486
rect 3582 486 3600 504
rect 3582 504 3600 522
rect 3582 522 3600 540
rect 3582 540 3600 558
rect 3582 558 3600 576
rect 3582 576 3600 594
rect 3582 594 3600 612
rect 3582 828 3600 846
rect 3582 846 3600 864
rect 3582 864 3600 882
rect 3582 882 3600 900
rect 3582 900 3600 918
rect 3582 918 3600 936
rect 3582 936 3600 954
rect 3582 954 3600 972
rect 3582 972 3600 990
rect 3582 990 3600 1008
rect 3582 1008 3600 1026
rect 3582 1026 3600 1044
rect 3582 1044 3600 1062
rect 3582 1062 3600 1080
rect 3582 1080 3600 1098
rect 3582 1098 3600 1116
rect 3582 1116 3600 1134
rect 3582 1134 3600 1152
rect 3582 1152 3600 1170
rect 3582 1170 3600 1188
rect 3582 1188 3600 1206
rect 3582 1206 3600 1224
rect 3582 1224 3600 1242
rect 3582 1242 3600 1260
rect 3582 1260 3600 1278
rect 3582 1494 3600 1512
rect 3582 1512 3600 1530
rect 3582 1530 3600 1548
rect 3582 1548 3600 1566
rect 3582 1566 3600 1584
rect 3582 1584 3600 1602
rect 3582 1602 3600 1620
rect 3582 1620 3600 1638
rect 3582 1638 3600 1656
rect 3582 1656 3600 1674
rect 3582 1674 3600 1692
rect 3582 1692 3600 1710
rect 3582 1710 3600 1728
rect 3582 1728 3600 1746
rect 3582 1746 3600 1764
rect 3582 1764 3600 1782
rect 3582 1782 3600 1800
rect 3582 1800 3600 1818
rect 3582 1818 3600 1836
rect 3582 1836 3600 1854
rect 3582 1854 3600 1872
rect 3582 1872 3600 1890
rect 3582 1890 3600 1908
rect 3582 1908 3600 1926
rect 3582 1926 3600 1944
rect 3582 1944 3600 1962
rect 3582 1962 3600 1980
rect 3582 1980 3600 1998
rect 3582 1998 3600 2016
rect 3582 2016 3600 2034
rect 3582 2034 3600 2052
rect 3582 2052 3600 2070
rect 3582 2070 3600 2088
rect 3582 2088 3600 2106
rect 3582 2106 3600 2124
rect 3582 2124 3600 2142
rect 3582 2142 3600 2160
rect 3582 2160 3600 2178
rect 3582 2178 3600 2196
rect 3582 2196 3600 2214
rect 3582 2214 3600 2232
rect 3582 2232 3600 2250
rect 3582 2250 3600 2268
rect 3582 2268 3600 2286
rect 3582 2286 3600 2304
rect 3582 2304 3600 2322
rect 3582 2322 3600 2340
rect 3582 2340 3600 2358
rect 3582 2358 3600 2376
rect 3582 2376 3600 2394
rect 3582 2394 3600 2412
rect 3582 2412 3600 2430
rect 3582 2430 3600 2448
rect 3582 2448 3600 2466
rect 3582 2718 3600 2736
rect 3582 2736 3600 2754
rect 3582 2754 3600 2772
rect 3582 2772 3600 2790
rect 3582 2790 3600 2808
rect 3582 2808 3600 2826
rect 3582 2826 3600 2844
rect 3582 2844 3600 2862
rect 3582 2862 3600 2880
rect 3582 2880 3600 2898
rect 3582 2898 3600 2916
rect 3582 2916 3600 2934
rect 3582 2934 3600 2952
rect 3582 2952 3600 2970
rect 3582 2970 3600 2988
rect 3582 2988 3600 3006
rect 3582 3006 3600 3024
rect 3582 3024 3600 3042
rect 3582 3042 3600 3060
rect 3582 3060 3600 3078
rect 3582 3078 3600 3096
rect 3582 3096 3600 3114
rect 3582 3114 3600 3132
rect 3582 3132 3600 3150
rect 3582 3150 3600 3168
rect 3582 3168 3600 3186
rect 3582 3186 3600 3204
rect 3582 3204 3600 3222
rect 3582 3222 3600 3240
rect 3582 3240 3600 3258
rect 3582 3258 3600 3276
rect 3582 3276 3600 3294
rect 3582 3294 3600 3312
rect 3582 3312 3600 3330
rect 3582 3330 3600 3348
rect 3582 3348 3600 3366
rect 3582 3366 3600 3384
rect 3582 3384 3600 3402
rect 3582 3402 3600 3420
rect 3582 3420 3600 3438
rect 3582 3438 3600 3456
rect 3582 3456 3600 3474
rect 3582 3474 3600 3492
rect 3582 3492 3600 3510
rect 3582 3510 3600 3528
rect 3582 3528 3600 3546
rect 3582 3546 3600 3564
rect 3582 3564 3600 3582
rect 3582 3582 3600 3600
rect 3582 3600 3600 3618
rect 3582 3618 3600 3636
rect 3582 3636 3600 3654
rect 3582 3654 3600 3672
rect 3582 3672 3600 3690
rect 3582 3690 3600 3708
rect 3582 3708 3600 3726
rect 3582 3726 3600 3744
rect 3582 3744 3600 3762
rect 3582 3762 3600 3780
rect 3582 3780 3600 3798
rect 3582 3798 3600 3816
rect 3582 3816 3600 3834
rect 3582 3834 3600 3852
rect 3582 3852 3600 3870
rect 3582 3870 3600 3888
rect 3582 3888 3600 3906
rect 3582 3906 3600 3924
rect 3582 3924 3600 3942
rect 3582 3942 3600 3960
rect 3582 3960 3600 3978
rect 3582 3978 3600 3996
rect 3582 3996 3600 4014
rect 3582 4014 3600 4032
rect 3582 4032 3600 4050
rect 3582 4050 3600 4068
rect 3582 4068 3600 4086
rect 3582 4086 3600 4104
rect 3582 4104 3600 4122
rect 3582 4122 3600 4140
rect 3582 4140 3600 4158
rect 3582 4158 3600 4176
rect 3582 4176 3600 4194
rect 3582 4194 3600 4212
rect 3582 4212 3600 4230
rect 3582 4230 3600 4248
rect 3582 4248 3600 4266
rect 3582 4266 3600 4284
rect 3582 4284 3600 4302
rect 3582 4302 3600 4320
rect 3582 4320 3600 4338
rect 3582 4338 3600 4356
rect 3582 4356 3600 4374
rect 3582 4374 3600 4392
rect 3582 4392 3600 4410
rect 3582 4410 3600 4428
rect 3582 4428 3600 4446
rect 3582 4446 3600 4464
rect 3582 4464 3600 4482
rect 3582 4482 3600 4500
rect 3582 4500 3600 4518
rect 3582 4518 3600 4536
rect 3582 4536 3600 4554
rect 3582 4554 3600 4572
rect 3582 4572 3600 4590
rect 3582 4590 3600 4608
rect 3582 4608 3600 4626
rect 3582 4626 3600 4644
rect 3582 4644 3600 4662
rect 3582 4662 3600 4680
rect 3582 4680 3600 4698
rect 3582 4698 3600 4716
rect 3582 4716 3600 4734
rect 3582 4734 3600 4752
rect 3582 4752 3600 4770
rect 3582 4770 3600 4788
rect 3582 4788 3600 4806
rect 3582 4806 3600 4824
rect 3582 4824 3600 4842
rect 3582 4842 3600 4860
rect 3582 4860 3600 4878
rect 3582 4878 3600 4896
rect 3582 4896 3600 4914
rect 3582 4914 3600 4932
rect 3582 4932 3600 4950
rect 3582 4950 3600 4968
rect 3582 4968 3600 4986
rect 3582 4986 3600 5004
rect 3582 5004 3600 5022
rect 3582 5022 3600 5040
rect 3582 5040 3600 5058
rect 3582 5058 3600 5076
rect 3582 5076 3600 5094
rect 3582 5094 3600 5112
rect 3582 6642 3600 6660
rect 3582 6660 3600 6678
rect 3582 6678 3600 6696
rect 3582 6696 3600 6714
rect 3582 6714 3600 6732
rect 3582 6732 3600 6750
rect 3582 6750 3600 6768
rect 3582 6768 3600 6786
rect 3582 6786 3600 6804
rect 3582 6804 3600 6822
rect 3582 6822 3600 6840
rect 3582 6840 3600 6858
rect 3582 6858 3600 6876
rect 3582 6876 3600 6894
rect 3582 6894 3600 6912
rect 3582 6912 3600 6930
rect 3582 6930 3600 6948
rect 3582 6948 3600 6966
rect 3582 6966 3600 6984
rect 3582 6984 3600 7002
rect 3582 7002 3600 7020
rect 3582 7020 3600 7038
rect 3582 7038 3600 7056
rect 3582 7056 3600 7074
rect 3582 7074 3600 7092
rect 3582 7092 3600 7110
rect 3582 7110 3600 7128
rect 3582 7128 3600 7146
rect 3582 7146 3600 7164
rect 3582 7164 3600 7182
rect 3582 7182 3600 7200
rect 3582 7200 3600 7218
rect 3582 7218 3600 7236
rect 3582 7236 3600 7254
rect 3582 7254 3600 7272
rect 3600 18 3618 36
rect 3600 36 3618 54
rect 3600 54 3618 72
rect 3600 72 3618 90
rect 3600 90 3618 108
rect 3600 108 3618 126
rect 3600 126 3618 144
rect 3600 144 3618 162
rect 3600 162 3618 180
rect 3600 180 3618 198
rect 3600 198 3618 216
rect 3600 216 3618 234
rect 3600 234 3618 252
rect 3600 252 3618 270
rect 3600 270 3618 288
rect 3600 288 3618 306
rect 3600 306 3618 324
rect 3600 324 3618 342
rect 3600 342 3618 360
rect 3600 360 3618 378
rect 3600 378 3618 396
rect 3600 396 3618 414
rect 3600 414 3618 432
rect 3600 432 3618 450
rect 3600 450 3618 468
rect 3600 468 3618 486
rect 3600 486 3618 504
rect 3600 504 3618 522
rect 3600 522 3618 540
rect 3600 540 3618 558
rect 3600 558 3618 576
rect 3600 576 3618 594
rect 3600 594 3618 612
rect 3600 846 3618 864
rect 3600 864 3618 882
rect 3600 882 3618 900
rect 3600 900 3618 918
rect 3600 918 3618 936
rect 3600 936 3618 954
rect 3600 954 3618 972
rect 3600 972 3618 990
rect 3600 990 3618 1008
rect 3600 1008 3618 1026
rect 3600 1026 3618 1044
rect 3600 1044 3618 1062
rect 3600 1062 3618 1080
rect 3600 1080 3618 1098
rect 3600 1098 3618 1116
rect 3600 1116 3618 1134
rect 3600 1134 3618 1152
rect 3600 1152 3618 1170
rect 3600 1170 3618 1188
rect 3600 1188 3618 1206
rect 3600 1206 3618 1224
rect 3600 1224 3618 1242
rect 3600 1242 3618 1260
rect 3600 1260 3618 1278
rect 3600 1278 3618 1296
rect 3600 1512 3618 1530
rect 3600 1530 3618 1548
rect 3600 1548 3618 1566
rect 3600 1566 3618 1584
rect 3600 1584 3618 1602
rect 3600 1602 3618 1620
rect 3600 1620 3618 1638
rect 3600 1638 3618 1656
rect 3600 1656 3618 1674
rect 3600 1674 3618 1692
rect 3600 1692 3618 1710
rect 3600 1710 3618 1728
rect 3600 1728 3618 1746
rect 3600 1746 3618 1764
rect 3600 1764 3618 1782
rect 3600 1782 3618 1800
rect 3600 1800 3618 1818
rect 3600 1818 3618 1836
rect 3600 1836 3618 1854
rect 3600 1854 3618 1872
rect 3600 1872 3618 1890
rect 3600 1890 3618 1908
rect 3600 1908 3618 1926
rect 3600 1926 3618 1944
rect 3600 1944 3618 1962
rect 3600 1962 3618 1980
rect 3600 1980 3618 1998
rect 3600 1998 3618 2016
rect 3600 2016 3618 2034
rect 3600 2034 3618 2052
rect 3600 2052 3618 2070
rect 3600 2070 3618 2088
rect 3600 2088 3618 2106
rect 3600 2106 3618 2124
rect 3600 2124 3618 2142
rect 3600 2142 3618 2160
rect 3600 2160 3618 2178
rect 3600 2178 3618 2196
rect 3600 2196 3618 2214
rect 3600 2214 3618 2232
rect 3600 2232 3618 2250
rect 3600 2250 3618 2268
rect 3600 2268 3618 2286
rect 3600 2286 3618 2304
rect 3600 2304 3618 2322
rect 3600 2322 3618 2340
rect 3600 2340 3618 2358
rect 3600 2358 3618 2376
rect 3600 2376 3618 2394
rect 3600 2394 3618 2412
rect 3600 2412 3618 2430
rect 3600 2430 3618 2448
rect 3600 2448 3618 2466
rect 3600 2466 3618 2484
rect 3600 2754 3618 2772
rect 3600 2772 3618 2790
rect 3600 2790 3618 2808
rect 3600 2808 3618 2826
rect 3600 2826 3618 2844
rect 3600 2844 3618 2862
rect 3600 2862 3618 2880
rect 3600 2880 3618 2898
rect 3600 2898 3618 2916
rect 3600 2916 3618 2934
rect 3600 2934 3618 2952
rect 3600 2952 3618 2970
rect 3600 2970 3618 2988
rect 3600 2988 3618 3006
rect 3600 3006 3618 3024
rect 3600 3024 3618 3042
rect 3600 3042 3618 3060
rect 3600 3060 3618 3078
rect 3600 3078 3618 3096
rect 3600 3096 3618 3114
rect 3600 3114 3618 3132
rect 3600 3132 3618 3150
rect 3600 3150 3618 3168
rect 3600 3168 3618 3186
rect 3600 3186 3618 3204
rect 3600 3204 3618 3222
rect 3600 3222 3618 3240
rect 3600 3240 3618 3258
rect 3600 3258 3618 3276
rect 3600 3276 3618 3294
rect 3600 3294 3618 3312
rect 3600 3312 3618 3330
rect 3600 3330 3618 3348
rect 3600 3348 3618 3366
rect 3600 3366 3618 3384
rect 3600 3384 3618 3402
rect 3600 3402 3618 3420
rect 3600 3420 3618 3438
rect 3600 3438 3618 3456
rect 3600 3456 3618 3474
rect 3600 3474 3618 3492
rect 3600 3492 3618 3510
rect 3600 3510 3618 3528
rect 3600 3528 3618 3546
rect 3600 3546 3618 3564
rect 3600 3564 3618 3582
rect 3600 3582 3618 3600
rect 3600 3600 3618 3618
rect 3600 3618 3618 3636
rect 3600 3636 3618 3654
rect 3600 3654 3618 3672
rect 3600 3672 3618 3690
rect 3600 3690 3618 3708
rect 3600 3708 3618 3726
rect 3600 3726 3618 3744
rect 3600 3744 3618 3762
rect 3600 3762 3618 3780
rect 3600 3780 3618 3798
rect 3600 3798 3618 3816
rect 3600 3816 3618 3834
rect 3600 3834 3618 3852
rect 3600 3852 3618 3870
rect 3600 3870 3618 3888
rect 3600 3888 3618 3906
rect 3600 3906 3618 3924
rect 3600 3924 3618 3942
rect 3600 3942 3618 3960
rect 3600 3960 3618 3978
rect 3600 3978 3618 3996
rect 3600 3996 3618 4014
rect 3600 4014 3618 4032
rect 3600 4032 3618 4050
rect 3600 4050 3618 4068
rect 3600 4068 3618 4086
rect 3600 4086 3618 4104
rect 3600 4104 3618 4122
rect 3600 4122 3618 4140
rect 3600 4140 3618 4158
rect 3600 4158 3618 4176
rect 3600 4176 3618 4194
rect 3600 4194 3618 4212
rect 3600 4212 3618 4230
rect 3600 4230 3618 4248
rect 3600 4248 3618 4266
rect 3600 4266 3618 4284
rect 3600 4284 3618 4302
rect 3600 4302 3618 4320
rect 3600 4320 3618 4338
rect 3600 4338 3618 4356
rect 3600 4356 3618 4374
rect 3600 4374 3618 4392
rect 3600 4392 3618 4410
rect 3600 4410 3618 4428
rect 3600 4428 3618 4446
rect 3600 4446 3618 4464
rect 3600 4464 3618 4482
rect 3600 4482 3618 4500
rect 3600 4500 3618 4518
rect 3600 4518 3618 4536
rect 3600 4536 3618 4554
rect 3600 4554 3618 4572
rect 3600 4572 3618 4590
rect 3600 4590 3618 4608
rect 3600 4608 3618 4626
rect 3600 4626 3618 4644
rect 3600 4644 3618 4662
rect 3600 4662 3618 4680
rect 3600 4680 3618 4698
rect 3600 4698 3618 4716
rect 3600 4716 3618 4734
rect 3600 4734 3618 4752
rect 3600 4752 3618 4770
rect 3600 4770 3618 4788
rect 3600 4788 3618 4806
rect 3600 4806 3618 4824
rect 3600 4824 3618 4842
rect 3600 4842 3618 4860
rect 3600 4860 3618 4878
rect 3600 4878 3618 4896
rect 3600 4896 3618 4914
rect 3600 4914 3618 4932
rect 3600 4932 3618 4950
rect 3600 4950 3618 4968
rect 3600 4968 3618 4986
rect 3600 4986 3618 5004
rect 3600 5004 3618 5022
rect 3600 5022 3618 5040
rect 3600 5040 3618 5058
rect 3600 5058 3618 5076
rect 3600 5076 3618 5094
rect 3600 5094 3618 5112
rect 3600 5112 3618 5130
rect 3600 5130 3618 5148
rect 3600 6642 3618 6660
rect 3600 6660 3618 6678
rect 3600 6678 3618 6696
rect 3600 6696 3618 6714
rect 3600 6714 3618 6732
rect 3600 6732 3618 6750
rect 3600 6750 3618 6768
rect 3600 6768 3618 6786
rect 3600 6786 3618 6804
rect 3600 6804 3618 6822
rect 3600 6822 3618 6840
rect 3600 6840 3618 6858
rect 3600 6858 3618 6876
rect 3600 6876 3618 6894
rect 3600 6894 3618 6912
rect 3600 6912 3618 6930
rect 3600 6930 3618 6948
rect 3600 6948 3618 6966
rect 3600 6966 3618 6984
rect 3600 6984 3618 7002
rect 3600 7002 3618 7020
rect 3600 7020 3618 7038
rect 3600 7038 3618 7056
rect 3600 7056 3618 7074
rect 3600 7074 3618 7092
rect 3600 7092 3618 7110
rect 3600 7110 3618 7128
rect 3600 7128 3618 7146
rect 3600 7146 3618 7164
rect 3600 7164 3618 7182
rect 3600 7182 3618 7200
rect 3600 7200 3618 7218
rect 3600 7218 3618 7236
rect 3600 7236 3618 7254
rect 3600 7254 3618 7272
rect 3618 18 3636 36
rect 3618 36 3636 54
rect 3618 54 3636 72
rect 3618 72 3636 90
rect 3618 90 3636 108
rect 3618 108 3636 126
rect 3618 126 3636 144
rect 3618 144 3636 162
rect 3618 162 3636 180
rect 3618 180 3636 198
rect 3618 198 3636 216
rect 3618 216 3636 234
rect 3618 234 3636 252
rect 3618 252 3636 270
rect 3618 270 3636 288
rect 3618 288 3636 306
rect 3618 306 3636 324
rect 3618 324 3636 342
rect 3618 342 3636 360
rect 3618 360 3636 378
rect 3618 378 3636 396
rect 3618 396 3636 414
rect 3618 414 3636 432
rect 3618 432 3636 450
rect 3618 450 3636 468
rect 3618 468 3636 486
rect 3618 486 3636 504
rect 3618 504 3636 522
rect 3618 522 3636 540
rect 3618 540 3636 558
rect 3618 558 3636 576
rect 3618 576 3636 594
rect 3618 594 3636 612
rect 3618 846 3636 864
rect 3618 864 3636 882
rect 3618 882 3636 900
rect 3618 900 3636 918
rect 3618 918 3636 936
rect 3618 936 3636 954
rect 3618 954 3636 972
rect 3618 972 3636 990
rect 3618 990 3636 1008
rect 3618 1008 3636 1026
rect 3618 1026 3636 1044
rect 3618 1044 3636 1062
rect 3618 1062 3636 1080
rect 3618 1080 3636 1098
rect 3618 1098 3636 1116
rect 3618 1116 3636 1134
rect 3618 1134 3636 1152
rect 3618 1152 3636 1170
rect 3618 1170 3636 1188
rect 3618 1188 3636 1206
rect 3618 1206 3636 1224
rect 3618 1224 3636 1242
rect 3618 1242 3636 1260
rect 3618 1260 3636 1278
rect 3618 1278 3636 1296
rect 3618 1296 3636 1314
rect 3618 1530 3636 1548
rect 3618 1548 3636 1566
rect 3618 1566 3636 1584
rect 3618 1584 3636 1602
rect 3618 1602 3636 1620
rect 3618 1620 3636 1638
rect 3618 1638 3636 1656
rect 3618 1656 3636 1674
rect 3618 1674 3636 1692
rect 3618 1692 3636 1710
rect 3618 1710 3636 1728
rect 3618 1728 3636 1746
rect 3618 1746 3636 1764
rect 3618 1764 3636 1782
rect 3618 1782 3636 1800
rect 3618 1800 3636 1818
rect 3618 1818 3636 1836
rect 3618 1836 3636 1854
rect 3618 1854 3636 1872
rect 3618 1872 3636 1890
rect 3618 1890 3636 1908
rect 3618 1908 3636 1926
rect 3618 1926 3636 1944
rect 3618 1944 3636 1962
rect 3618 1962 3636 1980
rect 3618 1980 3636 1998
rect 3618 1998 3636 2016
rect 3618 2016 3636 2034
rect 3618 2034 3636 2052
rect 3618 2052 3636 2070
rect 3618 2070 3636 2088
rect 3618 2088 3636 2106
rect 3618 2106 3636 2124
rect 3618 2124 3636 2142
rect 3618 2142 3636 2160
rect 3618 2160 3636 2178
rect 3618 2178 3636 2196
rect 3618 2196 3636 2214
rect 3618 2214 3636 2232
rect 3618 2232 3636 2250
rect 3618 2250 3636 2268
rect 3618 2268 3636 2286
rect 3618 2286 3636 2304
rect 3618 2304 3636 2322
rect 3618 2322 3636 2340
rect 3618 2340 3636 2358
rect 3618 2358 3636 2376
rect 3618 2376 3636 2394
rect 3618 2394 3636 2412
rect 3618 2412 3636 2430
rect 3618 2430 3636 2448
rect 3618 2448 3636 2466
rect 3618 2466 3636 2484
rect 3618 2484 3636 2502
rect 3618 2502 3636 2520
rect 3618 2772 3636 2790
rect 3618 2790 3636 2808
rect 3618 2808 3636 2826
rect 3618 2826 3636 2844
rect 3618 2844 3636 2862
rect 3618 2862 3636 2880
rect 3618 2880 3636 2898
rect 3618 2898 3636 2916
rect 3618 2916 3636 2934
rect 3618 2934 3636 2952
rect 3618 2952 3636 2970
rect 3618 2970 3636 2988
rect 3618 2988 3636 3006
rect 3618 3006 3636 3024
rect 3618 3024 3636 3042
rect 3618 3042 3636 3060
rect 3618 3060 3636 3078
rect 3618 3078 3636 3096
rect 3618 3096 3636 3114
rect 3618 3114 3636 3132
rect 3618 3132 3636 3150
rect 3618 3150 3636 3168
rect 3618 3168 3636 3186
rect 3618 3186 3636 3204
rect 3618 3204 3636 3222
rect 3618 3222 3636 3240
rect 3618 3240 3636 3258
rect 3618 3258 3636 3276
rect 3618 3276 3636 3294
rect 3618 3294 3636 3312
rect 3618 3312 3636 3330
rect 3618 3330 3636 3348
rect 3618 3348 3636 3366
rect 3618 3366 3636 3384
rect 3618 3384 3636 3402
rect 3618 3402 3636 3420
rect 3618 3420 3636 3438
rect 3618 3438 3636 3456
rect 3618 3456 3636 3474
rect 3618 3474 3636 3492
rect 3618 3492 3636 3510
rect 3618 3510 3636 3528
rect 3618 3528 3636 3546
rect 3618 3546 3636 3564
rect 3618 3564 3636 3582
rect 3618 3582 3636 3600
rect 3618 3600 3636 3618
rect 3618 3618 3636 3636
rect 3618 3636 3636 3654
rect 3618 3654 3636 3672
rect 3618 3672 3636 3690
rect 3618 3690 3636 3708
rect 3618 3708 3636 3726
rect 3618 3726 3636 3744
rect 3618 3744 3636 3762
rect 3618 3762 3636 3780
rect 3618 3780 3636 3798
rect 3618 3798 3636 3816
rect 3618 3816 3636 3834
rect 3618 3834 3636 3852
rect 3618 3852 3636 3870
rect 3618 3870 3636 3888
rect 3618 3888 3636 3906
rect 3618 3906 3636 3924
rect 3618 3924 3636 3942
rect 3618 3942 3636 3960
rect 3618 3960 3636 3978
rect 3618 3978 3636 3996
rect 3618 3996 3636 4014
rect 3618 4014 3636 4032
rect 3618 4032 3636 4050
rect 3618 4050 3636 4068
rect 3618 4068 3636 4086
rect 3618 4086 3636 4104
rect 3618 4104 3636 4122
rect 3618 4122 3636 4140
rect 3618 4140 3636 4158
rect 3618 4158 3636 4176
rect 3618 4176 3636 4194
rect 3618 4194 3636 4212
rect 3618 4212 3636 4230
rect 3618 4230 3636 4248
rect 3618 4248 3636 4266
rect 3618 4266 3636 4284
rect 3618 4284 3636 4302
rect 3618 4302 3636 4320
rect 3618 4320 3636 4338
rect 3618 4338 3636 4356
rect 3618 4356 3636 4374
rect 3618 4374 3636 4392
rect 3618 4392 3636 4410
rect 3618 4410 3636 4428
rect 3618 4428 3636 4446
rect 3618 4446 3636 4464
rect 3618 4464 3636 4482
rect 3618 4482 3636 4500
rect 3618 4500 3636 4518
rect 3618 4518 3636 4536
rect 3618 4536 3636 4554
rect 3618 4554 3636 4572
rect 3618 4572 3636 4590
rect 3618 4590 3636 4608
rect 3618 4608 3636 4626
rect 3618 4626 3636 4644
rect 3618 4644 3636 4662
rect 3618 4662 3636 4680
rect 3618 4680 3636 4698
rect 3618 4698 3636 4716
rect 3618 4716 3636 4734
rect 3618 4734 3636 4752
rect 3618 4752 3636 4770
rect 3618 4770 3636 4788
rect 3618 4788 3636 4806
rect 3618 4806 3636 4824
rect 3618 4824 3636 4842
rect 3618 4842 3636 4860
rect 3618 4860 3636 4878
rect 3618 4878 3636 4896
rect 3618 4896 3636 4914
rect 3618 4914 3636 4932
rect 3618 4932 3636 4950
rect 3618 4950 3636 4968
rect 3618 4968 3636 4986
rect 3618 4986 3636 5004
rect 3618 5004 3636 5022
rect 3618 5022 3636 5040
rect 3618 5040 3636 5058
rect 3618 5058 3636 5076
rect 3618 5076 3636 5094
rect 3618 5094 3636 5112
rect 3618 5112 3636 5130
rect 3618 5130 3636 5148
rect 3618 5148 3636 5166
rect 3618 5166 3636 5184
rect 3618 5184 3636 5202
rect 3618 6642 3636 6660
rect 3618 6660 3636 6678
rect 3618 6678 3636 6696
rect 3618 6696 3636 6714
rect 3618 6714 3636 6732
rect 3618 6732 3636 6750
rect 3618 6750 3636 6768
rect 3618 6768 3636 6786
rect 3618 6786 3636 6804
rect 3618 6804 3636 6822
rect 3618 6822 3636 6840
rect 3618 6840 3636 6858
rect 3618 6858 3636 6876
rect 3618 6876 3636 6894
rect 3618 6894 3636 6912
rect 3618 6912 3636 6930
rect 3618 6930 3636 6948
rect 3618 6948 3636 6966
rect 3618 6966 3636 6984
rect 3618 6984 3636 7002
rect 3618 7002 3636 7020
rect 3618 7020 3636 7038
rect 3618 7038 3636 7056
rect 3618 7056 3636 7074
rect 3618 7074 3636 7092
rect 3618 7092 3636 7110
rect 3618 7110 3636 7128
rect 3618 7128 3636 7146
rect 3618 7146 3636 7164
rect 3618 7164 3636 7182
rect 3618 7182 3636 7200
rect 3618 7200 3636 7218
rect 3618 7218 3636 7236
rect 3618 7236 3636 7254
rect 3618 7254 3636 7272
rect 3636 0 3654 18
rect 3636 18 3654 36
rect 3636 36 3654 54
rect 3636 54 3654 72
rect 3636 72 3654 90
rect 3636 90 3654 108
rect 3636 108 3654 126
rect 3636 126 3654 144
rect 3636 144 3654 162
rect 3636 162 3654 180
rect 3636 180 3654 198
rect 3636 198 3654 216
rect 3636 216 3654 234
rect 3636 234 3654 252
rect 3636 252 3654 270
rect 3636 270 3654 288
rect 3636 288 3654 306
rect 3636 306 3654 324
rect 3636 324 3654 342
rect 3636 342 3654 360
rect 3636 360 3654 378
rect 3636 378 3654 396
rect 3636 396 3654 414
rect 3636 414 3654 432
rect 3636 432 3654 450
rect 3636 450 3654 468
rect 3636 468 3654 486
rect 3636 486 3654 504
rect 3636 504 3654 522
rect 3636 522 3654 540
rect 3636 540 3654 558
rect 3636 558 3654 576
rect 3636 576 3654 594
rect 3636 594 3654 612
rect 3636 846 3654 864
rect 3636 864 3654 882
rect 3636 882 3654 900
rect 3636 900 3654 918
rect 3636 918 3654 936
rect 3636 936 3654 954
rect 3636 954 3654 972
rect 3636 972 3654 990
rect 3636 990 3654 1008
rect 3636 1008 3654 1026
rect 3636 1026 3654 1044
rect 3636 1044 3654 1062
rect 3636 1062 3654 1080
rect 3636 1080 3654 1098
rect 3636 1098 3654 1116
rect 3636 1116 3654 1134
rect 3636 1134 3654 1152
rect 3636 1152 3654 1170
rect 3636 1170 3654 1188
rect 3636 1188 3654 1206
rect 3636 1206 3654 1224
rect 3636 1224 3654 1242
rect 3636 1242 3654 1260
rect 3636 1260 3654 1278
rect 3636 1278 3654 1296
rect 3636 1296 3654 1314
rect 3636 1530 3654 1548
rect 3636 1548 3654 1566
rect 3636 1566 3654 1584
rect 3636 1584 3654 1602
rect 3636 1602 3654 1620
rect 3636 1620 3654 1638
rect 3636 1638 3654 1656
rect 3636 1656 3654 1674
rect 3636 1674 3654 1692
rect 3636 1692 3654 1710
rect 3636 1710 3654 1728
rect 3636 1728 3654 1746
rect 3636 1746 3654 1764
rect 3636 1764 3654 1782
rect 3636 1782 3654 1800
rect 3636 1800 3654 1818
rect 3636 1818 3654 1836
rect 3636 1836 3654 1854
rect 3636 1854 3654 1872
rect 3636 1872 3654 1890
rect 3636 1890 3654 1908
rect 3636 1908 3654 1926
rect 3636 1926 3654 1944
rect 3636 1944 3654 1962
rect 3636 1962 3654 1980
rect 3636 1980 3654 1998
rect 3636 1998 3654 2016
rect 3636 2016 3654 2034
rect 3636 2034 3654 2052
rect 3636 2052 3654 2070
rect 3636 2070 3654 2088
rect 3636 2088 3654 2106
rect 3636 2106 3654 2124
rect 3636 2124 3654 2142
rect 3636 2142 3654 2160
rect 3636 2160 3654 2178
rect 3636 2178 3654 2196
rect 3636 2196 3654 2214
rect 3636 2214 3654 2232
rect 3636 2232 3654 2250
rect 3636 2250 3654 2268
rect 3636 2268 3654 2286
rect 3636 2286 3654 2304
rect 3636 2304 3654 2322
rect 3636 2322 3654 2340
rect 3636 2340 3654 2358
rect 3636 2358 3654 2376
rect 3636 2376 3654 2394
rect 3636 2394 3654 2412
rect 3636 2412 3654 2430
rect 3636 2430 3654 2448
rect 3636 2448 3654 2466
rect 3636 2466 3654 2484
rect 3636 2484 3654 2502
rect 3636 2502 3654 2520
rect 3636 2520 3654 2538
rect 3636 2808 3654 2826
rect 3636 2826 3654 2844
rect 3636 2844 3654 2862
rect 3636 2862 3654 2880
rect 3636 2880 3654 2898
rect 3636 2898 3654 2916
rect 3636 2916 3654 2934
rect 3636 2934 3654 2952
rect 3636 2952 3654 2970
rect 3636 2970 3654 2988
rect 3636 2988 3654 3006
rect 3636 3006 3654 3024
rect 3636 3024 3654 3042
rect 3636 3042 3654 3060
rect 3636 3060 3654 3078
rect 3636 3078 3654 3096
rect 3636 3096 3654 3114
rect 3636 3114 3654 3132
rect 3636 3132 3654 3150
rect 3636 3150 3654 3168
rect 3636 3168 3654 3186
rect 3636 3186 3654 3204
rect 3636 3204 3654 3222
rect 3636 3222 3654 3240
rect 3636 3240 3654 3258
rect 3636 3258 3654 3276
rect 3636 3276 3654 3294
rect 3636 3294 3654 3312
rect 3636 3312 3654 3330
rect 3636 3330 3654 3348
rect 3636 3348 3654 3366
rect 3636 3366 3654 3384
rect 3636 3384 3654 3402
rect 3636 3402 3654 3420
rect 3636 3420 3654 3438
rect 3636 3438 3654 3456
rect 3636 3456 3654 3474
rect 3636 3474 3654 3492
rect 3636 3492 3654 3510
rect 3636 3510 3654 3528
rect 3636 3528 3654 3546
rect 3636 3546 3654 3564
rect 3636 3564 3654 3582
rect 3636 3582 3654 3600
rect 3636 3600 3654 3618
rect 3636 3618 3654 3636
rect 3636 3636 3654 3654
rect 3636 3654 3654 3672
rect 3636 3672 3654 3690
rect 3636 3690 3654 3708
rect 3636 3708 3654 3726
rect 3636 3726 3654 3744
rect 3636 3744 3654 3762
rect 3636 3762 3654 3780
rect 3636 3780 3654 3798
rect 3636 3798 3654 3816
rect 3636 3816 3654 3834
rect 3636 3834 3654 3852
rect 3636 3852 3654 3870
rect 3636 3870 3654 3888
rect 3636 3888 3654 3906
rect 3636 3906 3654 3924
rect 3636 3924 3654 3942
rect 3636 3942 3654 3960
rect 3636 3960 3654 3978
rect 3636 3978 3654 3996
rect 3636 3996 3654 4014
rect 3636 4014 3654 4032
rect 3636 4032 3654 4050
rect 3636 4050 3654 4068
rect 3636 4068 3654 4086
rect 3636 4086 3654 4104
rect 3636 4104 3654 4122
rect 3636 4122 3654 4140
rect 3636 4140 3654 4158
rect 3636 4158 3654 4176
rect 3636 4176 3654 4194
rect 3636 4194 3654 4212
rect 3636 4212 3654 4230
rect 3636 4230 3654 4248
rect 3636 4248 3654 4266
rect 3636 4266 3654 4284
rect 3636 4284 3654 4302
rect 3636 4302 3654 4320
rect 3636 4320 3654 4338
rect 3636 4338 3654 4356
rect 3636 4356 3654 4374
rect 3636 4374 3654 4392
rect 3636 4392 3654 4410
rect 3636 4410 3654 4428
rect 3636 4428 3654 4446
rect 3636 4446 3654 4464
rect 3636 4464 3654 4482
rect 3636 4482 3654 4500
rect 3636 4500 3654 4518
rect 3636 4518 3654 4536
rect 3636 4536 3654 4554
rect 3636 4554 3654 4572
rect 3636 4572 3654 4590
rect 3636 4590 3654 4608
rect 3636 4608 3654 4626
rect 3636 4626 3654 4644
rect 3636 4644 3654 4662
rect 3636 4662 3654 4680
rect 3636 4680 3654 4698
rect 3636 4698 3654 4716
rect 3636 4716 3654 4734
rect 3636 4734 3654 4752
rect 3636 4752 3654 4770
rect 3636 4770 3654 4788
rect 3636 4788 3654 4806
rect 3636 4806 3654 4824
rect 3636 4824 3654 4842
rect 3636 4842 3654 4860
rect 3636 4860 3654 4878
rect 3636 4878 3654 4896
rect 3636 4896 3654 4914
rect 3636 4914 3654 4932
rect 3636 4932 3654 4950
rect 3636 4950 3654 4968
rect 3636 4968 3654 4986
rect 3636 4986 3654 5004
rect 3636 5004 3654 5022
rect 3636 5022 3654 5040
rect 3636 5040 3654 5058
rect 3636 5058 3654 5076
rect 3636 5076 3654 5094
rect 3636 5094 3654 5112
rect 3636 5112 3654 5130
rect 3636 5130 3654 5148
rect 3636 5148 3654 5166
rect 3636 5166 3654 5184
rect 3636 5184 3654 5202
rect 3636 5202 3654 5220
rect 3636 5220 3654 5238
rect 3636 6642 3654 6660
rect 3636 6660 3654 6678
rect 3636 6678 3654 6696
rect 3636 6696 3654 6714
rect 3636 6714 3654 6732
rect 3636 6732 3654 6750
rect 3636 6750 3654 6768
rect 3636 6768 3654 6786
rect 3636 6786 3654 6804
rect 3636 6804 3654 6822
rect 3636 6822 3654 6840
rect 3636 6840 3654 6858
rect 3636 6858 3654 6876
rect 3636 6876 3654 6894
rect 3636 6894 3654 6912
rect 3636 6912 3654 6930
rect 3636 6930 3654 6948
rect 3636 6948 3654 6966
rect 3636 6966 3654 6984
rect 3636 6984 3654 7002
rect 3636 7002 3654 7020
rect 3636 7020 3654 7038
rect 3636 7038 3654 7056
rect 3636 7056 3654 7074
rect 3636 7074 3654 7092
rect 3636 7092 3654 7110
rect 3636 7110 3654 7128
rect 3636 7128 3654 7146
rect 3636 7146 3654 7164
rect 3636 7164 3654 7182
rect 3636 7182 3654 7200
rect 3636 7200 3654 7218
rect 3636 7218 3654 7236
rect 3636 7236 3654 7254
rect 3636 7254 3654 7272
rect 3654 0 3672 18
rect 3654 18 3672 36
rect 3654 36 3672 54
rect 3654 54 3672 72
rect 3654 72 3672 90
rect 3654 90 3672 108
rect 3654 108 3672 126
rect 3654 126 3672 144
rect 3654 144 3672 162
rect 3654 162 3672 180
rect 3654 180 3672 198
rect 3654 198 3672 216
rect 3654 216 3672 234
rect 3654 234 3672 252
rect 3654 252 3672 270
rect 3654 270 3672 288
rect 3654 288 3672 306
rect 3654 306 3672 324
rect 3654 324 3672 342
rect 3654 342 3672 360
rect 3654 360 3672 378
rect 3654 378 3672 396
rect 3654 396 3672 414
rect 3654 414 3672 432
rect 3654 432 3672 450
rect 3654 450 3672 468
rect 3654 468 3672 486
rect 3654 486 3672 504
rect 3654 504 3672 522
rect 3654 522 3672 540
rect 3654 540 3672 558
rect 3654 558 3672 576
rect 3654 576 3672 594
rect 3654 594 3672 612
rect 3654 846 3672 864
rect 3654 864 3672 882
rect 3654 882 3672 900
rect 3654 900 3672 918
rect 3654 918 3672 936
rect 3654 936 3672 954
rect 3654 954 3672 972
rect 3654 972 3672 990
rect 3654 990 3672 1008
rect 3654 1008 3672 1026
rect 3654 1026 3672 1044
rect 3654 1044 3672 1062
rect 3654 1062 3672 1080
rect 3654 1080 3672 1098
rect 3654 1098 3672 1116
rect 3654 1116 3672 1134
rect 3654 1134 3672 1152
rect 3654 1152 3672 1170
rect 3654 1170 3672 1188
rect 3654 1188 3672 1206
rect 3654 1206 3672 1224
rect 3654 1224 3672 1242
rect 3654 1242 3672 1260
rect 3654 1260 3672 1278
rect 3654 1278 3672 1296
rect 3654 1296 3672 1314
rect 3654 1314 3672 1332
rect 3654 1548 3672 1566
rect 3654 1566 3672 1584
rect 3654 1584 3672 1602
rect 3654 1602 3672 1620
rect 3654 1620 3672 1638
rect 3654 1638 3672 1656
rect 3654 1656 3672 1674
rect 3654 1674 3672 1692
rect 3654 1692 3672 1710
rect 3654 1710 3672 1728
rect 3654 1728 3672 1746
rect 3654 1746 3672 1764
rect 3654 1764 3672 1782
rect 3654 1782 3672 1800
rect 3654 1800 3672 1818
rect 3654 1818 3672 1836
rect 3654 1836 3672 1854
rect 3654 1854 3672 1872
rect 3654 1872 3672 1890
rect 3654 1890 3672 1908
rect 3654 1908 3672 1926
rect 3654 1926 3672 1944
rect 3654 1944 3672 1962
rect 3654 1962 3672 1980
rect 3654 1980 3672 1998
rect 3654 1998 3672 2016
rect 3654 2016 3672 2034
rect 3654 2034 3672 2052
rect 3654 2052 3672 2070
rect 3654 2070 3672 2088
rect 3654 2088 3672 2106
rect 3654 2106 3672 2124
rect 3654 2124 3672 2142
rect 3654 2142 3672 2160
rect 3654 2160 3672 2178
rect 3654 2178 3672 2196
rect 3654 2196 3672 2214
rect 3654 2214 3672 2232
rect 3654 2232 3672 2250
rect 3654 2250 3672 2268
rect 3654 2268 3672 2286
rect 3654 2286 3672 2304
rect 3654 2304 3672 2322
rect 3654 2322 3672 2340
rect 3654 2340 3672 2358
rect 3654 2358 3672 2376
rect 3654 2376 3672 2394
rect 3654 2394 3672 2412
rect 3654 2412 3672 2430
rect 3654 2430 3672 2448
rect 3654 2448 3672 2466
rect 3654 2466 3672 2484
rect 3654 2484 3672 2502
rect 3654 2502 3672 2520
rect 3654 2520 3672 2538
rect 3654 2538 3672 2556
rect 3654 2556 3672 2574
rect 3654 2826 3672 2844
rect 3654 2844 3672 2862
rect 3654 2862 3672 2880
rect 3654 2880 3672 2898
rect 3654 2898 3672 2916
rect 3654 2916 3672 2934
rect 3654 2934 3672 2952
rect 3654 2952 3672 2970
rect 3654 2970 3672 2988
rect 3654 2988 3672 3006
rect 3654 3006 3672 3024
rect 3654 3024 3672 3042
rect 3654 3042 3672 3060
rect 3654 3060 3672 3078
rect 3654 3078 3672 3096
rect 3654 3096 3672 3114
rect 3654 3114 3672 3132
rect 3654 3132 3672 3150
rect 3654 3150 3672 3168
rect 3654 3168 3672 3186
rect 3654 3186 3672 3204
rect 3654 3204 3672 3222
rect 3654 3222 3672 3240
rect 3654 3240 3672 3258
rect 3654 3258 3672 3276
rect 3654 3276 3672 3294
rect 3654 3294 3672 3312
rect 3654 3312 3672 3330
rect 3654 3330 3672 3348
rect 3654 3348 3672 3366
rect 3654 3366 3672 3384
rect 3654 3384 3672 3402
rect 3654 3402 3672 3420
rect 3654 3420 3672 3438
rect 3654 3438 3672 3456
rect 3654 3456 3672 3474
rect 3654 3474 3672 3492
rect 3654 3492 3672 3510
rect 3654 3510 3672 3528
rect 3654 3528 3672 3546
rect 3654 3546 3672 3564
rect 3654 3564 3672 3582
rect 3654 3582 3672 3600
rect 3654 3600 3672 3618
rect 3654 3618 3672 3636
rect 3654 3636 3672 3654
rect 3654 3654 3672 3672
rect 3654 3672 3672 3690
rect 3654 3690 3672 3708
rect 3654 3708 3672 3726
rect 3654 3726 3672 3744
rect 3654 3744 3672 3762
rect 3654 3762 3672 3780
rect 3654 3780 3672 3798
rect 3654 3798 3672 3816
rect 3654 3816 3672 3834
rect 3654 3834 3672 3852
rect 3654 3852 3672 3870
rect 3654 3870 3672 3888
rect 3654 3888 3672 3906
rect 3654 3906 3672 3924
rect 3654 3924 3672 3942
rect 3654 3942 3672 3960
rect 3654 3960 3672 3978
rect 3654 3978 3672 3996
rect 3654 3996 3672 4014
rect 3654 4014 3672 4032
rect 3654 4032 3672 4050
rect 3654 4050 3672 4068
rect 3654 4068 3672 4086
rect 3654 4086 3672 4104
rect 3654 4104 3672 4122
rect 3654 4122 3672 4140
rect 3654 4140 3672 4158
rect 3654 4158 3672 4176
rect 3654 4176 3672 4194
rect 3654 4194 3672 4212
rect 3654 4212 3672 4230
rect 3654 4230 3672 4248
rect 3654 4248 3672 4266
rect 3654 4266 3672 4284
rect 3654 4284 3672 4302
rect 3654 4302 3672 4320
rect 3654 4320 3672 4338
rect 3654 4338 3672 4356
rect 3654 4356 3672 4374
rect 3654 4374 3672 4392
rect 3654 4392 3672 4410
rect 3654 4410 3672 4428
rect 3654 4428 3672 4446
rect 3654 4446 3672 4464
rect 3654 4464 3672 4482
rect 3654 4482 3672 4500
rect 3654 4500 3672 4518
rect 3654 4518 3672 4536
rect 3654 4536 3672 4554
rect 3654 4554 3672 4572
rect 3654 4572 3672 4590
rect 3654 4590 3672 4608
rect 3654 4608 3672 4626
rect 3654 4626 3672 4644
rect 3654 4644 3672 4662
rect 3654 4662 3672 4680
rect 3654 4680 3672 4698
rect 3654 4698 3672 4716
rect 3654 4716 3672 4734
rect 3654 4734 3672 4752
rect 3654 4752 3672 4770
rect 3654 4770 3672 4788
rect 3654 4788 3672 4806
rect 3654 4806 3672 4824
rect 3654 4824 3672 4842
rect 3654 4842 3672 4860
rect 3654 4860 3672 4878
rect 3654 4878 3672 4896
rect 3654 4896 3672 4914
rect 3654 4914 3672 4932
rect 3654 4932 3672 4950
rect 3654 4950 3672 4968
rect 3654 4968 3672 4986
rect 3654 4986 3672 5004
rect 3654 5004 3672 5022
rect 3654 5022 3672 5040
rect 3654 5040 3672 5058
rect 3654 5058 3672 5076
rect 3654 5076 3672 5094
rect 3654 5094 3672 5112
rect 3654 5112 3672 5130
rect 3654 5130 3672 5148
rect 3654 5148 3672 5166
rect 3654 5166 3672 5184
rect 3654 5184 3672 5202
rect 3654 5202 3672 5220
rect 3654 5220 3672 5238
rect 3654 5238 3672 5256
rect 3654 5256 3672 5274
rect 3654 5274 3672 5292
rect 3654 6642 3672 6660
rect 3654 6660 3672 6678
rect 3654 6678 3672 6696
rect 3654 6696 3672 6714
rect 3654 6714 3672 6732
rect 3654 6732 3672 6750
rect 3654 6750 3672 6768
rect 3654 6768 3672 6786
rect 3654 6786 3672 6804
rect 3654 6804 3672 6822
rect 3654 6822 3672 6840
rect 3654 6840 3672 6858
rect 3654 6858 3672 6876
rect 3654 6876 3672 6894
rect 3654 6894 3672 6912
rect 3654 6912 3672 6930
rect 3654 6930 3672 6948
rect 3654 6948 3672 6966
rect 3654 6966 3672 6984
rect 3654 6984 3672 7002
rect 3654 7002 3672 7020
rect 3654 7020 3672 7038
rect 3654 7038 3672 7056
rect 3654 7056 3672 7074
rect 3654 7074 3672 7092
rect 3654 7092 3672 7110
rect 3654 7110 3672 7128
rect 3654 7128 3672 7146
rect 3654 7146 3672 7164
rect 3654 7164 3672 7182
rect 3654 7182 3672 7200
rect 3654 7200 3672 7218
rect 3654 7218 3672 7236
rect 3654 7236 3672 7254
rect 3654 7254 3672 7272
rect 3672 0 3690 18
rect 3672 18 3690 36
rect 3672 36 3690 54
rect 3672 54 3690 72
rect 3672 72 3690 90
rect 3672 90 3690 108
rect 3672 108 3690 126
rect 3672 126 3690 144
rect 3672 144 3690 162
rect 3672 162 3690 180
rect 3672 180 3690 198
rect 3672 198 3690 216
rect 3672 216 3690 234
rect 3672 234 3690 252
rect 3672 252 3690 270
rect 3672 270 3690 288
rect 3672 288 3690 306
rect 3672 306 3690 324
rect 3672 324 3690 342
rect 3672 342 3690 360
rect 3672 360 3690 378
rect 3672 378 3690 396
rect 3672 396 3690 414
rect 3672 414 3690 432
rect 3672 432 3690 450
rect 3672 450 3690 468
rect 3672 468 3690 486
rect 3672 486 3690 504
rect 3672 504 3690 522
rect 3672 522 3690 540
rect 3672 540 3690 558
rect 3672 558 3690 576
rect 3672 576 3690 594
rect 3672 594 3690 612
rect 3672 846 3690 864
rect 3672 864 3690 882
rect 3672 882 3690 900
rect 3672 900 3690 918
rect 3672 918 3690 936
rect 3672 936 3690 954
rect 3672 954 3690 972
rect 3672 972 3690 990
rect 3672 990 3690 1008
rect 3672 1008 3690 1026
rect 3672 1026 3690 1044
rect 3672 1044 3690 1062
rect 3672 1062 3690 1080
rect 3672 1080 3690 1098
rect 3672 1098 3690 1116
rect 3672 1116 3690 1134
rect 3672 1134 3690 1152
rect 3672 1152 3690 1170
rect 3672 1170 3690 1188
rect 3672 1188 3690 1206
rect 3672 1206 3690 1224
rect 3672 1224 3690 1242
rect 3672 1242 3690 1260
rect 3672 1260 3690 1278
rect 3672 1278 3690 1296
rect 3672 1296 3690 1314
rect 3672 1314 3690 1332
rect 3672 1332 3690 1350
rect 3672 1566 3690 1584
rect 3672 1584 3690 1602
rect 3672 1602 3690 1620
rect 3672 1620 3690 1638
rect 3672 1638 3690 1656
rect 3672 1656 3690 1674
rect 3672 1674 3690 1692
rect 3672 1692 3690 1710
rect 3672 1710 3690 1728
rect 3672 1728 3690 1746
rect 3672 1746 3690 1764
rect 3672 1764 3690 1782
rect 3672 1782 3690 1800
rect 3672 1800 3690 1818
rect 3672 1818 3690 1836
rect 3672 1836 3690 1854
rect 3672 1854 3690 1872
rect 3672 1872 3690 1890
rect 3672 1890 3690 1908
rect 3672 1908 3690 1926
rect 3672 1926 3690 1944
rect 3672 1944 3690 1962
rect 3672 1962 3690 1980
rect 3672 1980 3690 1998
rect 3672 1998 3690 2016
rect 3672 2016 3690 2034
rect 3672 2034 3690 2052
rect 3672 2052 3690 2070
rect 3672 2070 3690 2088
rect 3672 2088 3690 2106
rect 3672 2106 3690 2124
rect 3672 2124 3690 2142
rect 3672 2142 3690 2160
rect 3672 2160 3690 2178
rect 3672 2178 3690 2196
rect 3672 2196 3690 2214
rect 3672 2214 3690 2232
rect 3672 2232 3690 2250
rect 3672 2250 3690 2268
rect 3672 2268 3690 2286
rect 3672 2286 3690 2304
rect 3672 2304 3690 2322
rect 3672 2322 3690 2340
rect 3672 2340 3690 2358
rect 3672 2358 3690 2376
rect 3672 2376 3690 2394
rect 3672 2394 3690 2412
rect 3672 2412 3690 2430
rect 3672 2430 3690 2448
rect 3672 2448 3690 2466
rect 3672 2466 3690 2484
rect 3672 2484 3690 2502
rect 3672 2502 3690 2520
rect 3672 2520 3690 2538
rect 3672 2538 3690 2556
rect 3672 2556 3690 2574
rect 3672 2574 3690 2592
rect 3672 2592 3690 2610
rect 3672 2862 3690 2880
rect 3672 2880 3690 2898
rect 3672 2898 3690 2916
rect 3672 2916 3690 2934
rect 3672 2934 3690 2952
rect 3672 2952 3690 2970
rect 3672 2970 3690 2988
rect 3672 2988 3690 3006
rect 3672 3006 3690 3024
rect 3672 3024 3690 3042
rect 3672 3042 3690 3060
rect 3672 3060 3690 3078
rect 3672 3078 3690 3096
rect 3672 3096 3690 3114
rect 3672 3114 3690 3132
rect 3672 3132 3690 3150
rect 3672 3150 3690 3168
rect 3672 3168 3690 3186
rect 3672 3186 3690 3204
rect 3672 3204 3690 3222
rect 3672 3222 3690 3240
rect 3672 3240 3690 3258
rect 3672 3258 3690 3276
rect 3672 3276 3690 3294
rect 3672 3294 3690 3312
rect 3672 3312 3690 3330
rect 3672 3330 3690 3348
rect 3672 3348 3690 3366
rect 3672 3366 3690 3384
rect 3672 3384 3690 3402
rect 3672 3402 3690 3420
rect 3672 3420 3690 3438
rect 3672 3438 3690 3456
rect 3672 3456 3690 3474
rect 3672 3474 3690 3492
rect 3672 3492 3690 3510
rect 3672 3510 3690 3528
rect 3672 3528 3690 3546
rect 3672 3546 3690 3564
rect 3672 3564 3690 3582
rect 3672 3582 3690 3600
rect 3672 3600 3690 3618
rect 3672 3618 3690 3636
rect 3672 3636 3690 3654
rect 3672 3654 3690 3672
rect 3672 3672 3690 3690
rect 3672 3690 3690 3708
rect 3672 3708 3690 3726
rect 3672 3726 3690 3744
rect 3672 3744 3690 3762
rect 3672 3762 3690 3780
rect 3672 3780 3690 3798
rect 3672 3798 3690 3816
rect 3672 3816 3690 3834
rect 3672 3834 3690 3852
rect 3672 3852 3690 3870
rect 3672 3870 3690 3888
rect 3672 3888 3690 3906
rect 3672 3906 3690 3924
rect 3672 3924 3690 3942
rect 3672 3942 3690 3960
rect 3672 3960 3690 3978
rect 3672 3978 3690 3996
rect 3672 3996 3690 4014
rect 3672 4014 3690 4032
rect 3672 4032 3690 4050
rect 3672 4050 3690 4068
rect 3672 4068 3690 4086
rect 3672 4086 3690 4104
rect 3672 4104 3690 4122
rect 3672 4122 3690 4140
rect 3672 4140 3690 4158
rect 3672 4158 3690 4176
rect 3672 4176 3690 4194
rect 3672 4194 3690 4212
rect 3672 4212 3690 4230
rect 3672 4230 3690 4248
rect 3672 4248 3690 4266
rect 3672 4266 3690 4284
rect 3672 4284 3690 4302
rect 3672 4302 3690 4320
rect 3672 4320 3690 4338
rect 3672 4338 3690 4356
rect 3672 4356 3690 4374
rect 3672 4374 3690 4392
rect 3672 4392 3690 4410
rect 3672 4410 3690 4428
rect 3672 4428 3690 4446
rect 3672 4446 3690 4464
rect 3672 4464 3690 4482
rect 3672 4482 3690 4500
rect 3672 4500 3690 4518
rect 3672 4518 3690 4536
rect 3672 4536 3690 4554
rect 3672 4554 3690 4572
rect 3672 4572 3690 4590
rect 3672 4590 3690 4608
rect 3672 4608 3690 4626
rect 3672 4626 3690 4644
rect 3672 4644 3690 4662
rect 3672 4662 3690 4680
rect 3672 4680 3690 4698
rect 3672 4698 3690 4716
rect 3672 4716 3690 4734
rect 3672 4734 3690 4752
rect 3672 4752 3690 4770
rect 3672 4770 3690 4788
rect 3672 4788 3690 4806
rect 3672 4806 3690 4824
rect 3672 4824 3690 4842
rect 3672 4842 3690 4860
rect 3672 4860 3690 4878
rect 3672 4878 3690 4896
rect 3672 4896 3690 4914
rect 3672 4914 3690 4932
rect 3672 4932 3690 4950
rect 3672 4950 3690 4968
rect 3672 4968 3690 4986
rect 3672 4986 3690 5004
rect 3672 5004 3690 5022
rect 3672 5022 3690 5040
rect 3672 5040 3690 5058
rect 3672 5058 3690 5076
rect 3672 5076 3690 5094
rect 3672 5094 3690 5112
rect 3672 5112 3690 5130
rect 3672 5130 3690 5148
rect 3672 5148 3690 5166
rect 3672 5166 3690 5184
rect 3672 5184 3690 5202
rect 3672 5202 3690 5220
rect 3672 5220 3690 5238
rect 3672 5238 3690 5256
rect 3672 5256 3690 5274
rect 3672 5274 3690 5292
rect 3672 5292 3690 5310
rect 3672 5310 3690 5328
rect 3672 6642 3690 6660
rect 3672 6660 3690 6678
rect 3672 6678 3690 6696
rect 3672 6696 3690 6714
rect 3672 6714 3690 6732
rect 3672 6732 3690 6750
rect 3672 6750 3690 6768
rect 3672 6768 3690 6786
rect 3672 6786 3690 6804
rect 3672 6804 3690 6822
rect 3672 6822 3690 6840
rect 3672 6840 3690 6858
rect 3672 6858 3690 6876
rect 3672 6876 3690 6894
rect 3672 6894 3690 6912
rect 3672 6912 3690 6930
rect 3672 6930 3690 6948
rect 3672 6948 3690 6966
rect 3672 6966 3690 6984
rect 3672 6984 3690 7002
rect 3672 7002 3690 7020
rect 3672 7020 3690 7038
rect 3672 7038 3690 7056
rect 3672 7056 3690 7074
rect 3672 7074 3690 7092
rect 3672 7092 3690 7110
rect 3672 7110 3690 7128
rect 3672 7128 3690 7146
rect 3672 7146 3690 7164
rect 3672 7164 3690 7182
rect 3672 7182 3690 7200
rect 3672 7200 3690 7218
rect 3672 7218 3690 7236
rect 3672 7236 3690 7254
rect 3672 7254 3690 7272
rect 3690 0 3708 18
rect 3690 18 3708 36
rect 3690 36 3708 54
rect 3690 54 3708 72
rect 3690 72 3708 90
rect 3690 90 3708 108
rect 3690 108 3708 126
rect 3690 126 3708 144
rect 3690 144 3708 162
rect 3690 162 3708 180
rect 3690 180 3708 198
rect 3690 198 3708 216
rect 3690 216 3708 234
rect 3690 234 3708 252
rect 3690 252 3708 270
rect 3690 270 3708 288
rect 3690 288 3708 306
rect 3690 306 3708 324
rect 3690 324 3708 342
rect 3690 342 3708 360
rect 3690 360 3708 378
rect 3690 378 3708 396
rect 3690 396 3708 414
rect 3690 414 3708 432
rect 3690 432 3708 450
rect 3690 450 3708 468
rect 3690 468 3708 486
rect 3690 486 3708 504
rect 3690 504 3708 522
rect 3690 522 3708 540
rect 3690 540 3708 558
rect 3690 558 3708 576
rect 3690 576 3708 594
rect 3690 594 3708 612
rect 3690 846 3708 864
rect 3690 864 3708 882
rect 3690 882 3708 900
rect 3690 900 3708 918
rect 3690 918 3708 936
rect 3690 936 3708 954
rect 3690 954 3708 972
rect 3690 972 3708 990
rect 3690 990 3708 1008
rect 3690 1008 3708 1026
rect 3690 1026 3708 1044
rect 3690 1044 3708 1062
rect 3690 1062 3708 1080
rect 3690 1080 3708 1098
rect 3690 1098 3708 1116
rect 3690 1116 3708 1134
rect 3690 1134 3708 1152
rect 3690 1152 3708 1170
rect 3690 1170 3708 1188
rect 3690 1188 3708 1206
rect 3690 1206 3708 1224
rect 3690 1224 3708 1242
rect 3690 1242 3708 1260
rect 3690 1260 3708 1278
rect 3690 1278 3708 1296
rect 3690 1296 3708 1314
rect 3690 1314 3708 1332
rect 3690 1332 3708 1350
rect 3690 1584 3708 1602
rect 3690 1602 3708 1620
rect 3690 1620 3708 1638
rect 3690 1638 3708 1656
rect 3690 1656 3708 1674
rect 3690 1674 3708 1692
rect 3690 1692 3708 1710
rect 3690 1710 3708 1728
rect 3690 1728 3708 1746
rect 3690 1746 3708 1764
rect 3690 1764 3708 1782
rect 3690 1782 3708 1800
rect 3690 1800 3708 1818
rect 3690 1818 3708 1836
rect 3690 1836 3708 1854
rect 3690 1854 3708 1872
rect 3690 1872 3708 1890
rect 3690 1890 3708 1908
rect 3690 1908 3708 1926
rect 3690 1926 3708 1944
rect 3690 1944 3708 1962
rect 3690 1962 3708 1980
rect 3690 1980 3708 1998
rect 3690 1998 3708 2016
rect 3690 2016 3708 2034
rect 3690 2034 3708 2052
rect 3690 2052 3708 2070
rect 3690 2070 3708 2088
rect 3690 2088 3708 2106
rect 3690 2106 3708 2124
rect 3690 2124 3708 2142
rect 3690 2142 3708 2160
rect 3690 2160 3708 2178
rect 3690 2178 3708 2196
rect 3690 2196 3708 2214
rect 3690 2214 3708 2232
rect 3690 2232 3708 2250
rect 3690 2250 3708 2268
rect 3690 2268 3708 2286
rect 3690 2286 3708 2304
rect 3690 2304 3708 2322
rect 3690 2322 3708 2340
rect 3690 2340 3708 2358
rect 3690 2358 3708 2376
rect 3690 2376 3708 2394
rect 3690 2394 3708 2412
rect 3690 2412 3708 2430
rect 3690 2430 3708 2448
rect 3690 2448 3708 2466
rect 3690 2466 3708 2484
rect 3690 2484 3708 2502
rect 3690 2502 3708 2520
rect 3690 2520 3708 2538
rect 3690 2538 3708 2556
rect 3690 2556 3708 2574
rect 3690 2574 3708 2592
rect 3690 2592 3708 2610
rect 3690 2610 3708 2628
rect 3690 2880 3708 2898
rect 3690 2898 3708 2916
rect 3690 2916 3708 2934
rect 3690 2934 3708 2952
rect 3690 2952 3708 2970
rect 3690 2970 3708 2988
rect 3690 2988 3708 3006
rect 3690 3006 3708 3024
rect 3690 3024 3708 3042
rect 3690 3042 3708 3060
rect 3690 3060 3708 3078
rect 3690 3078 3708 3096
rect 3690 3096 3708 3114
rect 3690 3114 3708 3132
rect 3690 3132 3708 3150
rect 3690 3150 3708 3168
rect 3690 3168 3708 3186
rect 3690 3186 3708 3204
rect 3690 3204 3708 3222
rect 3690 3222 3708 3240
rect 3690 3240 3708 3258
rect 3690 3258 3708 3276
rect 3690 3276 3708 3294
rect 3690 3294 3708 3312
rect 3690 3312 3708 3330
rect 3690 3330 3708 3348
rect 3690 3348 3708 3366
rect 3690 3366 3708 3384
rect 3690 3384 3708 3402
rect 3690 3402 3708 3420
rect 3690 3420 3708 3438
rect 3690 3438 3708 3456
rect 3690 3456 3708 3474
rect 3690 3474 3708 3492
rect 3690 3492 3708 3510
rect 3690 3510 3708 3528
rect 3690 3528 3708 3546
rect 3690 3546 3708 3564
rect 3690 3564 3708 3582
rect 3690 3582 3708 3600
rect 3690 3600 3708 3618
rect 3690 3618 3708 3636
rect 3690 3636 3708 3654
rect 3690 3654 3708 3672
rect 3690 3672 3708 3690
rect 3690 3690 3708 3708
rect 3690 3708 3708 3726
rect 3690 3726 3708 3744
rect 3690 3744 3708 3762
rect 3690 3762 3708 3780
rect 3690 3780 3708 3798
rect 3690 3798 3708 3816
rect 3690 3816 3708 3834
rect 3690 3834 3708 3852
rect 3690 3852 3708 3870
rect 3690 3870 3708 3888
rect 3690 3888 3708 3906
rect 3690 3906 3708 3924
rect 3690 3924 3708 3942
rect 3690 3942 3708 3960
rect 3690 3960 3708 3978
rect 3690 3978 3708 3996
rect 3690 3996 3708 4014
rect 3690 4014 3708 4032
rect 3690 4032 3708 4050
rect 3690 4050 3708 4068
rect 3690 4068 3708 4086
rect 3690 4086 3708 4104
rect 3690 4104 3708 4122
rect 3690 4122 3708 4140
rect 3690 4140 3708 4158
rect 3690 4158 3708 4176
rect 3690 4176 3708 4194
rect 3690 4194 3708 4212
rect 3690 4212 3708 4230
rect 3690 4230 3708 4248
rect 3690 4248 3708 4266
rect 3690 4266 3708 4284
rect 3690 4284 3708 4302
rect 3690 4302 3708 4320
rect 3690 4320 3708 4338
rect 3690 4338 3708 4356
rect 3690 4356 3708 4374
rect 3690 4374 3708 4392
rect 3690 4392 3708 4410
rect 3690 4410 3708 4428
rect 3690 4428 3708 4446
rect 3690 4446 3708 4464
rect 3690 4464 3708 4482
rect 3690 4482 3708 4500
rect 3690 4500 3708 4518
rect 3690 4518 3708 4536
rect 3690 4536 3708 4554
rect 3690 4554 3708 4572
rect 3690 4572 3708 4590
rect 3690 4590 3708 4608
rect 3690 4608 3708 4626
rect 3690 4626 3708 4644
rect 3690 4644 3708 4662
rect 3690 4662 3708 4680
rect 3690 4680 3708 4698
rect 3690 4698 3708 4716
rect 3690 4716 3708 4734
rect 3690 4734 3708 4752
rect 3690 4752 3708 4770
rect 3690 4770 3708 4788
rect 3690 4788 3708 4806
rect 3690 4806 3708 4824
rect 3690 4824 3708 4842
rect 3690 4842 3708 4860
rect 3690 4860 3708 4878
rect 3690 4878 3708 4896
rect 3690 4896 3708 4914
rect 3690 4914 3708 4932
rect 3690 4932 3708 4950
rect 3690 4950 3708 4968
rect 3690 4968 3708 4986
rect 3690 4986 3708 5004
rect 3690 5004 3708 5022
rect 3690 5022 3708 5040
rect 3690 5040 3708 5058
rect 3690 5058 3708 5076
rect 3690 5076 3708 5094
rect 3690 5094 3708 5112
rect 3690 5112 3708 5130
rect 3690 5130 3708 5148
rect 3690 5148 3708 5166
rect 3690 5166 3708 5184
rect 3690 5184 3708 5202
rect 3690 5202 3708 5220
rect 3690 5220 3708 5238
rect 3690 5238 3708 5256
rect 3690 5256 3708 5274
rect 3690 5274 3708 5292
rect 3690 5292 3708 5310
rect 3690 5310 3708 5328
rect 3690 5328 3708 5346
rect 3690 5346 3708 5364
rect 3690 5364 3708 5382
rect 3690 6642 3708 6660
rect 3690 6660 3708 6678
rect 3690 6678 3708 6696
rect 3690 6696 3708 6714
rect 3690 6714 3708 6732
rect 3690 6732 3708 6750
rect 3690 6750 3708 6768
rect 3690 6768 3708 6786
rect 3690 6786 3708 6804
rect 3690 6804 3708 6822
rect 3690 6822 3708 6840
rect 3690 6840 3708 6858
rect 3690 6858 3708 6876
rect 3690 6876 3708 6894
rect 3690 6894 3708 6912
rect 3690 6912 3708 6930
rect 3690 6930 3708 6948
rect 3690 6948 3708 6966
rect 3690 6966 3708 6984
rect 3690 6984 3708 7002
rect 3690 7002 3708 7020
rect 3690 7020 3708 7038
rect 3690 7038 3708 7056
rect 3690 7056 3708 7074
rect 3690 7074 3708 7092
rect 3690 7092 3708 7110
rect 3690 7110 3708 7128
rect 3690 7128 3708 7146
rect 3690 7146 3708 7164
rect 3690 7164 3708 7182
rect 3690 7182 3708 7200
rect 3690 7200 3708 7218
rect 3690 7218 3708 7236
rect 3690 7236 3708 7254
rect 3690 7254 3708 7272
rect 3708 0 3726 18
rect 3708 18 3726 36
rect 3708 36 3726 54
rect 3708 54 3726 72
rect 3708 72 3726 90
rect 3708 90 3726 108
rect 3708 108 3726 126
rect 3708 126 3726 144
rect 3708 144 3726 162
rect 3708 162 3726 180
rect 3708 180 3726 198
rect 3708 198 3726 216
rect 3708 216 3726 234
rect 3708 234 3726 252
rect 3708 252 3726 270
rect 3708 270 3726 288
rect 3708 288 3726 306
rect 3708 306 3726 324
rect 3708 324 3726 342
rect 3708 342 3726 360
rect 3708 360 3726 378
rect 3708 378 3726 396
rect 3708 396 3726 414
rect 3708 414 3726 432
rect 3708 432 3726 450
rect 3708 450 3726 468
rect 3708 468 3726 486
rect 3708 486 3726 504
rect 3708 504 3726 522
rect 3708 522 3726 540
rect 3708 540 3726 558
rect 3708 558 3726 576
rect 3708 576 3726 594
rect 3708 594 3726 612
rect 3708 846 3726 864
rect 3708 864 3726 882
rect 3708 882 3726 900
rect 3708 900 3726 918
rect 3708 918 3726 936
rect 3708 936 3726 954
rect 3708 954 3726 972
rect 3708 972 3726 990
rect 3708 990 3726 1008
rect 3708 1008 3726 1026
rect 3708 1026 3726 1044
rect 3708 1044 3726 1062
rect 3708 1062 3726 1080
rect 3708 1080 3726 1098
rect 3708 1098 3726 1116
rect 3708 1116 3726 1134
rect 3708 1134 3726 1152
rect 3708 1152 3726 1170
rect 3708 1170 3726 1188
rect 3708 1188 3726 1206
rect 3708 1206 3726 1224
rect 3708 1224 3726 1242
rect 3708 1242 3726 1260
rect 3708 1260 3726 1278
rect 3708 1278 3726 1296
rect 3708 1296 3726 1314
rect 3708 1314 3726 1332
rect 3708 1332 3726 1350
rect 3708 1350 3726 1368
rect 3708 1584 3726 1602
rect 3708 1602 3726 1620
rect 3708 1620 3726 1638
rect 3708 1638 3726 1656
rect 3708 1656 3726 1674
rect 3708 1674 3726 1692
rect 3708 1692 3726 1710
rect 3708 1710 3726 1728
rect 3708 1728 3726 1746
rect 3708 1746 3726 1764
rect 3708 1764 3726 1782
rect 3708 1782 3726 1800
rect 3708 1800 3726 1818
rect 3708 1818 3726 1836
rect 3708 1836 3726 1854
rect 3708 1854 3726 1872
rect 3708 1872 3726 1890
rect 3708 1890 3726 1908
rect 3708 1908 3726 1926
rect 3708 1926 3726 1944
rect 3708 1944 3726 1962
rect 3708 1962 3726 1980
rect 3708 1980 3726 1998
rect 3708 1998 3726 2016
rect 3708 2016 3726 2034
rect 3708 2034 3726 2052
rect 3708 2052 3726 2070
rect 3708 2070 3726 2088
rect 3708 2088 3726 2106
rect 3708 2106 3726 2124
rect 3708 2124 3726 2142
rect 3708 2142 3726 2160
rect 3708 2160 3726 2178
rect 3708 2178 3726 2196
rect 3708 2196 3726 2214
rect 3708 2214 3726 2232
rect 3708 2232 3726 2250
rect 3708 2250 3726 2268
rect 3708 2268 3726 2286
rect 3708 2286 3726 2304
rect 3708 2304 3726 2322
rect 3708 2322 3726 2340
rect 3708 2340 3726 2358
rect 3708 2358 3726 2376
rect 3708 2376 3726 2394
rect 3708 2394 3726 2412
rect 3708 2412 3726 2430
rect 3708 2430 3726 2448
rect 3708 2448 3726 2466
rect 3708 2466 3726 2484
rect 3708 2484 3726 2502
rect 3708 2502 3726 2520
rect 3708 2520 3726 2538
rect 3708 2538 3726 2556
rect 3708 2556 3726 2574
rect 3708 2574 3726 2592
rect 3708 2592 3726 2610
rect 3708 2610 3726 2628
rect 3708 2628 3726 2646
rect 3708 2646 3726 2664
rect 3708 2916 3726 2934
rect 3708 2934 3726 2952
rect 3708 2952 3726 2970
rect 3708 2970 3726 2988
rect 3708 2988 3726 3006
rect 3708 3006 3726 3024
rect 3708 3024 3726 3042
rect 3708 3042 3726 3060
rect 3708 3060 3726 3078
rect 3708 3078 3726 3096
rect 3708 3096 3726 3114
rect 3708 3114 3726 3132
rect 3708 3132 3726 3150
rect 3708 3150 3726 3168
rect 3708 3168 3726 3186
rect 3708 3186 3726 3204
rect 3708 3204 3726 3222
rect 3708 3222 3726 3240
rect 3708 3240 3726 3258
rect 3708 3258 3726 3276
rect 3708 3276 3726 3294
rect 3708 3294 3726 3312
rect 3708 3312 3726 3330
rect 3708 3330 3726 3348
rect 3708 3348 3726 3366
rect 3708 3366 3726 3384
rect 3708 3384 3726 3402
rect 3708 3402 3726 3420
rect 3708 3420 3726 3438
rect 3708 3438 3726 3456
rect 3708 3456 3726 3474
rect 3708 3474 3726 3492
rect 3708 3492 3726 3510
rect 3708 3510 3726 3528
rect 3708 3528 3726 3546
rect 3708 3546 3726 3564
rect 3708 3564 3726 3582
rect 3708 3582 3726 3600
rect 3708 3600 3726 3618
rect 3708 3618 3726 3636
rect 3708 3636 3726 3654
rect 3708 3654 3726 3672
rect 3708 3672 3726 3690
rect 3708 3690 3726 3708
rect 3708 3708 3726 3726
rect 3708 3726 3726 3744
rect 3708 3744 3726 3762
rect 3708 3762 3726 3780
rect 3708 3780 3726 3798
rect 3708 3798 3726 3816
rect 3708 3816 3726 3834
rect 3708 3834 3726 3852
rect 3708 3852 3726 3870
rect 3708 3870 3726 3888
rect 3708 3888 3726 3906
rect 3708 3906 3726 3924
rect 3708 3924 3726 3942
rect 3708 3942 3726 3960
rect 3708 3960 3726 3978
rect 3708 3978 3726 3996
rect 3708 3996 3726 4014
rect 3708 4014 3726 4032
rect 3708 4032 3726 4050
rect 3708 4050 3726 4068
rect 3708 4068 3726 4086
rect 3708 4086 3726 4104
rect 3708 4104 3726 4122
rect 3708 4122 3726 4140
rect 3708 4140 3726 4158
rect 3708 4158 3726 4176
rect 3708 4176 3726 4194
rect 3708 4194 3726 4212
rect 3708 4212 3726 4230
rect 3708 4230 3726 4248
rect 3708 4248 3726 4266
rect 3708 4266 3726 4284
rect 3708 4284 3726 4302
rect 3708 4302 3726 4320
rect 3708 4320 3726 4338
rect 3708 4338 3726 4356
rect 3708 4356 3726 4374
rect 3708 4374 3726 4392
rect 3708 4392 3726 4410
rect 3708 4410 3726 4428
rect 3708 4428 3726 4446
rect 3708 4446 3726 4464
rect 3708 4464 3726 4482
rect 3708 4482 3726 4500
rect 3708 4500 3726 4518
rect 3708 4518 3726 4536
rect 3708 4536 3726 4554
rect 3708 4554 3726 4572
rect 3708 4572 3726 4590
rect 3708 4590 3726 4608
rect 3708 4608 3726 4626
rect 3708 4626 3726 4644
rect 3708 4644 3726 4662
rect 3708 4662 3726 4680
rect 3708 4680 3726 4698
rect 3708 4698 3726 4716
rect 3708 4716 3726 4734
rect 3708 4734 3726 4752
rect 3708 4752 3726 4770
rect 3708 4770 3726 4788
rect 3708 4788 3726 4806
rect 3708 4806 3726 4824
rect 3708 4824 3726 4842
rect 3708 4842 3726 4860
rect 3708 4860 3726 4878
rect 3708 4878 3726 4896
rect 3708 4896 3726 4914
rect 3708 4914 3726 4932
rect 3708 4932 3726 4950
rect 3708 4950 3726 4968
rect 3708 4968 3726 4986
rect 3708 4986 3726 5004
rect 3708 5004 3726 5022
rect 3708 5022 3726 5040
rect 3708 5040 3726 5058
rect 3708 5058 3726 5076
rect 3708 5076 3726 5094
rect 3708 5094 3726 5112
rect 3708 5112 3726 5130
rect 3708 5130 3726 5148
rect 3708 5148 3726 5166
rect 3708 5166 3726 5184
rect 3708 5184 3726 5202
rect 3708 5202 3726 5220
rect 3708 5220 3726 5238
rect 3708 5238 3726 5256
rect 3708 5256 3726 5274
rect 3708 5274 3726 5292
rect 3708 5292 3726 5310
rect 3708 5310 3726 5328
rect 3708 5328 3726 5346
rect 3708 5346 3726 5364
rect 3708 5364 3726 5382
rect 3708 5382 3726 5400
rect 3708 5400 3726 5418
rect 3708 6642 3726 6660
rect 3708 6660 3726 6678
rect 3708 6678 3726 6696
rect 3708 6696 3726 6714
rect 3708 6714 3726 6732
rect 3708 6732 3726 6750
rect 3708 6750 3726 6768
rect 3708 6768 3726 6786
rect 3708 6786 3726 6804
rect 3708 6804 3726 6822
rect 3708 6822 3726 6840
rect 3708 6840 3726 6858
rect 3708 6858 3726 6876
rect 3708 6876 3726 6894
rect 3708 6894 3726 6912
rect 3708 6912 3726 6930
rect 3708 6930 3726 6948
rect 3708 6948 3726 6966
rect 3708 6966 3726 6984
rect 3708 6984 3726 7002
rect 3708 7002 3726 7020
rect 3708 7020 3726 7038
rect 3708 7038 3726 7056
rect 3708 7056 3726 7074
rect 3708 7074 3726 7092
rect 3708 7092 3726 7110
rect 3708 7110 3726 7128
rect 3708 7128 3726 7146
rect 3708 7146 3726 7164
rect 3708 7164 3726 7182
rect 3708 7182 3726 7200
rect 3708 7200 3726 7218
rect 3708 7218 3726 7236
rect 3708 7236 3726 7254
rect 3708 7254 3726 7272
rect 3726 0 3744 18
rect 3726 18 3744 36
rect 3726 36 3744 54
rect 3726 54 3744 72
rect 3726 72 3744 90
rect 3726 90 3744 108
rect 3726 108 3744 126
rect 3726 126 3744 144
rect 3726 144 3744 162
rect 3726 162 3744 180
rect 3726 180 3744 198
rect 3726 198 3744 216
rect 3726 216 3744 234
rect 3726 234 3744 252
rect 3726 252 3744 270
rect 3726 270 3744 288
rect 3726 288 3744 306
rect 3726 306 3744 324
rect 3726 324 3744 342
rect 3726 342 3744 360
rect 3726 360 3744 378
rect 3726 378 3744 396
rect 3726 396 3744 414
rect 3726 414 3744 432
rect 3726 432 3744 450
rect 3726 450 3744 468
rect 3726 468 3744 486
rect 3726 486 3744 504
rect 3726 504 3744 522
rect 3726 522 3744 540
rect 3726 540 3744 558
rect 3726 558 3744 576
rect 3726 576 3744 594
rect 3726 594 3744 612
rect 3726 612 3744 630
rect 3726 864 3744 882
rect 3726 882 3744 900
rect 3726 900 3744 918
rect 3726 918 3744 936
rect 3726 936 3744 954
rect 3726 954 3744 972
rect 3726 972 3744 990
rect 3726 990 3744 1008
rect 3726 1008 3744 1026
rect 3726 1026 3744 1044
rect 3726 1044 3744 1062
rect 3726 1062 3744 1080
rect 3726 1080 3744 1098
rect 3726 1098 3744 1116
rect 3726 1116 3744 1134
rect 3726 1134 3744 1152
rect 3726 1152 3744 1170
rect 3726 1170 3744 1188
rect 3726 1188 3744 1206
rect 3726 1206 3744 1224
rect 3726 1224 3744 1242
rect 3726 1242 3744 1260
rect 3726 1260 3744 1278
rect 3726 1278 3744 1296
rect 3726 1296 3744 1314
rect 3726 1314 3744 1332
rect 3726 1332 3744 1350
rect 3726 1350 3744 1368
rect 3726 1368 3744 1386
rect 3726 1602 3744 1620
rect 3726 1620 3744 1638
rect 3726 1638 3744 1656
rect 3726 1656 3744 1674
rect 3726 1674 3744 1692
rect 3726 1692 3744 1710
rect 3726 1710 3744 1728
rect 3726 1728 3744 1746
rect 3726 1746 3744 1764
rect 3726 1764 3744 1782
rect 3726 1782 3744 1800
rect 3726 1800 3744 1818
rect 3726 1818 3744 1836
rect 3726 1836 3744 1854
rect 3726 1854 3744 1872
rect 3726 1872 3744 1890
rect 3726 1890 3744 1908
rect 3726 1908 3744 1926
rect 3726 1926 3744 1944
rect 3726 1944 3744 1962
rect 3726 1962 3744 1980
rect 3726 1980 3744 1998
rect 3726 1998 3744 2016
rect 3726 2016 3744 2034
rect 3726 2034 3744 2052
rect 3726 2052 3744 2070
rect 3726 2070 3744 2088
rect 3726 2088 3744 2106
rect 3726 2106 3744 2124
rect 3726 2124 3744 2142
rect 3726 2142 3744 2160
rect 3726 2160 3744 2178
rect 3726 2178 3744 2196
rect 3726 2196 3744 2214
rect 3726 2214 3744 2232
rect 3726 2232 3744 2250
rect 3726 2250 3744 2268
rect 3726 2268 3744 2286
rect 3726 2286 3744 2304
rect 3726 2304 3744 2322
rect 3726 2322 3744 2340
rect 3726 2340 3744 2358
rect 3726 2358 3744 2376
rect 3726 2376 3744 2394
rect 3726 2394 3744 2412
rect 3726 2412 3744 2430
rect 3726 2430 3744 2448
rect 3726 2448 3744 2466
rect 3726 2466 3744 2484
rect 3726 2484 3744 2502
rect 3726 2502 3744 2520
rect 3726 2520 3744 2538
rect 3726 2538 3744 2556
rect 3726 2556 3744 2574
rect 3726 2574 3744 2592
rect 3726 2592 3744 2610
rect 3726 2610 3744 2628
rect 3726 2628 3744 2646
rect 3726 2646 3744 2664
rect 3726 2664 3744 2682
rect 3726 2934 3744 2952
rect 3726 2952 3744 2970
rect 3726 2970 3744 2988
rect 3726 2988 3744 3006
rect 3726 3006 3744 3024
rect 3726 3024 3744 3042
rect 3726 3042 3744 3060
rect 3726 3060 3744 3078
rect 3726 3078 3744 3096
rect 3726 3096 3744 3114
rect 3726 3114 3744 3132
rect 3726 3132 3744 3150
rect 3726 3150 3744 3168
rect 3726 3168 3744 3186
rect 3726 3186 3744 3204
rect 3726 3204 3744 3222
rect 3726 3222 3744 3240
rect 3726 3240 3744 3258
rect 3726 3258 3744 3276
rect 3726 3276 3744 3294
rect 3726 3294 3744 3312
rect 3726 3312 3744 3330
rect 3726 3330 3744 3348
rect 3726 3348 3744 3366
rect 3726 3366 3744 3384
rect 3726 3384 3744 3402
rect 3726 3402 3744 3420
rect 3726 3420 3744 3438
rect 3726 3438 3744 3456
rect 3726 3456 3744 3474
rect 3726 3474 3744 3492
rect 3726 3492 3744 3510
rect 3726 3510 3744 3528
rect 3726 3528 3744 3546
rect 3726 3546 3744 3564
rect 3726 3564 3744 3582
rect 3726 3582 3744 3600
rect 3726 3600 3744 3618
rect 3726 3618 3744 3636
rect 3726 3636 3744 3654
rect 3726 3654 3744 3672
rect 3726 3672 3744 3690
rect 3726 3690 3744 3708
rect 3726 3708 3744 3726
rect 3726 3726 3744 3744
rect 3726 3744 3744 3762
rect 3726 3762 3744 3780
rect 3726 3780 3744 3798
rect 3726 3798 3744 3816
rect 3726 3816 3744 3834
rect 3726 3834 3744 3852
rect 3726 3852 3744 3870
rect 3726 3870 3744 3888
rect 3726 3888 3744 3906
rect 3726 3906 3744 3924
rect 3726 3924 3744 3942
rect 3726 3942 3744 3960
rect 3726 3960 3744 3978
rect 3726 3978 3744 3996
rect 3726 3996 3744 4014
rect 3726 4014 3744 4032
rect 3726 4032 3744 4050
rect 3726 4050 3744 4068
rect 3726 4068 3744 4086
rect 3726 4086 3744 4104
rect 3726 4104 3744 4122
rect 3726 4122 3744 4140
rect 3726 4140 3744 4158
rect 3726 4158 3744 4176
rect 3726 4176 3744 4194
rect 3726 4194 3744 4212
rect 3726 4212 3744 4230
rect 3726 4230 3744 4248
rect 3726 4248 3744 4266
rect 3726 4266 3744 4284
rect 3726 4284 3744 4302
rect 3726 4302 3744 4320
rect 3726 4320 3744 4338
rect 3726 4338 3744 4356
rect 3726 4356 3744 4374
rect 3726 4374 3744 4392
rect 3726 4392 3744 4410
rect 3726 4410 3744 4428
rect 3726 4428 3744 4446
rect 3726 4446 3744 4464
rect 3726 4464 3744 4482
rect 3726 4482 3744 4500
rect 3726 4500 3744 4518
rect 3726 4518 3744 4536
rect 3726 4536 3744 4554
rect 3726 4554 3744 4572
rect 3726 4572 3744 4590
rect 3726 4590 3744 4608
rect 3726 4608 3744 4626
rect 3726 4626 3744 4644
rect 3726 4644 3744 4662
rect 3726 4662 3744 4680
rect 3726 4680 3744 4698
rect 3726 4698 3744 4716
rect 3726 4716 3744 4734
rect 3726 4734 3744 4752
rect 3726 4752 3744 4770
rect 3726 4770 3744 4788
rect 3726 4788 3744 4806
rect 3726 4806 3744 4824
rect 3726 4824 3744 4842
rect 3726 4842 3744 4860
rect 3726 4860 3744 4878
rect 3726 4878 3744 4896
rect 3726 4896 3744 4914
rect 3726 4914 3744 4932
rect 3726 4932 3744 4950
rect 3726 4950 3744 4968
rect 3726 4968 3744 4986
rect 3726 4986 3744 5004
rect 3726 5004 3744 5022
rect 3726 5022 3744 5040
rect 3726 5040 3744 5058
rect 3726 5058 3744 5076
rect 3726 5076 3744 5094
rect 3726 5094 3744 5112
rect 3726 5112 3744 5130
rect 3726 5130 3744 5148
rect 3726 5148 3744 5166
rect 3726 5166 3744 5184
rect 3726 5184 3744 5202
rect 3726 5202 3744 5220
rect 3726 5220 3744 5238
rect 3726 5238 3744 5256
rect 3726 5256 3744 5274
rect 3726 5274 3744 5292
rect 3726 5292 3744 5310
rect 3726 5310 3744 5328
rect 3726 5328 3744 5346
rect 3726 5346 3744 5364
rect 3726 5364 3744 5382
rect 3726 5382 3744 5400
rect 3726 5400 3744 5418
rect 3726 5418 3744 5436
rect 3726 5436 3744 5454
rect 3726 5454 3744 5472
rect 3726 6642 3744 6660
rect 3726 6660 3744 6678
rect 3726 6678 3744 6696
rect 3726 6696 3744 6714
rect 3726 6714 3744 6732
rect 3726 6732 3744 6750
rect 3726 6750 3744 6768
rect 3726 6768 3744 6786
rect 3726 6786 3744 6804
rect 3726 6804 3744 6822
rect 3726 6822 3744 6840
rect 3726 6840 3744 6858
rect 3726 6858 3744 6876
rect 3726 6876 3744 6894
rect 3726 6894 3744 6912
rect 3726 6912 3744 6930
rect 3726 6930 3744 6948
rect 3726 6948 3744 6966
rect 3726 6966 3744 6984
rect 3726 6984 3744 7002
rect 3726 7002 3744 7020
rect 3726 7020 3744 7038
rect 3726 7038 3744 7056
rect 3726 7056 3744 7074
rect 3726 7074 3744 7092
rect 3726 7092 3744 7110
rect 3726 7110 3744 7128
rect 3726 7128 3744 7146
rect 3726 7146 3744 7164
rect 3726 7164 3744 7182
rect 3726 7182 3744 7200
rect 3726 7200 3744 7218
rect 3726 7218 3744 7236
rect 3726 7236 3744 7254
rect 3726 7254 3744 7272
rect 3744 0 3762 18
rect 3744 18 3762 36
rect 3744 36 3762 54
rect 3744 54 3762 72
rect 3744 72 3762 90
rect 3744 90 3762 108
rect 3744 108 3762 126
rect 3744 126 3762 144
rect 3744 144 3762 162
rect 3744 162 3762 180
rect 3744 180 3762 198
rect 3744 198 3762 216
rect 3744 216 3762 234
rect 3744 234 3762 252
rect 3744 252 3762 270
rect 3744 270 3762 288
rect 3744 288 3762 306
rect 3744 306 3762 324
rect 3744 324 3762 342
rect 3744 342 3762 360
rect 3744 360 3762 378
rect 3744 378 3762 396
rect 3744 396 3762 414
rect 3744 414 3762 432
rect 3744 432 3762 450
rect 3744 450 3762 468
rect 3744 468 3762 486
rect 3744 486 3762 504
rect 3744 504 3762 522
rect 3744 522 3762 540
rect 3744 540 3762 558
rect 3744 558 3762 576
rect 3744 576 3762 594
rect 3744 594 3762 612
rect 3744 612 3762 630
rect 3744 864 3762 882
rect 3744 882 3762 900
rect 3744 900 3762 918
rect 3744 918 3762 936
rect 3744 936 3762 954
rect 3744 954 3762 972
rect 3744 972 3762 990
rect 3744 990 3762 1008
rect 3744 1008 3762 1026
rect 3744 1026 3762 1044
rect 3744 1044 3762 1062
rect 3744 1062 3762 1080
rect 3744 1080 3762 1098
rect 3744 1098 3762 1116
rect 3744 1116 3762 1134
rect 3744 1134 3762 1152
rect 3744 1152 3762 1170
rect 3744 1170 3762 1188
rect 3744 1188 3762 1206
rect 3744 1206 3762 1224
rect 3744 1224 3762 1242
rect 3744 1242 3762 1260
rect 3744 1260 3762 1278
rect 3744 1278 3762 1296
rect 3744 1296 3762 1314
rect 3744 1314 3762 1332
rect 3744 1332 3762 1350
rect 3744 1350 3762 1368
rect 3744 1368 3762 1386
rect 3744 1620 3762 1638
rect 3744 1638 3762 1656
rect 3744 1656 3762 1674
rect 3744 1674 3762 1692
rect 3744 1692 3762 1710
rect 3744 1710 3762 1728
rect 3744 1728 3762 1746
rect 3744 1746 3762 1764
rect 3744 1764 3762 1782
rect 3744 1782 3762 1800
rect 3744 1800 3762 1818
rect 3744 1818 3762 1836
rect 3744 1836 3762 1854
rect 3744 1854 3762 1872
rect 3744 1872 3762 1890
rect 3744 1890 3762 1908
rect 3744 1908 3762 1926
rect 3744 1926 3762 1944
rect 3744 1944 3762 1962
rect 3744 1962 3762 1980
rect 3744 1980 3762 1998
rect 3744 1998 3762 2016
rect 3744 2016 3762 2034
rect 3744 2034 3762 2052
rect 3744 2052 3762 2070
rect 3744 2070 3762 2088
rect 3744 2088 3762 2106
rect 3744 2106 3762 2124
rect 3744 2124 3762 2142
rect 3744 2142 3762 2160
rect 3744 2160 3762 2178
rect 3744 2178 3762 2196
rect 3744 2196 3762 2214
rect 3744 2214 3762 2232
rect 3744 2232 3762 2250
rect 3744 2250 3762 2268
rect 3744 2268 3762 2286
rect 3744 2286 3762 2304
rect 3744 2304 3762 2322
rect 3744 2322 3762 2340
rect 3744 2340 3762 2358
rect 3744 2358 3762 2376
rect 3744 2376 3762 2394
rect 3744 2394 3762 2412
rect 3744 2412 3762 2430
rect 3744 2430 3762 2448
rect 3744 2448 3762 2466
rect 3744 2466 3762 2484
rect 3744 2484 3762 2502
rect 3744 2502 3762 2520
rect 3744 2520 3762 2538
rect 3744 2538 3762 2556
rect 3744 2556 3762 2574
rect 3744 2574 3762 2592
rect 3744 2592 3762 2610
rect 3744 2610 3762 2628
rect 3744 2628 3762 2646
rect 3744 2646 3762 2664
rect 3744 2664 3762 2682
rect 3744 2682 3762 2700
rect 3744 2700 3762 2718
rect 3744 2970 3762 2988
rect 3744 2988 3762 3006
rect 3744 3006 3762 3024
rect 3744 3024 3762 3042
rect 3744 3042 3762 3060
rect 3744 3060 3762 3078
rect 3744 3078 3762 3096
rect 3744 3096 3762 3114
rect 3744 3114 3762 3132
rect 3744 3132 3762 3150
rect 3744 3150 3762 3168
rect 3744 3168 3762 3186
rect 3744 3186 3762 3204
rect 3744 3204 3762 3222
rect 3744 3222 3762 3240
rect 3744 3240 3762 3258
rect 3744 3258 3762 3276
rect 3744 3276 3762 3294
rect 3744 3294 3762 3312
rect 3744 3312 3762 3330
rect 3744 3330 3762 3348
rect 3744 3348 3762 3366
rect 3744 3366 3762 3384
rect 3744 3384 3762 3402
rect 3744 3402 3762 3420
rect 3744 3420 3762 3438
rect 3744 3438 3762 3456
rect 3744 3456 3762 3474
rect 3744 3474 3762 3492
rect 3744 3492 3762 3510
rect 3744 3510 3762 3528
rect 3744 3528 3762 3546
rect 3744 3546 3762 3564
rect 3744 3564 3762 3582
rect 3744 3582 3762 3600
rect 3744 3600 3762 3618
rect 3744 3618 3762 3636
rect 3744 3636 3762 3654
rect 3744 3654 3762 3672
rect 3744 3672 3762 3690
rect 3744 3690 3762 3708
rect 3744 3708 3762 3726
rect 3744 3726 3762 3744
rect 3744 3744 3762 3762
rect 3744 3762 3762 3780
rect 3744 3780 3762 3798
rect 3744 3798 3762 3816
rect 3744 3816 3762 3834
rect 3744 3834 3762 3852
rect 3744 3852 3762 3870
rect 3744 3870 3762 3888
rect 3744 3888 3762 3906
rect 3744 3906 3762 3924
rect 3744 3924 3762 3942
rect 3744 3942 3762 3960
rect 3744 3960 3762 3978
rect 3744 3978 3762 3996
rect 3744 3996 3762 4014
rect 3744 4014 3762 4032
rect 3744 4032 3762 4050
rect 3744 4050 3762 4068
rect 3744 4068 3762 4086
rect 3744 4086 3762 4104
rect 3744 4104 3762 4122
rect 3744 4122 3762 4140
rect 3744 4140 3762 4158
rect 3744 4158 3762 4176
rect 3744 4176 3762 4194
rect 3744 4194 3762 4212
rect 3744 4212 3762 4230
rect 3744 4230 3762 4248
rect 3744 4248 3762 4266
rect 3744 4266 3762 4284
rect 3744 4284 3762 4302
rect 3744 4302 3762 4320
rect 3744 4320 3762 4338
rect 3744 4338 3762 4356
rect 3744 4356 3762 4374
rect 3744 4374 3762 4392
rect 3744 4392 3762 4410
rect 3744 4410 3762 4428
rect 3744 4428 3762 4446
rect 3744 4446 3762 4464
rect 3744 4464 3762 4482
rect 3744 4482 3762 4500
rect 3744 4500 3762 4518
rect 3744 4518 3762 4536
rect 3744 4536 3762 4554
rect 3744 4554 3762 4572
rect 3744 4572 3762 4590
rect 3744 4590 3762 4608
rect 3744 4608 3762 4626
rect 3744 4626 3762 4644
rect 3744 4644 3762 4662
rect 3744 4662 3762 4680
rect 3744 4680 3762 4698
rect 3744 4698 3762 4716
rect 3744 4716 3762 4734
rect 3744 4734 3762 4752
rect 3744 4752 3762 4770
rect 3744 4770 3762 4788
rect 3744 4788 3762 4806
rect 3744 4806 3762 4824
rect 3744 4824 3762 4842
rect 3744 4842 3762 4860
rect 3744 4860 3762 4878
rect 3744 4878 3762 4896
rect 3744 4896 3762 4914
rect 3744 4914 3762 4932
rect 3744 4932 3762 4950
rect 3744 4950 3762 4968
rect 3744 4968 3762 4986
rect 3744 4986 3762 5004
rect 3744 5004 3762 5022
rect 3744 5022 3762 5040
rect 3744 5040 3762 5058
rect 3744 5058 3762 5076
rect 3744 5076 3762 5094
rect 3744 5094 3762 5112
rect 3744 5112 3762 5130
rect 3744 5130 3762 5148
rect 3744 5148 3762 5166
rect 3744 5166 3762 5184
rect 3744 5184 3762 5202
rect 3744 5202 3762 5220
rect 3744 5220 3762 5238
rect 3744 5238 3762 5256
rect 3744 5256 3762 5274
rect 3744 5274 3762 5292
rect 3744 5292 3762 5310
rect 3744 5310 3762 5328
rect 3744 5328 3762 5346
rect 3744 5346 3762 5364
rect 3744 5364 3762 5382
rect 3744 5382 3762 5400
rect 3744 5400 3762 5418
rect 3744 5418 3762 5436
rect 3744 5436 3762 5454
rect 3744 5454 3762 5472
rect 3744 5472 3762 5490
rect 3744 5490 3762 5508
rect 3744 6642 3762 6660
rect 3744 6660 3762 6678
rect 3744 6678 3762 6696
rect 3744 6696 3762 6714
rect 3744 6714 3762 6732
rect 3744 6732 3762 6750
rect 3744 6750 3762 6768
rect 3744 6768 3762 6786
rect 3744 6786 3762 6804
rect 3744 6804 3762 6822
rect 3744 6822 3762 6840
rect 3744 6840 3762 6858
rect 3744 6858 3762 6876
rect 3744 6876 3762 6894
rect 3744 6894 3762 6912
rect 3744 6912 3762 6930
rect 3744 6930 3762 6948
rect 3744 6948 3762 6966
rect 3744 6966 3762 6984
rect 3744 6984 3762 7002
rect 3744 7002 3762 7020
rect 3744 7020 3762 7038
rect 3744 7038 3762 7056
rect 3744 7056 3762 7074
rect 3744 7074 3762 7092
rect 3744 7092 3762 7110
rect 3744 7110 3762 7128
rect 3744 7128 3762 7146
rect 3744 7146 3762 7164
rect 3744 7164 3762 7182
rect 3744 7182 3762 7200
rect 3744 7200 3762 7218
rect 3744 7218 3762 7236
rect 3744 7236 3762 7254
rect 3744 7254 3762 7272
rect 3762 0 3780 18
rect 3762 18 3780 36
rect 3762 36 3780 54
rect 3762 54 3780 72
rect 3762 72 3780 90
rect 3762 90 3780 108
rect 3762 108 3780 126
rect 3762 126 3780 144
rect 3762 144 3780 162
rect 3762 162 3780 180
rect 3762 180 3780 198
rect 3762 198 3780 216
rect 3762 216 3780 234
rect 3762 234 3780 252
rect 3762 252 3780 270
rect 3762 270 3780 288
rect 3762 288 3780 306
rect 3762 306 3780 324
rect 3762 324 3780 342
rect 3762 342 3780 360
rect 3762 360 3780 378
rect 3762 378 3780 396
rect 3762 396 3780 414
rect 3762 414 3780 432
rect 3762 432 3780 450
rect 3762 450 3780 468
rect 3762 468 3780 486
rect 3762 486 3780 504
rect 3762 504 3780 522
rect 3762 522 3780 540
rect 3762 540 3780 558
rect 3762 558 3780 576
rect 3762 576 3780 594
rect 3762 594 3780 612
rect 3762 612 3780 630
rect 3762 864 3780 882
rect 3762 882 3780 900
rect 3762 900 3780 918
rect 3762 918 3780 936
rect 3762 936 3780 954
rect 3762 954 3780 972
rect 3762 972 3780 990
rect 3762 990 3780 1008
rect 3762 1008 3780 1026
rect 3762 1026 3780 1044
rect 3762 1044 3780 1062
rect 3762 1062 3780 1080
rect 3762 1080 3780 1098
rect 3762 1098 3780 1116
rect 3762 1116 3780 1134
rect 3762 1134 3780 1152
rect 3762 1152 3780 1170
rect 3762 1170 3780 1188
rect 3762 1188 3780 1206
rect 3762 1206 3780 1224
rect 3762 1224 3780 1242
rect 3762 1242 3780 1260
rect 3762 1260 3780 1278
rect 3762 1278 3780 1296
rect 3762 1296 3780 1314
rect 3762 1314 3780 1332
rect 3762 1332 3780 1350
rect 3762 1350 3780 1368
rect 3762 1368 3780 1386
rect 3762 1386 3780 1404
rect 3762 1638 3780 1656
rect 3762 1656 3780 1674
rect 3762 1674 3780 1692
rect 3762 1692 3780 1710
rect 3762 1710 3780 1728
rect 3762 1728 3780 1746
rect 3762 1746 3780 1764
rect 3762 1764 3780 1782
rect 3762 1782 3780 1800
rect 3762 1800 3780 1818
rect 3762 1818 3780 1836
rect 3762 1836 3780 1854
rect 3762 1854 3780 1872
rect 3762 1872 3780 1890
rect 3762 1890 3780 1908
rect 3762 1908 3780 1926
rect 3762 1926 3780 1944
rect 3762 1944 3780 1962
rect 3762 1962 3780 1980
rect 3762 1980 3780 1998
rect 3762 1998 3780 2016
rect 3762 2016 3780 2034
rect 3762 2034 3780 2052
rect 3762 2052 3780 2070
rect 3762 2070 3780 2088
rect 3762 2088 3780 2106
rect 3762 2106 3780 2124
rect 3762 2124 3780 2142
rect 3762 2142 3780 2160
rect 3762 2160 3780 2178
rect 3762 2178 3780 2196
rect 3762 2196 3780 2214
rect 3762 2214 3780 2232
rect 3762 2232 3780 2250
rect 3762 2250 3780 2268
rect 3762 2268 3780 2286
rect 3762 2286 3780 2304
rect 3762 2304 3780 2322
rect 3762 2322 3780 2340
rect 3762 2340 3780 2358
rect 3762 2358 3780 2376
rect 3762 2376 3780 2394
rect 3762 2394 3780 2412
rect 3762 2412 3780 2430
rect 3762 2430 3780 2448
rect 3762 2448 3780 2466
rect 3762 2466 3780 2484
rect 3762 2484 3780 2502
rect 3762 2502 3780 2520
rect 3762 2520 3780 2538
rect 3762 2538 3780 2556
rect 3762 2556 3780 2574
rect 3762 2574 3780 2592
rect 3762 2592 3780 2610
rect 3762 2610 3780 2628
rect 3762 2628 3780 2646
rect 3762 2646 3780 2664
rect 3762 2664 3780 2682
rect 3762 2682 3780 2700
rect 3762 2700 3780 2718
rect 3762 2718 3780 2736
rect 3762 2988 3780 3006
rect 3762 3006 3780 3024
rect 3762 3024 3780 3042
rect 3762 3042 3780 3060
rect 3762 3060 3780 3078
rect 3762 3078 3780 3096
rect 3762 3096 3780 3114
rect 3762 3114 3780 3132
rect 3762 3132 3780 3150
rect 3762 3150 3780 3168
rect 3762 3168 3780 3186
rect 3762 3186 3780 3204
rect 3762 3204 3780 3222
rect 3762 3222 3780 3240
rect 3762 3240 3780 3258
rect 3762 3258 3780 3276
rect 3762 3276 3780 3294
rect 3762 3294 3780 3312
rect 3762 3312 3780 3330
rect 3762 3330 3780 3348
rect 3762 3348 3780 3366
rect 3762 3366 3780 3384
rect 3762 3384 3780 3402
rect 3762 3402 3780 3420
rect 3762 3420 3780 3438
rect 3762 3438 3780 3456
rect 3762 3456 3780 3474
rect 3762 3474 3780 3492
rect 3762 3492 3780 3510
rect 3762 3510 3780 3528
rect 3762 3528 3780 3546
rect 3762 3546 3780 3564
rect 3762 3564 3780 3582
rect 3762 3582 3780 3600
rect 3762 3600 3780 3618
rect 3762 3618 3780 3636
rect 3762 3636 3780 3654
rect 3762 3654 3780 3672
rect 3762 3672 3780 3690
rect 3762 3690 3780 3708
rect 3762 3708 3780 3726
rect 3762 3726 3780 3744
rect 3762 3744 3780 3762
rect 3762 3762 3780 3780
rect 3762 3780 3780 3798
rect 3762 3798 3780 3816
rect 3762 3816 3780 3834
rect 3762 3834 3780 3852
rect 3762 3852 3780 3870
rect 3762 3870 3780 3888
rect 3762 3888 3780 3906
rect 3762 3906 3780 3924
rect 3762 3924 3780 3942
rect 3762 3942 3780 3960
rect 3762 3960 3780 3978
rect 3762 3978 3780 3996
rect 3762 3996 3780 4014
rect 3762 4014 3780 4032
rect 3762 4032 3780 4050
rect 3762 4050 3780 4068
rect 3762 4068 3780 4086
rect 3762 4086 3780 4104
rect 3762 4104 3780 4122
rect 3762 4122 3780 4140
rect 3762 4140 3780 4158
rect 3762 4158 3780 4176
rect 3762 4176 3780 4194
rect 3762 4194 3780 4212
rect 3762 4212 3780 4230
rect 3762 4230 3780 4248
rect 3762 4248 3780 4266
rect 3762 4266 3780 4284
rect 3762 4284 3780 4302
rect 3762 4302 3780 4320
rect 3762 4320 3780 4338
rect 3762 4338 3780 4356
rect 3762 4356 3780 4374
rect 3762 4374 3780 4392
rect 3762 4392 3780 4410
rect 3762 4410 3780 4428
rect 3762 4428 3780 4446
rect 3762 4446 3780 4464
rect 3762 4464 3780 4482
rect 3762 4482 3780 4500
rect 3762 4500 3780 4518
rect 3762 4518 3780 4536
rect 3762 4536 3780 4554
rect 3762 4554 3780 4572
rect 3762 4572 3780 4590
rect 3762 4590 3780 4608
rect 3762 4608 3780 4626
rect 3762 4626 3780 4644
rect 3762 4644 3780 4662
rect 3762 4662 3780 4680
rect 3762 4680 3780 4698
rect 3762 4698 3780 4716
rect 3762 4716 3780 4734
rect 3762 4734 3780 4752
rect 3762 4752 3780 4770
rect 3762 4770 3780 4788
rect 3762 4788 3780 4806
rect 3762 4806 3780 4824
rect 3762 4824 3780 4842
rect 3762 4842 3780 4860
rect 3762 4860 3780 4878
rect 3762 4878 3780 4896
rect 3762 4896 3780 4914
rect 3762 4914 3780 4932
rect 3762 4932 3780 4950
rect 3762 4950 3780 4968
rect 3762 4968 3780 4986
rect 3762 4986 3780 5004
rect 3762 5004 3780 5022
rect 3762 5022 3780 5040
rect 3762 5040 3780 5058
rect 3762 5058 3780 5076
rect 3762 5076 3780 5094
rect 3762 5094 3780 5112
rect 3762 5112 3780 5130
rect 3762 5130 3780 5148
rect 3762 5148 3780 5166
rect 3762 5166 3780 5184
rect 3762 5184 3780 5202
rect 3762 5202 3780 5220
rect 3762 5220 3780 5238
rect 3762 5238 3780 5256
rect 3762 5256 3780 5274
rect 3762 5274 3780 5292
rect 3762 5292 3780 5310
rect 3762 5310 3780 5328
rect 3762 5328 3780 5346
rect 3762 5346 3780 5364
rect 3762 5364 3780 5382
rect 3762 5382 3780 5400
rect 3762 5400 3780 5418
rect 3762 5418 3780 5436
rect 3762 5436 3780 5454
rect 3762 5454 3780 5472
rect 3762 5472 3780 5490
rect 3762 5490 3780 5508
rect 3762 5508 3780 5526
rect 3762 5526 3780 5544
rect 3762 6642 3780 6660
rect 3762 6660 3780 6678
rect 3762 6678 3780 6696
rect 3762 6696 3780 6714
rect 3762 6714 3780 6732
rect 3762 6732 3780 6750
rect 3762 6750 3780 6768
rect 3762 6768 3780 6786
rect 3762 6786 3780 6804
rect 3762 6804 3780 6822
rect 3762 6822 3780 6840
rect 3762 6840 3780 6858
rect 3762 6858 3780 6876
rect 3762 6876 3780 6894
rect 3762 6894 3780 6912
rect 3762 6912 3780 6930
rect 3762 6930 3780 6948
rect 3762 6948 3780 6966
rect 3762 6966 3780 6984
rect 3762 6984 3780 7002
rect 3762 7002 3780 7020
rect 3762 7020 3780 7038
rect 3762 7038 3780 7056
rect 3762 7056 3780 7074
rect 3762 7074 3780 7092
rect 3762 7092 3780 7110
rect 3762 7110 3780 7128
rect 3762 7128 3780 7146
rect 3762 7146 3780 7164
rect 3762 7164 3780 7182
rect 3762 7182 3780 7200
rect 3762 7200 3780 7218
rect 3762 7218 3780 7236
rect 3762 7236 3780 7254
rect 3762 7254 3780 7272
rect 3780 0 3798 18
rect 3780 18 3798 36
rect 3780 36 3798 54
rect 3780 54 3798 72
rect 3780 72 3798 90
rect 3780 90 3798 108
rect 3780 108 3798 126
rect 3780 126 3798 144
rect 3780 144 3798 162
rect 3780 162 3798 180
rect 3780 180 3798 198
rect 3780 198 3798 216
rect 3780 216 3798 234
rect 3780 234 3798 252
rect 3780 252 3798 270
rect 3780 270 3798 288
rect 3780 288 3798 306
rect 3780 306 3798 324
rect 3780 324 3798 342
rect 3780 342 3798 360
rect 3780 360 3798 378
rect 3780 378 3798 396
rect 3780 396 3798 414
rect 3780 414 3798 432
rect 3780 432 3798 450
rect 3780 450 3798 468
rect 3780 468 3798 486
rect 3780 486 3798 504
rect 3780 504 3798 522
rect 3780 522 3798 540
rect 3780 540 3798 558
rect 3780 558 3798 576
rect 3780 576 3798 594
rect 3780 594 3798 612
rect 3780 612 3798 630
rect 3780 864 3798 882
rect 3780 882 3798 900
rect 3780 900 3798 918
rect 3780 918 3798 936
rect 3780 936 3798 954
rect 3780 954 3798 972
rect 3780 972 3798 990
rect 3780 990 3798 1008
rect 3780 1008 3798 1026
rect 3780 1026 3798 1044
rect 3780 1044 3798 1062
rect 3780 1062 3798 1080
rect 3780 1080 3798 1098
rect 3780 1098 3798 1116
rect 3780 1116 3798 1134
rect 3780 1134 3798 1152
rect 3780 1152 3798 1170
rect 3780 1170 3798 1188
rect 3780 1188 3798 1206
rect 3780 1206 3798 1224
rect 3780 1224 3798 1242
rect 3780 1242 3798 1260
rect 3780 1260 3798 1278
rect 3780 1278 3798 1296
rect 3780 1296 3798 1314
rect 3780 1314 3798 1332
rect 3780 1332 3798 1350
rect 3780 1350 3798 1368
rect 3780 1368 3798 1386
rect 3780 1386 3798 1404
rect 3780 1404 3798 1422
rect 3780 1638 3798 1656
rect 3780 1656 3798 1674
rect 3780 1674 3798 1692
rect 3780 1692 3798 1710
rect 3780 1710 3798 1728
rect 3780 1728 3798 1746
rect 3780 1746 3798 1764
rect 3780 1764 3798 1782
rect 3780 1782 3798 1800
rect 3780 1800 3798 1818
rect 3780 1818 3798 1836
rect 3780 1836 3798 1854
rect 3780 1854 3798 1872
rect 3780 1872 3798 1890
rect 3780 1890 3798 1908
rect 3780 1908 3798 1926
rect 3780 1926 3798 1944
rect 3780 1944 3798 1962
rect 3780 1962 3798 1980
rect 3780 1980 3798 1998
rect 3780 1998 3798 2016
rect 3780 2016 3798 2034
rect 3780 2034 3798 2052
rect 3780 2052 3798 2070
rect 3780 2070 3798 2088
rect 3780 2088 3798 2106
rect 3780 2106 3798 2124
rect 3780 2124 3798 2142
rect 3780 2142 3798 2160
rect 3780 2160 3798 2178
rect 3780 2178 3798 2196
rect 3780 2196 3798 2214
rect 3780 2214 3798 2232
rect 3780 2232 3798 2250
rect 3780 2250 3798 2268
rect 3780 2268 3798 2286
rect 3780 2286 3798 2304
rect 3780 2304 3798 2322
rect 3780 2322 3798 2340
rect 3780 2340 3798 2358
rect 3780 2358 3798 2376
rect 3780 2376 3798 2394
rect 3780 2394 3798 2412
rect 3780 2412 3798 2430
rect 3780 2430 3798 2448
rect 3780 2448 3798 2466
rect 3780 2466 3798 2484
rect 3780 2484 3798 2502
rect 3780 2502 3798 2520
rect 3780 2520 3798 2538
rect 3780 2538 3798 2556
rect 3780 2556 3798 2574
rect 3780 2574 3798 2592
rect 3780 2592 3798 2610
rect 3780 2610 3798 2628
rect 3780 2628 3798 2646
rect 3780 2646 3798 2664
rect 3780 2664 3798 2682
rect 3780 2682 3798 2700
rect 3780 2700 3798 2718
rect 3780 2718 3798 2736
rect 3780 2736 3798 2754
rect 3780 2754 3798 2772
rect 3780 3024 3798 3042
rect 3780 3042 3798 3060
rect 3780 3060 3798 3078
rect 3780 3078 3798 3096
rect 3780 3096 3798 3114
rect 3780 3114 3798 3132
rect 3780 3132 3798 3150
rect 3780 3150 3798 3168
rect 3780 3168 3798 3186
rect 3780 3186 3798 3204
rect 3780 3204 3798 3222
rect 3780 3222 3798 3240
rect 3780 3240 3798 3258
rect 3780 3258 3798 3276
rect 3780 3276 3798 3294
rect 3780 3294 3798 3312
rect 3780 3312 3798 3330
rect 3780 3330 3798 3348
rect 3780 3348 3798 3366
rect 3780 3366 3798 3384
rect 3780 3384 3798 3402
rect 3780 3402 3798 3420
rect 3780 3420 3798 3438
rect 3780 3438 3798 3456
rect 3780 3456 3798 3474
rect 3780 3474 3798 3492
rect 3780 3492 3798 3510
rect 3780 3510 3798 3528
rect 3780 3528 3798 3546
rect 3780 3546 3798 3564
rect 3780 3564 3798 3582
rect 3780 3582 3798 3600
rect 3780 3600 3798 3618
rect 3780 3618 3798 3636
rect 3780 3636 3798 3654
rect 3780 3654 3798 3672
rect 3780 3672 3798 3690
rect 3780 3690 3798 3708
rect 3780 3708 3798 3726
rect 3780 3726 3798 3744
rect 3780 3744 3798 3762
rect 3780 3762 3798 3780
rect 3780 3780 3798 3798
rect 3780 3798 3798 3816
rect 3780 3816 3798 3834
rect 3780 3834 3798 3852
rect 3780 3852 3798 3870
rect 3780 3870 3798 3888
rect 3780 3888 3798 3906
rect 3780 3906 3798 3924
rect 3780 3924 3798 3942
rect 3780 3942 3798 3960
rect 3780 3960 3798 3978
rect 3780 3978 3798 3996
rect 3780 3996 3798 4014
rect 3780 4014 3798 4032
rect 3780 4032 3798 4050
rect 3780 4050 3798 4068
rect 3780 4068 3798 4086
rect 3780 4086 3798 4104
rect 3780 4104 3798 4122
rect 3780 4122 3798 4140
rect 3780 4140 3798 4158
rect 3780 4158 3798 4176
rect 3780 4176 3798 4194
rect 3780 4194 3798 4212
rect 3780 4212 3798 4230
rect 3780 4230 3798 4248
rect 3780 4248 3798 4266
rect 3780 4266 3798 4284
rect 3780 4284 3798 4302
rect 3780 4302 3798 4320
rect 3780 4320 3798 4338
rect 3780 4338 3798 4356
rect 3780 4356 3798 4374
rect 3780 4374 3798 4392
rect 3780 4392 3798 4410
rect 3780 4410 3798 4428
rect 3780 4428 3798 4446
rect 3780 4446 3798 4464
rect 3780 4464 3798 4482
rect 3780 4482 3798 4500
rect 3780 4500 3798 4518
rect 3780 4518 3798 4536
rect 3780 4536 3798 4554
rect 3780 4554 3798 4572
rect 3780 4572 3798 4590
rect 3780 4590 3798 4608
rect 3780 4608 3798 4626
rect 3780 4626 3798 4644
rect 3780 4644 3798 4662
rect 3780 4662 3798 4680
rect 3780 4680 3798 4698
rect 3780 4698 3798 4716
rect 3780 4716 3798 4734
rect 3780 4734 3798 4752
rect 3780 4752 3798 4770
rect 3780 4770 3798 4788
rect 3780 4788 3798 4806
rect 3780 4806 3798 4824
rect 3780 4824 3798 4842
rect 3780 4842 3798 4860
rect 3780 4860 3798 4878
rect 3780 4878 3798 4896
rect 3780 4896 3798 4914
rect 3780 4914 3798 4932
rect 3780 4932 3798 4950
rect 3780 4950 3798 4968
rect 3780 4968 3798 4986
rect 3780 4986 3798 5004
rect 3780 5004 3798 5022
rect 3780 5022 3798 5040
rect 3780 5040 3798 5058
rect 3780 5058 3798 5076
rect 3780 5076 3798 5094
rect 3780 5094 3798 5112
rect 3780 5112 3798 5130
rect 3780 5130 3798 5148
rect 3780 5148 3798 5166
rect 3780 5166 3798 5184
rect 3780 5184 3798 5202
rect 3780 5202 3798 5220
rect 3780 5220 3798 5238
rect 3780 5238 3798 5256
rect 3780 5256 3798 5274
rect 3780 5274 3798 5292
rect 3780 5292 3798 5310
rect 3780 5310 3798 5328
rect 3780 5328 3798 5346
rect 3780 5346 3798 5364
rect 3780 5364 3798 5382
rect 3780 5382 3798 5400
rect 3780 5400 3798 5418
rect 3780 5418 3798 5436
rect 3780 5436 3798 5454
rect 3780 5454 3798 5472
rect 3780 5472 3798 5490
rect 3780 5490 3798 5508
rect 3780 5508 3798 5526
rect 3780 5526 3798 5544
rect 3780 5544 3798 5562
rect 3780 5562 3798 5580
rect 3780 5580 3798 5598
rect 3780 6642 3798 6660
rect 3780 6660 3798 6678
rect 3780 6678 3798 6696
rect 3780 6696 3798 6714
rect 3780 6714 3798 6732
rect 3780 6732 3798 6750
rect 3780 6750 3798 6768
rect 3780 6768 3798 6786
rect 3780 6786 3798 6804
rect 3780 6804 3798 6822
rect 3780 6822 3798 6840
rect 3780 6840 3798 6858
rect 3780 6858 3798 6876
rect 3780 6876 3798 6894
rect 3780 6894 3798 6912
rect 3780 6912 3798 6930
rect 3780 6930 3798 6948
rect 3780 6948 3798 6966
rect 3780 6966 3798 6984
rect 3780 6984 3798 7002
rect 3780 7002 3798 7020
rect 3780 7020 3798 7038
rect 3780 7038 3798 7056
rect 3780 7056 3798 7074
rect 3780 7074 3798 7092
rect 3780 7092 3798 7110
rect 3780 7110 3798 7128
rect 3780 7128 3798 7146
rect 3780 7146 3798 7164
rect 3780 7164 3798 7182
rect 3780 7182 3798 7200
rect 3780 7200 3798 7218
rect 3780 7218 3798 7236
rect 3780 7236 3798 7254
rect 3780 7254 3798 7272
rect 3798 0 3816 18
rect 3798 18 3816 36
rect 3798 36 3816 54
rect 3798 54 3816 72
rect 3798 72 3816 90
rect 3798 90 3816 108
rect 3798 108 3816 126
rect 3798 126 3816 144
rect 3798 144 3816 162
rect 3798 162 3816 180
rect 3798 180 3816 198
rect 3798 198 3816 216
rect 3798 216 3816 234
rect 3798 234 3816 252
rect 3798 252 3816 270
rect 3798 270 3816 288
rect 3798 288 3816 306
rect 3798 306 3816 324
rect 3798 324 3816 342
rect 3798 342 3816 360
rect 3798 360 3816 378
rect 3798 378 3816 396
rect 3798 396 3816 414
rect 3798 414 3816 432
rect 3798 432 3816 450
rect 3798 450 3816 468
rect 3798 468 3816 486
rect 3798 486 3816 504
rect 3798 504 3816 522
rect 3798 522 3816 540
rect 3798 540 3816 558
rect 3798 558 3816 576
rect 3798 576 3816 594
rect 3798 594 3816 612
rect 3798 612 3816 630
rect 3798 864 3816 882
rect 3798 882 3816 900
rect 3798 900 3816 918
rect 3798 918 3816 936
rect 3798 936 3816 954
rect 3798 954 3816 972
rect 3798 972 3816 990
rect 3798 990 3816 1008
rect 3798 1008 3816 1026
rect 3798 1026 3816 1044
rect 3798 1044 3816 1062
rect 3798 1062 3816 1080
rect 3798 1080 3816 1098
rect 3798 1098 3816 1116
rect 3798 1116 3816 1134
rect 3798 1134 3816 1152
rect 3798 1152 3816 1170
rect 3798 1170 3816 1188
rect 3798 1188 3816 1206
rect 3798 1206 3816 1224
rect 3798 1224 3816 1242
rect 3798 1242 3816 1260
rect 3798 1260 3816 1278
rect 3798 1278 3816 1296
rect 3798 1296 3816 1314
rect 3798 1314 3816 1332
rect 3798 1332 3816 1350
rect 3798 1350 3816 1368
rect 3798 1368 3816 1386
rect 3798 1386 3816 1404
rect 3798 1404 3816 1422
rect 3798 1422 3816 1440
rect 3798 1656 3816 1674
rect 3798 1674 3816 1692
rect 3798 1692 3816 1710
rect 3798 1710 3816 1728
rect 3798 1728 3816 1746
rect 3798 1746 3816 1764
rect 3798 1764 3816 1782
rect 3798 1782 3816 1800
rect 3798 1800 3816 1818
rect 3798 1818 3816 1836
rect 3798 1836 3816 1854
rect 3798 1854 3816 1872
rect 3798 1872 3816 1890
rect 3798 1890 3816 1908
rect 3798 1908 3816 1926
rect 3798 1926 3816 1944
rect 3798 1944 3816 1962
rect 3798 1962 3816 1980
rect 3798 1980 3816 1998
rect 3798 1998 3816 2016
rect 3798 2016 3816 2034
rect 3798 2034 3816 2052
rect 3798 2052 3816 2070
rect 3798 2070 3816 2088
rect 3798 2088 3816 2106
rect 3798 2106 3816 2124
rect 3798 2124 3816 2142
rect 3798 2142 3816 2160
rect 3798 2160 3816 2178
rect 3798 2178 3816 2196
rect 3798 2196 3816 2214
rect 3798 2214 3816 2232
rect 3798 2232 3816 2250
rect 3798 2250 3816 2268
rect 3798 2268 3816 2286
rect 3798 2286 3816 2304
rect 3798 2304 3816 2322
rect 3798 2322 3816 2340
rect 3798 2340 3816 2358
rect 3798 2358 3816 2376
rect 3798 2376 3816 2394
rect 3798 2394 3816 2412
rect 3798 2412 3816 2430
rect 3798 2430 3816 2448
rect 3798 2448 3816 2466
rect 3798 2466 3816 2484
rect 3798 2484 3816 2502
rect 3798 2502 3816 2520
rect 3798 2520 3816 2538
rect 3798 2538 3816 2556
rect 3798 2556 3816 2574
rect 3798 2574 3816 2592
rect 3798 2592 3816 2610
rect 3798 2610 3816 2628
rect 3798 2628 3816 2646
rect 3798 2646 3816 2664
rect 3798 2664 3816 2682
rect 3798 2682 3816 2700
rect 3798 2700 3816 2718
rect 3798 2718 3816 2736
rect 3798 2736 3816 2754
rect 3798 2754 3816 2772
rect 3798 2772 3816 2790
rect 3798 3042 3816 3060
rect 3798 3060 3816 3078
rect 3798 3078 3816 3096
rect 3798 3096 3816 3114
rect 3798 3114 3816 3132
rect 3798 3132 3816 3150
rect 3798 3150 3816 3168
rect 3798 3168 3816 3186
rect 3798 3186 3816 3204
rect 3798 3204 3816 3222
rect 3798 3222 3816 3240
rect 3798 3240 3816 3258
rect 3798 3258 3816 3276
rect 3798 3276 3816 3294
rect 3798 3294 3816 3312
rect 3798 3312 3816 3330
rect 3798 3330 3816 3348
rect 3798 3348 3816 3366
rect 3798 3366 3816 3384
rect 3798 3384 3816 3402
rect 3798 3402 3816 3420
rect 3798 3420 3816 3438
rect 3798 3438 3816 3456
rect 3798 3456 3816 3474
rect 3798 3474 3816 3492
rect 3798 3492 3816 3510
rect 3798 3510 3816 3528
rect 3798 3528 3816 3546
rect 3798 3546 3816 3564
rect 3798 3564 3816 3582
rect 3798 3582 3816 3600
rect 3798 3600 3816 3618
rect 3798 3618 3816 3636
rect 3798 3636 3816 3654
rect 3798 3654 3816 3672
rect 3798 3672 3816 3690
rect 3798 3690 3816 3708
rect 3798 3708 3816 3726
rect 3798 3726 3816 3744
rect 3798 3744 3816 3762
rect 3798 3762 3816 3780
rect 3798 3780 3816 3798
rect 3798 3798 3816 3816
rect 3798 3816 3816 3834
rect 3798 3834 3816 3852
rect 3798 3852 3816 3870
rect 3798 3870 3816 3888
rect 3798 3888 3816 3906
rect 3798 3906 3816 3924
rect 3798 3924 3816 3942
rect 3798 3942 3816 3960
rect 3798 3960 3816 3978
rect 3798 3978 3816 3996
rect 3798 3996 3816 4014
rect 3798 4014 3816 4032
rect 3798 4032 3816 4050
rect 3798 4050 3816 4068
rect 3798 4068 3816 4086
rect 3798 4086 3816 4104
rect 3798 4104 3816 4122
rect 3798 4122 3816 4140
rect 3798 4140 3816 4158
rect 3798 4158 3816 4176
rect 3798 4176 3816 4194
rect 3798 4194 3816 4212
rect 3798 4212 3816 4230
rect 3798 4230 3816 4248
rect 3798 4248 3816 4266
rect 3798 4266 3816 4284
rect 3798 4284 3816 4302
rect 3798 4302 3816 4320
rect 3798 4320 3816 4338
rect 3798 4338 3816 4356
rect 3798 4356 3816 4374
rect 3798 4374 3816 4392
rect 3798 4392 3816 4410
rect 3798 4410 3816 4428
rect 3798 4428 3816 4446
rect 3798 4446 3816 4464
rect 3798 4464 3816 4482
rect 3798 4482 3816 4500
rect 3798 4500 3816 4518
rect 3798 4518 3816 4536
rect 3798 4536 3816 4554
rect 3798 4554 3816 4572
rect 3798 4572 3816 4590
rect 3798 4590 3816 4608
rect 3798 4608 3816 4626
rect 3798 4626 3816 4644
rect 3798 4644 3816 4662
rect 3798 4662 3816 4680
rect 3798 4680 3816 4698
rect 3798 4698 3816 4716
rect 3798 4716 3816 4734
rect 3798 4734 3816 4752
rect 3798 4752 3816 4770
rect 3798 4770 3816 4788
rect 3798 4788 3816 4806
rect 3798 4806 3816 4824
rect 3798 4824 3816 4842
rect 3798 4842 3816 4860
rect 3798 4860 3816 4878
rect 3798 4878 3816 4896
rect 3798 4896 3816 4914
rect 3798 4914 3816 4932
rect 3798 4932 3816 4950
rect 3798 4950 3816 4968
rect 3798 4968 3816 4986
rect 3798 4986 3816 5004
rect 3798 5004 3816 5022
rect 3798 5022 3816 5040
rect 3798 5040 3816 5058
rect 3798 5058 3816 5076
rect 3798 5076 3816 5094
rect 3798 5094 3816 5112
rect 3798 5112 3816 5130
rect 3798 5130 3816 5148
rect 3798 5148 3816 5166
rect 3798 5166 3816 5184
rect 3798 5184 3816 5202
rect 3798 5202 3816 5220
rect 3798 5220 3816 5238
rect 3798 5238 3816 5256
rect 3798 5256 3816 5274
rect 3798 5274 3816 5292
rect 3798 5292 3816 5310
rect 3798 5310 3816 5328
rect 3798 5328 3816 5346
rect 3798 5346 3816 5364
rect 3798 5364 3816 5382
rect 3798 5382 3816 5400
rect 3798 5400 3816 5418
rect 3798 5418 3816 5436
rect 3798 5436 3816 5454
rect 3798 5454 3816 5472
rect 3798 5472 3816 5490
rect 3798 5490 3816 5508
rect 3798 5508 3816 5526
rect 3798 5526 3816 5544
rect 3798 5544 3816 5562
rect 3798 5562 3816 5580
rect 3798 5580 3816 5598
rect 3798 5598 3816 5616
rect 3798 5616 3816 5634
rect 3798 6642 3816 6660
rect 3798 6660 3816 6678
rect 3798 6678 3816 6696
rect 3798 6696 3816 6714
rect 3798 6714 3816 6732
rect 3798 6732 3816 6750
rect 3798 6750 3816 6768
rect 3798 6768 3816 6786
rect 3798 6786 3816 6804
rect 3798 6804 3816 6822
rect 3798 6822 3816 6840
rect 3798 6840 3816 6858
rect 3798 6858 3816 6876
rect 3798 6876 3816 6894
rect 3798 6894 3816 6912
rect 3798 6912 3816 6930
rect 3798 6930 3816 6948
rect 3798 6948 3816 6966
rect 3798 6966 3816 6984
rect 3798 6984 3816 7002
rect 3798 7002 3816 7020
rect 3798 7020 3816 7038
rect 3798 7038 3816 7056
rect 3798 7056 3816 7074
rect 3798 7074 3816 7092
rect 3798 7092 3816 7110
rect 3798 7110 3816 7128
rect 3798 7128 3816 7146
rect 3798 7146 3816 7164
rect 3798 7164 3816 7182
rect 3798 7182 3816 7200
rect 3798 7200 3816 7218
rect 3798 7218 3816 7236
rect 3798 7236 3816 7254
rect 3798 7254 3816 7272
rect 3816 0 3834 18
rect 3816 18 3834 36
rect 3816 36 3834 54
rect 3816 54 3834 72
rect 3816 72 3834 90
rect 3816 90 3834 108
rect 3816 108 3834 126
rect 3816 126 3834 144
rect 3816 144 3834 162
rect 3816 162 3834 180
rect 3816 180 3834 198
rect 3816 198 3834 216
rect 3816 216 3834 234
rect 3816 234 3834 252
rect 3816 252 3834 270
rect 3816 270 3834 288
rect 3816 288 3834 306
rect 3816 306 3834 324
rect 3816 324 3834 342
rect 3816 342 3834 360
rect 3816 360 3834 378
rect 3816 378 3834 396
rect 3816 396 3834 414
rect 3816 414 3834 432
rect 3816 432 3834 450
rect 3816 450 3834 468
rect 3816 468 3834 486
rect 3816 486 3834 504
rect 3816 504 3834 522
rect 3816 522 3834 540
rect 3816 540 3834 558
rect 3816 558 3834 576
rect 3816 576 3834 594
rect 3816 594 3834 612
rect 3816 612 3834 630
rect 3816 864 3834 882
rect 3816 882 3834 900
rect 3816 900 3834 918
rect 3816 918 3834 936
rect 3816 936 3834 954
rect 3816 954 3834 972
rect 3816 972 3834 990
rect 3816 990 3834 1008
rect 3816 1008 3834 1026
rect 3816 1026 3834 1044
rect 3816 1044 3834 1062
rect 3816 1062 3834 1080
rect 3816 1080 3834 1098
rect 3816 1098 3834 1116
rect 3816 1116 3834 1134
rect 3816 1134 3834 1152
rect 3816 1152 3834 1170
rect 3816 1170 3834 1188
rect 3816 1188 3834 1206
rect 3816 1206 3834 1224
rect 3816 1224 3834 1242
rect 3816 1242 3834 1260
rect 3816 1260 3834 1278
rect 3816 1278 3834 1296
rect 3816 1296 3834 1314
rect 3816 1314 3834 1332
rect 3816 1332 3834 1350
rect 3816 1350 3834 1368
rect 3816 1368 3834 1386
rect 3816 1386 3834 1404
rect 3816 1404 3834 1422
rect 3816 1422 3834 1440
rect 3816 1674 3834 1692
rect 3816 1692 3834 1710
rect 3816 1710 3834 1728
rect 3816 1728 3834 1746
rect 3816 1746 3834 1764
rect 3816 1764 3834 1782
rect 3816 1782 3834 1800
rect 3816 1800 3834 1818
rect 3816 1818 3834 1836
rect 3816 1836 3834 1854
rect 3816 1854 3834 1872
rect 3816 1872 3834 1890
rect 3816 1890 3834 1908
rect 3816 1908 3834 1926
rect 3816 1926 3834 1944
rect 3816 1944 3834 1962
rect 3816 1962 3834 1980
rect 3816 1980 3834 1998
rect 3816 1998 3834 2016
rect 3816 2016 3834 2034
rect 3816 2034 3834 2052
rect 3816 2052 3834 2070
rect 3816 2070 3834 2088
rect 3816 2088 3834 2106
rect 3816 2106 3834 2124
rect 3816 2124 3834 2142
rect 3816 2142 3834 2160
rect 3816 2160 3834 2178
rect 3816 2178 3834 2196
rect 3816 2196 3834 2214
rect 3816 2214 3834 2232
rect 3816 2232 3834 2250
rect 3816 2250 3834 2268
rect 3816 2268 3834 2286
rect 3816 2286 3834 2304
rect 3816 2304 3834 2322
rect 3816 2322 3834 2340
rect 3816 2340 3834 2358
rect 3816 2358 3834 2376
rect 3816 2376 3834 2394
rect 3816 2394 3834 2412
rect 3816 2412 3834 2430
rect 3816 2430 3834 2448
rect 3816 2448 3834 2466
rect 3816 2466 3834 2484
rect 3816 2484 3834 2502
rect 3816 2502 3834 2520
rect 3816 2520 3834 2538
rect 3816 2538 3834 2556
rect 3816 2556 3834 2574
rect 3816 2574 3834 2592
rect 3816 2592 3834 2610
rect 3816 2610 3834 2628
rect 3816 2628 3834 2646
rect 3816 2646 3834 2664
rect 3816 2664 3834 2682
rect 3816 2682 3834 2700
rect 3816 2700 3834 2718
rect 3816 2718 3834 2736
rect 3816 2736 3834 2754
rect 3816 2754 3834 2772
rect 3816 2772 3834 2790
rect 3816 2790 3834 2808
rect 3816 2808 3834 2826
rect 3816 3060 3834 3078
rect 3816 3078 3834 3096
rect 3816 3096 3834 3114
rect 3816 3114 3834 3132
rect 3816 3132 3834 3150
rect 3816 3150 3834 3168
rect 3816 3168 3834 3186
rect 3816 3186 3834 3204
rect 3816 3204 3834 3222
rect 3816 3222 3834 3240
rect 3816 3240 3834 3258
rect 3816 3258 3834 3276
rect 3816 3276 3834 3294
rect 3816 3294 3834 3312
rect 3816 3312 3834 3330
rect 3816 3330 3834 3348
rect 3816 3348 3834 3366
rect 3816 3366 3834 3384
rect 3816 3384 3834 3402
rect 3816 3402 3834 3420
rect 3816 3420 3834 3438
rect 3816 3438 3834 3456
rect 3816 3456 3834 3474
rect 3816 3474 3834 3492
rect 3816 3492 3834 3510
rect 3816 3510 3834 3528
rect 3816 3528 3834 3546
rect 3816 3546 3834 3564
rect 3816 3564 3834 3582
rect 3816 3582 3834 3600
rect 3816 3600 3834 3618
rect 3816 3618 3834 3636
rect 3816 3636 3834 3654
rect 3816 3654 3834 3672
rect 3816 3672 3834 3690
rect 3816 3690 3834 3708
rect 3816 3708 3834 3726
rect 3816 3726 3834 3744
rect 3816 3744 3834 3762
rect 3816 3762 3834 3780
rect 3816 3780 3834 3798
rect 3816 3798 3834 3816
rect 3816 3816 3834 3834
rect 3816 3834 3834 3852
rect 3816 3852 3834 3870
rect 3816 3870 3834 3888
rect 3816 3888 3834 3906
rect 3816 3906 3834 3924
rect 3816 3924 3834 3942
rect 3816 3942 3834 3960
rect 3816 3960 3834 3978
rect 3816 3978 3834 3996
rect 3816 3996 3834 4014
rect 3816 4014 3834 4032
rect 3816 4032 3834 4050
rect 3816 4050 3834 4068
rect 3816 4068 3834 4086
rect 3816 4086 3834 4104
rect 3816 4104 3834 4122
rect 3816 4122 3834 4140
rect 3816 4140 3834 4158
rect 3816 4158 3834 4176
rect 3816 4176 3834 4194
rect 3816 4194 3834 4212
rect 3816 4212 3834 4230
rect 3816 4230 3834 4248
rect 3816 4248 3834 4266
rect 3816 4266 3834 4284
rect 3816 4284 3834 4302
rect 3816 4302 3834 4320
rect 3816 4320 3834 4338
rect 3816 4338 3834 4356
rect 3816 4356 3834 4374
rect 3816 4374 3834 4392
rect 3816 4392 3834 4410
rect 3816 4410 3834 4428
rect 3816 4428 3834 4446
rect 3816 4446 3834 4464
rect 3816 4464 3834 4482
rect 3816 4482 3834 4500
rect 3816 4500 3834 4518
rect 3816 4518 3834 4536
rect 3816 4536 3834 4554
rect 3816 4554 3834 4572
rect 3816 4572 3834 4590
rect 3816 4590 3834 4608
rect 3816 4608 3834 4626
rect 3816 4626 3834 4644
rect 3816 4644 3834 4662
rect 3816 4662 3834 4680
rect 3816 4680 3834 4698
rect 3816 4698 3834 4716
rect 3816 4716 3834 4734
rect 3816 4734 3834 4752
rect 3816 4752 3834 4770
rect 3816 4770 3834 4788
rect 3816 4788 3834 4806
rect 3816 4806 3834 4824
rect 3816 4824 3834 4842
rect 3816 4842 3834 4860
rect 3816 4860 3834 4878
rect 3816 4878 3834 4896
rect 3816 4896 3834 4914
rect 3816 4914 3834 4932
rect 3816 4932 3834 4950
rect 3816 4950 3834 4968
rect 3816 4968 3834 4986
rect 3816 4986 3834 5004
rect 3816 5004 3834 5022
rect 3816 5022 3834 5040
rect 3816 5040 3834 5058
rect 3816 5058 3834 5076
rect 3816 5076 3834 5094
rect 3816 5094 3834 5112
rect 3816 5112 3834 5130
rect 3816 5130 3834 5148
rect 3816 5148 3834 5166
rect 3816 5166 3834 5184
rect 3816 5184 3834 5202
rect 3816 5202 3834 5220
rect 3816 5220 3834 5238
rect 3816 5238 3834 5256
rect 3816 5256 3834 5274
rect 3816 5274 3834 5292
rect 3816 5292 3834 5310
rect 3816 5310 3834 5328
rect 3816 5328 3834 5346
rect 3816 5346 3834 5364
rect 3816 5364 3834 5382
rect 3816 5382 3834 5400
rect 3816 5400 3834 5418
rect 3816 5418 3834 5436
rect 3816 5436 3834 5454
rect 3816 5454 3834 5472
rect 3816 5472 3834 5490
rect 3816 5490 3834 5508
rect 3816 5508 3834 5526
rect 3816 5526 3834 5544
rect 3816 5544 3834 5562
rect 3816 5562 3834 5580
rect 3816 5580 3834 5598
rect 3816 5598 3834 5616
rect 3816 5616 3834 5634
rect 3816 5634 3834 5652
rect 3816 5652 3834 5670
rect 3816 5670 3834 5688
rect 3816 6642 3834 6660
rect 3816 6660 3834 6678
rect 3816 6678 3834 6696
rect 3816 6696 3834 6714
rect 3816 6714 3834 6732
rect 3816 6732 3834 6750
rect 3816 6750 3834 6768
rect 3816 6768 3834 6786
rect 3816 6786 3834 6804
rect 3816 6804 3834 6822
rect 3816 6822 3834 6840
rect 3816 6840 3834 6858
rect 3816 6858 3834 6876
rect 3816 6876 3834 6894
rect 3816 6894 3834 6912
rect 3816 6912 3834 6930
rect 3816 6930 3834 6948
rect 3816 6948 3834 6966
rect 3816 6966 3834 6984
rect 3816 6984 3834 7002
rect 3816 7002 3834 7020
rect 3816 7020 3834 7038
rect 3816 7038 3834 7056
rect 3816 7056 3834 7074
rect 3816 7074 3834 7092
rect 3816 7092 3834 7110
rect 3816 7110 3834 7128
rect 3816 7128 3834 7146
rect 3816 7146 3834 7164
rect 3816 7164 3834 7182
rect 3816 7182 3834 7200
rect 3816 7200 3834 7218
rect 3816 7218 3834 7236
rect 3816 7236 3834 7254
rect 3816 7254 3834 7272
rect 3834 0 3852 18
rect 3834 18 3852 36
rect 3834 36 3852 54
rect 3834 54 3852 72
rect 3834 72 3852 90
rect 3834 90 3852 108
rect 3834 108 3852 126
rect 3834 126 3852 144
rect 3834 144 3852 162
rect 3834 162 3852 180
rect 3834 180 3852 198
rect 3834 198 3852 216
rect 3834 216 3852 234
rect 3834 234 3852 252
rect 3834 252 3852 270
rect 3834 270 3852 288
rect 3834 288 3852 306
rect 3834 306 3852 324
rect 3834 324 3852 342
rect 3834 342 3852 360
rect 3834 360 3852 378
rect 3834 378 3852 396
rect 3834 396 3852 414
rect 3834 414 3852 432
rect 3834 432 3852 450
rect 3834 450 3852 468
rect 3834 468 3852 486
rect 3834 486 3852 504
rect 3834 504 3852 522
rect 3834 522 3852 540
rect 3834 540 3852 558
rect 3834 558 3852 576
rect 3834 576 3852 594
rect 3834 594 3852 612
rect 3834 612 3852 630
rect 3834 864 3852 882
rect 3834 882 3852 900
rect 3834 900 3852 918
rect 3834 918 3852 936
rect 3834 936 3852 954
rect 3834 954 3852 972
rect 3834 972 3852 990
rect 3834 990 3852 1008
rect 3834 1008 3852 1026
rect 3834 1026 3852 1044
rect 3834 1044 3852 1062
rect 3834 1062 3852 1080
rect 3834 1080 3852 1098
rect 3834 1098 3852 1116
rect 3834 1116 3852 1134
rect 3834 1134 3852 1152
rect 3834 1152 3852 1170
rect 3834 1170 3852 1188
rect 3834 1188 3852 1206
rect 3834 1206 3852 1224
rect 3834 1224 3852 1242
rect 3834 1242 3852 1260
rect 3834 1260 3852 1278
rect 3834 1278 3852 1296
rect 3834 1296 3852 1314
rect 3834 1314 3852 1332
rect 3834 1332 3852 1350
rect 3834 1350 3852 1368
rect 3834 1368 3852 1386
rect 3834 1386 3852 1404
rect 3834 1404 3852 1422
rect 3834 1422 3852 1440
rect 3834 1440 3852 1458
rect 3834 1692 3852 1710
rect 3834 1710 3852 1728
rect 3834 1728 3852 1746
rect 3834 1746 3852 1764
rect 3834 1764 3852 1782
rect 3834 1782 3852 1800
rect 3834 1800 3852 1818
rect 3834 1818 3852 1836
rect 3834 1836 3852 1854
rect 3834 1854 3852 1872
rect 3834 1872 3852 1890
rect 3834 1890 3852 1908
rect 3834 1908 3852 1926
rect 3834 1926 3852 1944
rect 3834 1944 3852 1962
rect 3834 1962 3852 1980
rect 3834 1980 3852 1998
rect 3834 1998 3852 2016
rect 3834 2016 3852 2034
rect 3834 2034 3852 2052
rect 3834 2052 3852 2070
rect 3834 2070 3852 2088
rect 3834 2088 3852 2106
rect 3834 2106 3852 2124
rect 3834 2124 3852 2142
rect 3834 2142 3852 2160
rect 3834 2160 3852 2178
rect 3834 2178 3852 2196
rect 3834 2196 3852 2214
rect 3834 2214 3852 2232
rect 3834 2232 3852 2250
rect 3834 2250 3852 2268
rect 3834 2268 3852 2286
rect 3834 2286 3852 2304
rect 3834 2304 3852 2322
rect 3834 2322 3852 2340
rect 3834 2340 3852 2358
rect 3834 2358 3852 2376
rect 3834 2376 3852 2394
rect 3834 2394 3852 2412
rect 3834 2412 3852 2430
rect 3834 2430 3852 2448
rect 3834 2448 3852 2466
rect 3834 2466 3852 2484
rect 3834 2484 3852 2502
rect 3834 2502 3852 2520
rect 3834 2520 3852 2538
rect 3834 2538 3852 2556
rect 3834 2556 3852 2574
rect 3834 2574 3852 2592
rect 3834 2592 3852 2610
rect 3834 2610 3852 2628
rect 3834 2628 3852 2646
rect 3834 2646 3852 2664
rect 3834 2664 3852 2682
rect 3834 2682 3852 2700
rect 3834 2700 3852 2718
rect 3834 2718 3852 2736
rect 3834 2736 3852 2754
rect 3834 2754 3852 2772
rect 3834 2772 3852 2790
rect 3834 2790 3852 2808
rect 3834 2808 3852 2826
rect 3834 2826 3852 2844
rect 3834 3096 3852 3114
rect 3834 3114 3852 3132
rect 3834 3132 3852 3150
rect 3834 3150 3852 3168
rect 3834 3168 3852 3186
rect 3834 3186 3852 3204
rect 3834 3204 3852 3222
rect 3834 3222 3852 3240
rect 3834 3240 3852 3258
rect 3834 3258 3852 3276
rect 3834 3276 3852 3294
rect 3834 3294 3852 3312
rect 3834 3312 3852 3330
rect 3834 3330 3852 3348
rect 3834 3348 3852 3366
rect 3834 3366 3852 3384
rect 3834 3384 3852 3402
rect 3834 3402 3852 3420
rect 3834 3420 3852 3438
rect 3834 3438 3852 3456
rect 3834 3456 3852 3474
rect 3834 3474 3852 3492
rect 3834 3492 3852 3510
rect 3834 3510 3852 3528
rect 3834 3528 3852 3546
rect 3834 3546 3852 3564
rect 3834 3564 3852 3582
rect 3834 3582 3852 3600
rect 3834 3600 3852 3618
rect 3834 3618 3852 3636
rect 3834 3636 3852 3654
rect 3834 3654 3852 3672
rect 3834 3672 3852 3690
rect 3834 3690 3852 3708
rect 3834 3708 3852 3726
rect 3834 3726 3852 3744
rect 3834 3744 3852 3762
rect 3834 3762 3852 3780
rect 3834 3780 3852 3798
rect 3834 3798 3852 3816
rect 3834 3816 3852 3834
rect 3834 3834 3852 3852
rect 3834 3852 3852 3870
rect 3834 3870 3852 3888
rect 3834 3888 3852 3906
rect 3834 3906 3852 3924
rect 3834 3924 3852 3942
rect 3834 3942 3852 3960
rect 3834 3960 3852 3978
rect 3834 3978 3852 3996
rect 3834 3996 3852 4014
rect 3834 4014 3852 4032
rect 3834 4032 3852 4050
rect 3834 4050 3852 4068
rect 3834 4068 3852 4086
rect 3834 4086 3852 4104
rect 3834 4104 3852 4122
rect 3834 4122 3852 4140
rect 3834 4140 3852 4158
rect 3834 4158 3852 4176
rect 3834 4176 3852 4194
rect 3834 4194 3852 4212
rect 3834 4212 3852 4230
rect 3834 4230 3852 4248
rect 3834 4248 3852 4266
rect 3834 4266 3852 4284
rect 3834 4284 3852 4302
rect 3834 4302 3852 4320
rect 3834 4320 3852 4338
rect 3834 4338 3852 4356
rect 3834 4356 3852 4374
rect 3834 4374 3852 4392
rect 3834 4392 3852 4410
rect 3834 4410 3852 4428
rect 3834 4428 3852 4446
rect 3834 4446 3852 4464
rect 3834 4464 3852 4482
rect 3834 4482 3852 4500
rect 3834 4500 3852 4518
rect 3834 4518 3852 4536
rect 3834 4536 3852 4554
rect 3834 4554 3852 4572
rect 3834 4572 3852 4590
rect 3834 4590 3852 4608
rect 3834 4608 3852 4626
rect 3834 4626 3852 4644
rect 3834 4644 3852 4662
rect 3834 4662 3852 4680
rect 3834 4680 3852 4698
rect 3834 4698 3852 4716
rect 3834 4716 3852 4734
rect 3834 4734 3852 4752
rect 3834 4752 3852 4770
rect 3834 4770 3852 4788
rect 3834 4788 3852 4806
rect 3834 4806 3852 4824
rect 3834 4824 3852 4842
rect 3834 4842 3852 4860
rect 3834 4860 3852 4878
rect 3834 4878 3852 4896
rect 3834 4896 3852 4914
rect 3834 4914 3852 4932
rect 3834 4932 3852 4950
rect 3834 4950 3852 4968
rect 3834 4968 3852 4986
rect 3834 4986 3852 5004
rect 3834 5004 3852 5022
rect 3834 5022 3852 5040
rect 3834 5040 3852 5058
rect 3834 5058 3852 5076
rect 3834 5076 3852 5094
rect 3834 5094 3852 5112
rect 3834 5112 3852 5130
rect 3834 5130 3852 5148
rect 3834 5148 3852 5166
rect 3834 5166 3852 5184
rect 3834 5184 3852 5202
rect 3834 5202 3852 5220
rect 3834 5220 3852 5238
rect 3834 5238 3852 5256
rect 3834 5256 3852 5274
rect 3834 5274 3852 5292
rect 3834 5292 3852 5310
rect 3834 5310 3852 5328
rect 3834 5328 3852 5346
rect 3834 5346 3852 5364
rect 3834 5364 3852 5382
rect 3834 5382 3852 5400
rect 3834 5400 3852 5418
rect 3834 5418 3852 5436
rect 3834 5436 3852 5454
rect 3834 5454 3852 5472
rect 3834 5472 3852 5490
rect 3834 5490 3852 5508
rect 3834 5508 3852 5526
rect 3834 5526 3852 5544
rect 3834 5544 3852 5562
rect 3834 5562 3852 5580
rect 3834 5580 3852 5598
rect 3834 5598 3852 5616
rect 3834 5616 3852 5634
rect 3834 5634 3852 5652
rect 3834 5652 3852 5670
rect 3834 5670 3852 5688
rect 3834 5688 3852 5706
rect 3834 5706 3852 5724
rect 3834 6642 3852 6660
rect 3834 6660 3852 6678
rect 3834 6678 3852 6696
rect 3834 6696 3852 6714
rect 3834 6714 3852 6732
rect 3834 6732 3852 6750
rect 3834 6750 3852 6768
rect 3834 6768 3852 6786
rect 3834 6786 3852 6804
rect 3834 6804 3852 6822
rect 3834 6822 3852 6840
rect 3834 6840 3852 6858
rect 3834 6858 3852 6876
rect 3834 6876 3852 6894
rect 3834 6894 3852 6912
rect 3834 6912 3852 6930
rect 3834 6930 3852 6948
rect 3834 6948 3852 6966
rect 3834 6966 3852 6984
rect 3834 6984 3852 7002
rect 3834 7002 3852 7020
rect 3834 7020 3852 7038
rect 3834 7038 3852 7056
rect 3834 7056 3852 7074
rect 3834 7074 3852 7092
rect 3834 7092 3852 7110
rect 3834 7110 3852 7128
rect 3834 7128 3852 7146
rect 3834 7146 3852 7164
rect 3834 7164 3852 7182
rect 3834 7182 3852 7200
rect 3834 7200 3852 7218
rect 3834 7218 3852 7236
rect 3834 7236 3852 7254
rect 3834 7254 3852 7272
rect 3852 18 3870 36
rect 3852 36 3870 54
rect 3852 54 3870 72
rect 3852 72 3870 90
rect 3852 90 3870 108
rect 3852 108 3870 126
rect 3852 126 3870 144
rect 3852 144 3870 162
rect 3852 162 3870 180
rect 3852 180 3870 198
rect 3852 198 3870 216
rect 3852 216 3870 234
rect 3852 234 3870 252
rect 3852 252 3870 270
rect 3852 270 3870 288
rect 3852 288 3870 306
rect 3852 306 3870 324
rect 3852 324 3870 342
rect 3852 342 3870 360
rect 3852 360 3870 378
rect 3852 378 3870 396
rect 3852 396 3870 414
rect 3852 414 3870 432
rect 3852 432 3870 450
rect 3852 450 3870 468
rect 3852 468 3870 486
rect 3852 486 3870 504
rect 3852 504 3870 522
rect 3852 522 3870 540
rect 3852 540 3870 558
rect 3852 558 3870 576
rect 3852 576 3870 594
rect 3852 594 3870 612
rect 3852 612 3870 630
rect 3852 864 3870 882
rect 3852 882 3870 900
rect 3852 900 3870 918
rect 3852 918 3870 936
rect 3852 936 3870 954
rect 3852 954 3870 972
rect 3852 972 3870 990
rect 3852 990 3870 1008
rect 3852 1008 3870 1026
rect 3852 1026 3870 1044
rect 3852 1044 3870 1062
rect 3852 1062 3870 1080
rect 3852 1080 3870 1098
rect 3852 1098 3870 1116
rect 3852 1116 3870 1134
rect 3852 1134 3870 1152
rect 3852 1152 3870 1170
rect 3852 1170 3870 1188
rect 3852 1188 3870 1206
rect 3852 1206 3870 1224
rect 3852 1224 3870 1242
rect 3852 1242 3870 1260
rect 3852 1260 3870 1278
rect 3852 1278 3870 1296
rect 3852 1296 3870 1314
rect 3852 1314 3870 1332
rect 3852 1332 3870 1350
rect 3852 1350 3870 1368
rect 3852 1368 3870 1386
rect 3852 1386 3870 1404
rect 3852 1404 3870 1422
rect 3852 1422 3870 1440
rect 3852 1440 3870 1458
rect 3852 1458 3870 1476
rect 3852 1692 3870 1710
rect 3852 1710 3870 1728
rect 3852 1728 3870 1746
rect 3852 1746 3870 1764
rect 3852 1764 3870 1782
rect 3852 1782 3870 1800
rect 3852 1800 3870 1818
rect 3852 1818 3870 1836
rect 3852 1836 3870 1854
rect 3852 1854 3870 1872
rect 3852 1872 3870 1890
rect 3852 1890 3870 1908
rect 3852 1908 3870 1926
rect 3852 1926 3870 1944
rect 3852 1944 3870 1962
rect 3852 1962 3870 1980
rect 3852 1980 3870 1998
rect 3852 1998 3870 2016
rect 3852 2016 3870 2034
rect 3852 2034 3870 2052
rect 3852 2052 3870 2070
rect 3852 2070 3870 2088
rect 3852 2088 3870 2106
rect 3852 2106 3870 2124
rect 3852 2124 3870 2142
rect 3852 2142 3870 2160
rect 3852 2160 3870 2178
rect 3852 2178 3870 2196
rect 3852 2196 3870 2214
rect 3852 2214 3870 2232
rect 3852 2232 3870 2250
rect 3852 2250 3870 2268
rect 3852 2268 3870 2286
rect 3852 2286 3870 2304
rect 3852 2304 3870 2322
rect 3852 2322 3870 2340
rect 3852 2340 3870 2358
rect 3852 2358 3870 2376
rect 3852 2376 3870 2394
rect 3852 2394 3870 2412
rect 3852 2412 3870 2430
rect 3852 2430 3870 2448
rect 3852 2448 3870 2466
rect 3852 2466 3870 2484
rect 3852 2484 3870 2502
rect 3852 2502 3870 2520
rect 3852 2520 3870 2538
rect 3852 2538 3870 2556
rect 3852 2556 3870 2574
rect 3852 2574 3870 2592
rect 3852 2592 3870 2610
rect 3852 2610 3870 2628
rect 3852 2628 3870 2646
rect 3852 2646 3870 2664
rect 3852 2664 3870 2682
rect 3852 2682 3870 2700
rect 3852 2700 3870 2718
rect 3852 2718 3870 2736
rect 3852 2736 3870 2754
rect 3852 2754 3870 2772
rect 3852 2772 3870 2790
rect 3852 2790 3870 2808
rect 3852 2808 3870 2826
rect 3852 2826 3870 2844
rect 3852 2844 3870 2862
rect 3852 2862 3870 2880
rect 3852 3114 3870 3132
rect 3852 3132 3870 3150
rect 3852 3150 3870 3168
rect 3852 3168 3870 3186
rect 3852 3186 3870 3204
rect 3852 3204 3870 3222
rect 3852 3222 3870 3240
rect 3852 3240 3870 3258
rect 3852 3258 3870 3276
rect 3852 3276 3870 3294
rect 3852 3294 3870 3312
rect 3852 3312 3870 3330
rect 3852 3330 3870 3348
rect 3852 3348 3870 3366
rect 3852 3366 3870 3384
rect 3852 3384 3870 3402
rect 3852 3402 3870 3420
rect 3852 3420 3870 3438
rect 3852 3438 3870 3456
rect 3852 3456 3870 3474
rect 3852 3474 3870 3492
rect 3852 3492 3870 3510
rect 3852 3510 3870 3528
rect 3852 3528 3870 3546
rect 3852 3546 3870 3564
rect 3852 3564 3870 3582
rect 3852 3582 3870 3600
rect 3852 3600 3870 3618
rect 3852 3618 3870 3636
rect 3852 3636 3870 3654
rect 3852 3654 3870 3672
rect 3852 3672 3870 3690
rect 3852 3690 3870 3708
rect 3852 3708 3870 3726
rect 3852 3726 3870 3744
rect 3852 3744 3870 3762
rect 3852 3762 3870 3780
rect 3852 3780 3870 3798
rect 3852 3798 3870 3816
rect 3852 3816 3870 3834
rect 3852 3834 3870 3852
rect 3852 3852 3870 3870
rect 3852 3870 3870 3888
rect 3852 3888 3870 3906
rect 3852 3906 3870 3924
rect 3852 3924 3870 3942
rect 3852 3942 3870 3960
rect 3852 3960 3870 3978
rect 3852 3978 3870 3996
rect 3852 3996 3870 4014
rect 3852 4014 3870 4032
rect 3852 4032 3870 4050
rect 3852 4050 3870 4068
rect 3852 4068 3870 4086
rect 3852 4086 3870 4104
rect 3852 4104 3870 4122
rect 3852 4122 3870 4140
rect 3852 4140 3870 4158
rect 3852 4158 3870 4176
rect 3852 4176 3870 4194
rect 3852 4194 3870 4212
rect 3852 4212 3870 4230
rect 3852 4230 3870 4248
rect 3852 4248 3870 4266
rect 3852 4266 3870 4284
rect 3852 4284 3870 4302
rect 3852 4302 3870 4320
rect 3852 4320 3870 4338
rect 3852 4338 3870 4356
rect 3852 4356 3870 4374
rect 3852 4374 3870 4392
rect 3852 4392 3870 4410
rect 3852 4410 3870 4428
rect 3852 4428 3870 4446
rect 3852 4446 3870 4464
rect 3852 4464 3870 4482
rect 3852 4482 3870 4500
rect 3852 4500 3870 4518
rect 3852 4518 3870 4536
rect 3852 4536 3870 4554
rect 3852 4554 3870 4572
rect 3852 4572 3870 4590
rect 3852 4590 3870 4608
rect 3852 4608 3870 4626
rect 3852 4626 3870 4644
rect 3852 4644 3870 4662
rect 3852 4662 3870 4680
rect 3852 4680 3870 4698
rect 3852 4698 3870 4716
rect 3852 4716 3870 4734
rect 3852 4734 3870 4752
rect 3852 4752 3870 4770
rect 3852 4770 3870 4788
rect 3852 4788 3870 4806
rect 3852 4806 3870 4824
rect 3852 4824 3870 4842
rect 3852 4842 3870 4860
rect 3852 4860 3870 4878
rect 3852 4878 3870 4896
rect 3852 4896 3870 4914
rect 3852 4914 3870 4932
rect 3852 4932 3870 4950
rect 3852 4950 3870 4968
rect 3852 4968 3870 4986
rect 3852 4986 3870 5004
rect 3852 5004 3870 5022
rect 3852 5022 3870 5040
rect 3852 5040 3870 5058
rect 3852 5058 3870 5076
rect 3852 5076 3870 5094
rect 3852 5094 3870 5112
rect 3852 5112 3870 5130
rect 3852 5130 3870 5148
rect 3852 5148 3870 5166
rect 3852 5166 3870 5184
rect 3852 5184 3870 5202
rect 3852 5202 3870 5220
rect 3852 5220 3870 5238
rect 3852 5238 3870 5256
rect 3852 5256 3870 5274
rect 3852 5274 3870 5292
rect 3852 5292 3870 5310
rect 3852 5310 3870 5328
rect 3852 5328 3870 5346
rect 3852 5346 3870 5364
rect 3852 5364 3870 5382
rect 3852 5382 3870 5400
rect 3852 5400 3870 5418
rect 3852 5418 3870 5436
rect 3852 5436 3870 5454
rect 3852 5454 3870 5472
rect 3852 5472 3870 5490
rect 3852 5490 3870 5508
rect 3852 5508 3870 5526
rect 3852 5526 3870 5544
rect 3852 5544 3870 5562
rect 3852 5562 3870 5580
rect 3852 5580 3870 5598
rect 3852 5598 3870 5616
rect 3852 5616 3870 5634
rect 3852 5634 3870 5652
rect 3852 5652 3870 5670
rect 3852 5670 3870 5688
rect 3852 5688 3870 5706
rect 3852 5706 3870 5724
rect 3852 5724 3870 5742
rect 3852 5742 3870 5760
rect 3852 6642 3870 6660
rect 3852 6660 3870 6678
rect 3852 6678 3870 6696
rect 3852 6696 3870 6714
rect 3852 6714 3870 6732
rect 3852 6732 3870 6750
rect 3852 6750 3870 6768
rect 3852 6768 3870 6786
rect 3852 6786 3870 6804
rect 3852 6804 3870 6822
rect 3852 6822 3870 6840
rect 3852 6840 3870 6858
rect 3852 6858 3870 6876
rect 3852 6876 3870 6894
rect 3852 6894 3870 6912
rect 3852 6912 3870 6930
rect 3852 6930 3870 6948
rect 3852 6948 3870 6966
rect 3852 6966 3870 6984
rect 3852 6984 3870 7002
rect 3852 7002 3870 7020
rect 3852 7020 3870 7038
rect 3852 7038 3870 7056
rect 3852 7056 3870 7074
rect 3852 7074 3870 7092
rect 3852 7092 3870 7110
rect 3852 7110 3870 7128
rect 3852 7128 3870 7146
rect 3852 7146 3870 7164
rect 3852 7164 3870 7182
rect 3852 7182 3870 7200
rect 3852 7200 3870 7218
rect 3852 7218 3870 7236
rect 3852 7236 3870 7254
rect 3852 7254 3870 7272
rect 3870 18 3888 36
rect 3870 36 3888 54
rect 3870 54 3888 72
rect 3870 72 3888 90
rect 3870 90 3888 108
rect 3870 108 3888 126
rect 3870 126 3888 144
rect 3870 144 3888 162
rect 3870 162 3888 180
rect 3870 180 3888 198
rect 3870 198 3888 216
rect 3870 216 3888 234
rect 3870 234 3888 252
rect 3870 252 3888 270
rect 3870 270 3888 288
rect 3870 288 3888 306
rect 3870 306 3888 324
rect 3870 324 3888 342
rect 3870 342 3888 360
rect 3870 360 3888 378
rect 3870 378 3888 396
rect 3870 396 3888 414
rect 3870 414 3888 432
rect 3870 432 3888 450
rect 3870 450 3888 468
rect 3870 468 3888 486
rect 3870 486 3888 504
rect 3870 504 3888 522
rect 3870 522 3888 540
rect 3870 540 3888 558
rect 3870 558 3888 576
rect 3870 576 3888 594
rect 3870 594 3888 612
rect 3870 612 3888 630
rect 3870 864 3888 882
rect 3870 882 3888 900
rect 3870 900 3888 918
rect 3870 918 3888 936
rect 3870 936 3888 954
rect 3870 954 3888 972
rect 3870 972 3888 990
rect 3870 990 3888 1008
rect 3870 1008 3888 1026
rect 3870 1026 3888 1044
rect 3870 1044 3888 1062
rect 3870 1062 3888 1080
rect 3870 1080 3888 1098
rect 3870 1098 3888 1116
rect 3870 1116 3888 1134
rect 3870 1134 3888 1152
rect 3870 1152 3888 1170
rect 3870 1170 3888 1188
rect 3870 1188 3888 1206
rect 3870 1206 3888 1224
rect 3870 1224 3888 1242
rect 3870 1242 3888 1260
rect 3870 1260 3888 1278
rect 3870 1278 3888 1296
rect 3870 1296 3888 1314
rect 3870 1314 3888 1332
rect 3870 1332 3888 1350
rect 3870 1350 3888 1368
rect 3870 1368 3888 1386
rect 3870 1386 3888 1404
rect 3870 1404 3888 1422
rect 3870 1422 3888 1440
rect 3870 1440 3888 1458
rect 3870 1458 3888 1476
rect 3870 1710 3888 1728
rect 3870 1728 3888 1746
rect 3870 1746 3888 1764
rect 3870 1764 3888 1782
rect 3870 1782 3888 1800
rect 3870 1800 3888 1818
rect 3870 1818 3888 1836
rect 3870 1836 3888 1854
rect 3870 1854 3888 1872
rect 3870 1872 3888 1890
rect 3870 1890 3888 1908
rect 3870 1908 3888 1926
rect 3870 1926 3888 1944
rect 3870 1944 3888 1962
rect 3870 1962 3888 1980
rect 3870 1980 3888 1998
rect 3870 1998 3888 2016
rect 3870 2016 3888 2034
rect 3870 2034 3888 2052
rect 3870 2052 3888 2070
rect 3870 2070 3888 2088
rect 3870 2088 3888 2106
rect 3870 2106 3888 2124
rect 3870 2124 3888 2142
rect 3870 2142 3888 2160
rect 3870 2160 3888 2178
rect 3870 2178 3888 2196
rect 3870 2196 3888 2214
rect 3870 2214 3888 2232
rect 3870 2232 3888 2250
rect 3870 2250 3888 2268
rect 3870 2268 3888 2286
rect 3870 2286 3888 2304
rect 3870 2304 3888 2322
rect 3870 2322 3888 2340
rect 3870 2340 3888 2358
rect 3870 2358 3888 2376
rect 3870 2376 3888 2394
rect 3870 2394 3888 2412
rect 3870 2412 3888 2430
rect 3870 2430 3888 2448
rect 3870 2448 3888 2466
rect 3870 2466 3888 2484
rect 3870 2484 3888 2502
rect 3870 2502 3888 2520
rect 3870 2520 3888 2538
rect 3870 2538 3888 2556
rect 3870 2556 3888 2574
rect 3870 2574 3888 2592
rect 3870 2592 3888 2610
rect 3870 2610 3888 2628
rect 3870 2628 3888 2646
rect 3870 2646 3888 2664
rect 3870 2664 3888 2682
rect 3870 2682 3888 2700
rect 3870 2700 3888 2718
rect 3870 2718 3888 2736
rect 3870 2736 3888 2754
rect 3870 2754 3888 2772
rect 3870 2772 3888 2790
rect 3870 2790 3888 2808
rect 3870 2808 3888 2826
rect 3870 2826 3888 2844
rect 3870 2844 3888 2862
rect 3870 2862 3888 2880
rect 3870 2880 3888 2898
rect 3870 3150 3888 3168
rect 3870 3168 3888 3186
rect 3870 3186 3888 3204
rect 3870 3204 3888 3222
rect 3870 3222 3888 3240
rect 3870 3240 3888 3258
rect 3870 3258 3888 3276
rect 3870 3276 3888 3294
rect 3870 3294 3888 3312
rect 3870 3312 3888 3330
rect 3870 3330 3888 3348
rect 3870 3348 3888 3366
rect 3870 3366 3888 3384
rect 3870 3384 3888 3402
rect 3870 3402 3888 3420
rect 3870 3420 3888 3438
rect 3870 3438 3888 3456
rect 3870 3456 3888 3474
rect 3870 3474 3888 3492
rect 3870 3492 3888 3510
rect 3870 3510 3888 3528
rect 3870 3528 3888 3546
rect 3870 3546 3888 3564
rect 3870 3564 3888 3582
rect 3870 3582 3888 3600
rect 3870 3600 3888 3618
rect 3870 3618 3888 3636
rect 3870 3636 3888 3654
rect 3870 3654 3888 3672
rect 3870 3672 3888 3690
rect 3870 3690 3888 3708
rect 3870 3708 3888 3726
rect 3870 3726 3888 3744
rect 3870 3744 3888 3762
rect 3870 3762 3888 3780
rect 3870 3780 3888 3798
rect 3870 3798 3888 3816
rect 3870 3816 3888 3834
rect 3870 3834 3888 3852
rect 3870 3852 3888 3870
rect 3870 3870 3888 3888
rect 3870 3888 3888 3906
rect 3870 3906 3888 3924
rect 3870 3924 3888 3942
rect 3870 3942 3888 3960
rect 3870 3960 3888 3978
rect 3870 3978 3888 3996
rect 3870 3996 3888 4014
rect 3870 4014 3888 4032
rect 3870 4032 3888 4050
rect 3870 4050 3888 4068
rect 3870 4068 3888 4086
rect 3870 4086 3888 4104
rect 3870 4104 3888 4122
rect 3870 4122 3888 4140
rect 3870 4140 3888 4158
rect 3870 4158 3888 4176
rect 3870 4176 3888 4194
rect 3870 4194 3888 4212
rect 3870 4212 3888 4230
rect 3870 4230 3888 4248
rect 3870 4248 3888 4266
rect 3870 4266 3888 4284
rect 3870 4284 3888 4302
rect 3870 4302 3888 4320
rect 3870 4320 3888 4338
rect 3870 4338 3888 4356
rect 3870 4356 3888 4374
rect 3870 4374 3888 4392
rect 3870 4392 3888 4410
rect 3870 4410 3888 4428
rect 3870 4428 3888 4446
rect 3870 4446 3888 4464
rect 3870 4464 3888 4482
rect 3870 4482 3888 4500
rect 3870 4500 3888 4518
rect 3870 4518 3888 4536
rect 3870 4536 3888 4554
rect 3870 4554 3888 4572
rect 3870 4572 3888 4590
rect 3870 4590 3888 4608
rect 3870 4608 3888 4626
rect 3870 4626 3888 4644
rect 3870 4644 3888 4662
rect 3870 4662 3888 4680
rect 3870 4680 3888 4698
rect 3870 4698 3888 4716
rect 3870 4716 3888 4734
rect 3870 4734 3888 4752
rect 3870 4752 3888 4770
rect 3870 4770 3888 4788
rect 3870 4788 3888 4806
rect 3870 4806 3888 4824
rect 3870 4824 3888 4842
rect 3870 4842 3888 4860
rect 3870 4860 3888 4878
rect 3870 4878 3888 4896
rect 3870 4896 3888 4914
rect 3870 4914 3888 4932
rect 3870 4932 3888 4950
rect 3870 4950 3888 4968
rect 3870 4968 3888 4986
rect 3870 4986 3888 5004
rect 3870 5004 3888 5022
rect 3870 5022 3888 5040
rect 3870 5040 3888 5058
rect 3870 5058 3888 5076
rect 3870 5076 3888 5094
rect 3870 5094 3888 5112
rect 3870 5112 3888 5130
rect 3870 5130 3888 5148
rect 3870 5148 3888 5166
rect 3870 5166 3888 5184
rect 3870 5184 3888 5202
rect 3870 5202 3888 5220
rect 3870 5220 3888 5238
rect 3870 5238 3888 5256
rect 3870 5256 3888 5274
rect 3870 5274 3888 5292
rect 3870 5292 3888 5310
rect 3870 5310 3888 5328
rect 3870 5328 3888 5346
rect 3870 5346 3888 5364
rect 3870 5364 3888 5382
rect 3870 5382 3888 5400
rect 3870 5400 3888 5418
rect 3870 5418 3888 5436
rect 3870 5436 3888 5454
rect 3870 5454 3888 5472
rect 3870 5472 3888 5490
rect 3870 5490 3888 5508
rect 3870 5508 3888 5526
rect 3870 5526 3888 5544
rect 3870 5544 3888 5562
rect 3870 5562 3888 5580
rect 3870 5580 3888 5598
rect 3870 5598 3888 5616
rect 3870 5616 3888 5634
rect 3870 5634 3888 5652
rect 3870 5652 3888 5670
rect 3870 5670 3888 5688
rect 3870 5688 3888 5706
rect 3870 5706 3888 5724
rect 3870 5724 3888 5742
rect 3870 5742 3888 5760
rect 3870 5760 3888 5778
rect 3870 5778 3888 5796
rect 3870 6642 3888 6660
rect 3870 6660 3888 6678
rect 3870 6678 3888 6696
rect 3870 6696 3888 6714
rect 3870 6714 3888 6732
rect 3870 6732 3888 6750
rect 3870 6750 3888 6768
rect 3870 6768 3888 6786
rect 3870 6786 3888 6804
rect 3870 6804 3888 6822
rect 3870 6822 3888 6840
rect 3870 6840 3888 6858
rect 3870 6858 3888 6876
rect 3870 6876 3888 6894
rect 3870 6894 3888 6912
rect 3870 6912 3888 6930
rect 3870 6930 3888 6948
rect 3870 6948 3888 6966
rect 3870 6966 3888 6984
rect 3870 6984 3888 7002
rect 3870 7002 3888 7020
rect 3870 7020 3888 7038
rect 3870 7038 3888 7056
rect 3870 7056 3888 7074
rect 3870 7074 3888 7092
rect 3870 7092 3888 7110
rect 3870 7110 3888 7128
rect 3870 7128 3888 7146
rect 3870 7146 3888 7164
rect 3870 7164 3888 7182
rect 3870 7182 3888 7200
rect 3870 7200 3888 7218
rect 3870 7218 3888 7236
rect 3870 7236 3888 7254
rect 3888 18 3906 36
rect 3888 36 3906 54
rect 3888 54 3906 72
rect 3888 72 3906 90
rect 3888 90 3906 108
rect 3888 108 3906 126
rect 3888 126 3906 144
rect 3888 144 3906 162
rect 3888 162 3906 180
rect 3888 180 3906 198
rect 3888 198 3906 216
rect 3888 216 3906 234
rect 3888 234 3906 252
rect 3888 252 3906 270
rect 3888 270 3906 288
rect 3888 288 3906 306
rect 3888 306 3906 324
rect 3888 324 3906 342
rect 3888 342 3906 360
rect 3888 360 3906 378
rect 3888 378 3906 396
rect 3888 396 3906 414
rect 3888 414 3906 432
rect 3888 432 3906 450
rect 3888 450 3906 468
rect 3888 468 3906 486
rect 3888 486 3906 504
rect 3888 504 3906 522
rect 3888 522 3906 540
rect 3888 540 3906 558
rect 3888 558 3906 576
rect 3888 576 3906 594
rect 3888 594 3906 612
rect 3888 612 3906 630
rect 3888 864 3906 882
rect 3888 882 3906 900
rect 3888 900 3906 918
rect 3888 918 3906 936
rect 3888 936 3906 954
rect 3888 954 3906 972
rect 3888 972 3906 990
rect 3888 990 3906 1008
rect 3888 1008 3906 1026
rect 3888 1026 3906 1044
rect 3888 1044 3906 1062
rect 3888 1062 3906 1080
rect 3888 1080 3906 1098
rect 3888 1098 3906 1116
rect 3888 1116 3906 1134
rect 3888 1134 3906 1152
rect 3888 1152 3906 1170
rect 3888 1170 3906 1188
rect 3888 1188 3906 1206
rect 3888 1206 3906 1224
rect 3888 1224 3906 1242
rect 3888 1242 3906 1260
rect 3888 1260 3906 1278
rect 3888 1278 3906 1296
rect 3888 1296 3906 1314
rect 3888 1314 3906 1332
rect 3888 1332 3906 1350
rect 3888 1350 3906 1368
rect 3888 1368 3906 1386
rect 3888 1386 3906 1404
rect 3888 1404 3906 1422
rect 3888 1422 3906 1440
rect 3888 1440 3906 1458
rect 3888 1458 3906 1476
rect 3888 1476 3906 1494
rect 3888 1728 3906 1746
rect 3888 1746 3906 1764
rect 3888 1764 3906 1782
rect 3888 1782 3906 1800
rect 3888 1800 3906 1818
rect 3888 1818 3906 1836
rect 3888 1836 3906 1854
rect 3888 1854 3906 1872
rect 3888 1872 3906 1890
rect 3888 1890 3906 1908
rect 3888 1908 3906 1926
rect 3888 1926 3906 1944
rect 3888 1944 3906 1962
rect 3888 1962 3906 1980
rect 3888 1980 3906 1998
rect 3888 1998 3906 2016
rect 3888 2016 3906 2034
rect 3888 2034 3906 2052
rect 3888 2052 3906 2070
rect 3888 2070 3906 2088
rect 3888 2088 3906 2106
rect 3888 2106 3906 2124
rect 3888 2124 3906 2142
rect 3888 2142 3906 2160
rect 3888 2160 3906 2178
rect 3888 2178 3906 2196
rect 3888 2196 3906 2214
rect 3888 2214 3906 2232
rect 3888 2232 3906 2250
rect 3888 2250 3906 2268
rect 3888 2268 3906 2286
rect 3888 2286 3906 2304
rect 3888 2304 3906 2322
rect 3888 2322 3906 2340
rect 3888 2340 3906 2358
rect 3888 2358 3906 2376
rect 3888 2376 3906 2394
rect 3888 2394 3906 2412
rect 3888 2412 3906 2430
rect 3888 2430 3906 2448
rect 3888 2448 3906 2466
rect 3888 2466 3906 2484
rect 3888 2484 3906 2502
rect 3888 2502 3906 2520
rect 3888 2520 3906 2538
rect 3888 2538 3906 2556
rect 3888 2556 3906 2574
rect 3888 2574 3906 2592
rect 3888 2592 3906 2610
rect 3888 2610 3906 2628
rect 3888 2628 3906 2646
rect 3888 2646 3906 2664
rect 3888 2664 3906 2682
rect 3888 2682 3906 2700
rect 3888 2700 3906 2718
rect 3888 2718 3906 2736
rect 3888 2736 3906 2754
rect 3888 2754 3906 2772
rect 3888 2772 3906 2790
rect 3888 2790 3906 2808
rect 3888 2808 3906 2826
rect 3888 2826 3906 2844
rect 3888 2844 3906 2862
rect 3888 2862 3906 2880
rect 3888 2880 3906 2898
rect 3888 2898 3906 2916
rect 3888 2916 3906 2934
rect 3888 3168 3906 3186
rect 3888 3186 3906 3204
rect 3888 3204 3906 3222
rect 3888 3222 3906 3240
rect 3888 3240 3906 3258
rect 3888 3258 3906 3276
rect 3888 3276 3906 3294
rect 3888 3294 3906 3312
rect 3888 3312 3906 3330
rect 3888 3330 3906 3348
rect 3888 3348 3906 3366
rect 3888 3366 3906 3384
rect 3888 3384 3906 3402
rect 3888 3402 3906 3420
rect 3888 3420 3906 3438
rect 3888 3438 3906 3456
rect 3888 3456 3906 3474
rect 3888 3474 3906 3492
rect 3888 3492 3906 3510
rect 3888 3510 3906 3528
rect 3888 3528 3906 3546
rect 3888 3546 3906 3564
rect 3888 3564 3906 3582
rect 3888 3582 3906 3600
rect 3888 3600 3906 3618
rect 3888 3618 3906 3636
rect 3888 3636 3906 3654
rect 3888 3654 3906 3672
rect 3888 3672 3906 3690
rect 3888 3690 3906 3708
rect 3888 3708 3906 3726
rect 3888 3726 3906 3744
rect 3888 3744 3906 3762
rect 3888 3762 3906 3780
rect 3888 3780 3906 3798
rect 3888 3798 3906 3816
rect 3888 3816 3906 3834
rect 3888 3834 3906 3852
rect 3888 3852 3906 3870
rect 3888 3870 3906 3888
rect 3888 3888 3906 3906
rect 3888 3906 3906 3924
rect 3888 3924 3906 3942
rect 3888 3942 3906 3960
rect 3888 3960 3906 3978
rect 3888 3978 3906 3996
rect 3888 3996 3906 4014
rect 3888 4014 3906 4032
rect 3888 4032 3906 4050
rect 3888 4050 3906 4068
rect 3888 4068 3906 4086
rect 3888 4086 3906 4104
rect 3888 4104 3906 4122
rect 3888 4122 3906 4140
rect 3888 4140 3906 4158
rect 3888 4158 3906 4176
rect 3888 4176 3906 4194
rect 3888 4194 3906 4212
rect 3888 4212 3906 4230
rect 3888 4230 3906 4248
rect 3888 4248 3906 4266
rect 3888 4266 3906 4284
rect 3888 4284 3906 4302
rect 3888 4302 3906 4320
rect 3888 4320 3906 4338
rect 3888 4338 3906 4356
rect 3888 4356 3906 4374
rect 3888 4374 3906 4392
rect 3888 4392 3906 4410
rect 3888 4410 3906 4428
rect 3888 4428 3906 4446
rect 3888 4446 3906 4464
rect 3888 4464 3906 4482
rect 3888 4482 3906 4500
rect 3888 4500 3906 4518
rect 3888 4518 3906 4536
rect 3888 4536 3906 4554
rect 3888 4554 3906 4572
rect 3888 4572 3906 4590
rect 3888 4590 3906 4608
rect 3888 4608 3906 4626
rect 3888 4626 3906 4644
rect 3888 4644 3906 4662
rect 3888 4662 3906 4680
rect 3888 4680 3906 4698
rect 3888 4698 3906 4716
rect 3888 4716 3906 4734
rect 3888 4734 3906 4752
rect 3888 4752 3906 4770
rect 3888 4770 3906 4788
rect 3888 4788 3906 4806
rect 3888 4806 3906 4824
rect 3888 4824 3906 4842
rect 3888 4842 3906 4860
rect 3888 4860 3906 4878
rect 3888 4878 3906 4896
rect 3888 4896 3906 4914
rect 3888 4914 3906 4932
rect 3888 4932 3906 4950
rect 3888 4950 3906 4968
rect 3888 4968 3906 4986
rect 3888 4986 3906 5004
rect 3888 5004 3906 5022
rect 3888 5022 3906 5040
rect 3888 5040 3906 5058
rect 3888 5058 3906 5076
rect 3888 5076 3906 5094
rect 3888 5094 3906 5112
rect 3888 5112 3906 5130
rect 3888 5130 3906 5148
rect 3888 5148 3906 5166
rect 3888 5166 3906 5184
rect 3888 5184 3906 5202
rect 3888 5202 3906 5220
rect 3888 5220 3906 5238
rect 3888 5238 3906 5256
rect 3888 5256 3906 5274
rect 3888 5274 3906 5292
rect 3888 5292 3906 5310
rect 3888 5310 3906 5328
rect 3888 5328 3906 5346
rect 3888 5346 3906 5364
rect 3888 5364 3906 5382
rect 3888 5382 3906 5400
rect 3888 5400 3906 5418
rect 3888 5418 3906 5436
rect 3888 5436 3906 5454
rect 3888 5454 3906 5472
rect 3888 5472 3906 5490
rect 3888 5490 3906 5508
rect 3888 5508 3906 5526
rect 3888 5526 3906 5544
rect 3888 5544 3906 5562
rect 3888 5562 3906 5580
rect 3888 5580 3906 5598
rect 3888 5598 3906 5616
rect 3888 5616 3906 5634
rect 3888 5634 3906 5652
rect 3888 5652 3906 5670
rect 3888 5670 3906 5688
rect 3888 5688 3906 5706
rect 3888 5706 3906 5724
rect 3888 5724 3906 5742
rect 3888 5742 3906 5760
rect 3888 5760 3906 5778
rect 3888 5778 3906 5796
rect 3888 5796 3906 5814
rect 3888 5814 3906 5832
rect 3888 5832 3906 5850
rect 3888 6642 3906 6660
rect 3888 6660 3906 6678
rect 3888 6678 3906 6696
rect 3888 6696 3906 6714
rect 3888 6714 3906 6732
rect 3888 6732 3906 6750
rect 3888 6750 3906 6768
rect 3888 6768 3906 6786
rect 3888 6786 3906 6804
rect 3888 6804 3906 6822
rect 3888 6822 3906 6840
rect 3888 6840 3906 6858
rect 3888 6858 3906 6876
rect 3888 6876 3906 6894
rect 3888 6894 3906 6912
rect 3888 6912 3906 6930
rect 3888 6930 3906 6948
rect 3888 6948 3906 6966
rect 3888 6966 3906 6984
rect 3888 6984 3906 7002
rect 3888 7002 3906 7020
rect 3888 7020 3906 7038
rect 3888 7038 3906 7056
rect 3888 7056 3906 7074
rect 3888 7074 3906 7092
rect 3888 7092 3906 7110
rect 3888 7110 3906 7128
rect 3888 7128 3906 7146
rect 3888 7146 3906 7164
rect 3888 7164 3906 7182
rect 3888 7182 3906 7200
rect 3888 7200 3906 7218
rect 3888 7218 3906 7236
rect 3888 7236 3906 7254
rect 3906 18 3924 36
rect 3906 36 3924 54
rect 3906 54 3924 72
rect 3906 72 3924 90
rect 3906 90 3924 108
rect 3906 108 3924 126
rect 3906 126 3924 144
rect 3906 144 3924 162
rect 3906 162 3924 180
rect 3906 180 3924 198
rect 3906 198 3924 216
rect 3906 216 3924 234
rect 3906 234 3924 252
rect 3906 252 3924 270
rect 3906 270 3924 288
rect 3906 288 3924 306
rect 3906 306 3924 324
rect 3906 324 3924 342
rect 3906 342 3924 360
rect 3906 360 3924 378
rect 3906 378 3924 396
rect 3906 396 3924 414
rect 3906 414 3924 432
rect 3906 432 3924 450
rect 3906 450 3924 468
rect 3906 468 3924 486
rect 3906 486 3924 504
rect 3906 504 3924 522
rect 3906 522 3924 540
rect 3906 540 3924 558
rect 3906 558 3924 576
rect 3906 576 3924 594
rect 3906 594 3924 612
rect 3906 612 3924 630
rect 3906 864 3924 882
rect 3906 882 3924 900
rect 3906 900 3924 918
rect 3906 918 3924 936
rect 3906 936 3924 954
rect 3906 954 3924 972
rect 3906 972 3924 990
rect 3906 990 3924 1008
rect 3906 1008 3924 1026
rect 3906 1026 3924 1044
rect 3906 1044 3924 1062
rect 3906 1062 3924 1080
rect 3906 1080 3924 1098
rect 3906 1098 3924 1116
rect 3906 1116 3924 1134
rect 3906 1134 3924 1152
rect 3906 1152 3924 1170
rect 3906 1170 3924 1188
rect 3906 1188 3924 1206
rect 3906 1206 3924 1224
rect 3906 1224 3924 1242
rect 3906 1242 3924 1260
rect 3906 1260 3924 1278
rect 3906 1278 3924 1296
rect 3906 1296 3924 1314
rect 3906 1314 3924 1332
rect 3906 1332 3924 1350
rect 3906 1350 3924 1368
rect 3906 1368 3924 1386
rect 3906 1386 3924 1404
rect 3906 1404 3924 1422
rect 3906 1422 3924 1440
rect 3906 1440 3924 1458
rect 3906 1458 3924 1476
rect 3906 1476 3924 1494
rect 3906 1494 3924 1512
rect 3906 1728 3924 1746
rect 3906 1746 3924 1764
rect 3906 1764 3924 1782
rect 3906 1782 3924 1800
rect 3906 1800 3924 1818
rect 3906 1818 3924 1836
rect 3906 1836 3924 1854
rect 3906 1854 3924 1872
rect 3906 1872 3924 1890
rect 3906 1890 3924 1908
rect 3906 1908 3924 1926
rect 3906 1926 3924 1944
rect 3906 1944 3924 1962
rect 3906 1962 3924 1980
rect 3906 1980 3924 1998
rect 3906 1998 3924 2016
rect 3906 2016 3924 2034
rect 3906 2034 3924 2052
rect 3906 2052 3924 2070
rect 3906 2070 3924 2088
rect 3906 2088 3924 2106
rect 3906 2106 3924 2124
rect 3906 2124 3924 2142
rect 3906 2142 3924 2160
rect 3906 2160 3924 2178
rect 3906 2178 3924 2196
rect 3906 2196 3924 2214
rect 3906 2214 3924 2232
rect 3906 2232 3924 2250
rect 3906 2250 3924 2268
rect 3906 2268 3924 2286
rect 3906 2286 3924 2304
rect 3906 2304 3924 2322
rect 3906 2322 3924 2340
rect 3906 2340 3924 2358
rect 3906 2358 3924 2376
rect 3906 2376 3924 2394
rect 3906 2394 3924 2412
rect 3906 2412 3924 2430
rect 3906 2430 3924 2448
rect 3906 2448 3924 2466
rect 3906 2466 3924 2484
rect 3906 2484 3924 2502
rect 3906 2502 3924 2520
rect 3906 2520 3924 2538
rect 3906 2538 3924 2556
rect 3906 2556 3924 2574
rect 3906 2574 3924 2592
rect 3906 2592 3924 2610
rect 3906 2610 3924 2628
rect 3906 2628 3924 2646
rect 3906 2646 3924 2664
rect 3906 2664 3924 2682
rect 3906 2682 3924 2700
rect 3906 2700 3924 2718
rect 3906 2718 3924 2736
rect 3906 2736 3924 2754
rect 3906 2754 3924 2772
rect 3906 2772 3924 2790
rect 3906 2790 3924 2808
rect 3906 2808 3924 2826
rect 3906 2826 3924 2844
rect 3906 2844 3924 2862
rect 3906 2862 3924 2880
rect 3906 2880 3924 2898
rect 3906 2898 3924 2916
rect 3906 2916 3924 2934
rect 3906 2934 3924 2952
rect 3906 3204 3924 3222
rect 3906 3222 3924 3240
rect 3906 3240 3924 3258
rect 3906 3258 3924 3276
rect 3906 3276 3924 3294
rect 3906 3294 3924 3312
rect 3906 3312 3924 3330
rect 3906 3330 3924 3348
rect 3906 3348 3924 3366
rect 3906 3366 3924 3384
rect 3906 3384 3924 3402
rect 3906 3402 3924 3420
rect 3906 3420 3924 3438
rect 3906 3438 3924 3456
rect 3906 3456 3924 3474
rect 3906 3474 3924 3492
rect 3906 3492 3924 3510
rect 3906 3510 3924 3528
rect 3906 3528 3924 3546
rect 3906 3546 3924 3564
rect 3906 3564 3924 3582
rect 3906 3582 3924 3600
rect 3906 3600 3924 3618
rect 3906 3618 3924 3636
rect 3906 3636 3924 3654
rect 3906 3654 3924 3672
rect 3906 3672 3924 3690
rect 3906 3690 3924 3708
rect 3906 3708 3924 3726
rect 3906 3726 3924 3744
rect 3906 3744 3924 3762
rect 3906 3762 3924 3780
rect 3906 3780 3924 3798
rect 3906 3798 3924 3816
rect 3906 3816 3924 3834
rect 3906 3834 3924 3852
rect 3906 3852 3924 3870
rect 3906 3870 3924 3888
rect 3906 3888 3924 3906
rect 3906 3906 3924 3924
rect 3906 3924 3924 3942
rect 3906 3942 3924 3960
rect 3906 3960 3924 3978
rect 3906 3978 3924 3996
rect 3906 3996 3924 4014
rect 3906 4014 3924 4032
rect 3906 4032 3924 4050
rect 3906 4050 3924 4068
rect 3906 4068 3924 4086
rect 3906 4086 3924 4104
rect 3906 4104 3924 4122
rect 3906 4122 3924 4140
rect 3906 4140 3924 4158
rect 3906 4158 3924 4176
rect 3906 4176 3924 4194
rect 3906 4194 3924 4212
rect 3906 4212 3924 4230
rect 3906 4230 3924 4248
rect 3906 4248 3924 4266
rect 3906 4266 3924 4284
rect 3906 4284 3924 4302
rect 3906 4302 3924 4320
rect 3906 4320 3924 4338
rect 3906 4338 3924 4356
rect 3906 4356 3924 4374
rect 3906 4374 3924 4392
rect 3906 4392 3924 4410
rect 3906 4410 3924 4428
rect 3906 4428 3924 4446
rect 3906 4446 3924 4464
rect 3906 4464 3924 4482
rect 3906 4482 3924 4500
rect 3906 4500 3924 4518
rect 3906 4518 3924 4536
rect 3906 4536 3924 4554
rect 3906 4554 3924 4572
rect 3906 4572 3924 4590
rect 3906 4590 3924 4608
rect 3906 4608 3924 4626
rect 3906 4626 3924 4644
rect 3906 4644 3924 4662
rect 3906 4662 3924 4680
rect 3906 4680 3924 4698
rect 3906 4698 3924 4716
rect 3906 4716 3924 4734
rect 3906 4734 3924 4752
rect 3906 4752 3924 4770
rect 3906 4770 3924 4788
rect 3906 4788 3924 4806
rect 3906 4806 3924 4824
rect 3906 4824 3924 4842
rect 3906 4842 3924 4860
rect 3906 4860 3924 4878
rect 3906 4878 3924 4896
rect 3906 4896 3924 4914
rect 3906 4914 3924 4932
rect 3906 4932 3924 4950
rect 3906 4950 3924 4968
rect 3906 4968 3924 4986
rect 3906 4986 3924 5004
rect 3906 5004 3924 5022
rect 3906 5022 3924 5040
rect 3906 5040 3924 5058
rect 3906 5058 3924 5076
rect 3906 5076 3924 5094
rect 3906 5094 3924 5112
rect 3906 5112 3924 5130
rect 3906 5130 3924 5148
rect 3906 5148 3924 5166
rect 3906 5166 3924 5184
rect 3906 5184 3924 5202
rect 3906 5202 3924 5220
rect 3906 5220 3924 5238
rect 3906 5238 3924 5256
rect 3906 5256 3924 5274
rect 3906 5274 3924 5292
rect 3906 5292 3924 5310
rect 3906 5310 3924 5328
rect 3906 5328 3924 5346
rect 3906 5346 3924 5364
rect 3906 5364 3924 5382
rect 3906 5382 3924 5400
rect 3906 5400 3924 5418
rect 3906 5418 3924 5436
rect 3906 5436 3924 5454
rect 3906 5454 3924 5472
rect 3906 5472 3924 5490
rect 3906 5490 3924 5508
rect 3906 5508 3924 5526
rect 3906 5526 3924 5544
rect 3906 5544 3924 5562
rect 3906 5562 3924 5580
rect 3906 5580 3924 5598
rect 3906 5598 3924 5616
rect 3906 5616 3924 5634
rect 3906 5634 3924 5652
rect 3906 5652 3924 5670
rect 3906 5670 3924 5688
rect 3906 5688 3924 5706
rect 3906 5706 3924 5724
rect 3906 5724 3924 5742
rect 3906 5742 3924 5760
rect 3906 5760 3924 5778
rect 3906 5778 3924 5796
rect 3906 5796 3924 5814
rect 3906 5814 3924 5832
rect 3906 5832 3924 5850
rect 3906 5850 3924 5868
rect 3906 5868 3924 5886
rect 3906 6642 3924 6660
rect 3906 6660 3924 6678
rect 3906 6678 3924 6696
rect 3906 6696 3924 6714
rect 3906 6714 3924 6732
rect 3906 6732 3924 6750
rect 3906 6750 3924 6768
rect 3906 6768 3924 6786
rect 3906 6786 3924 6804
rect 3906 6804 3924 6822
rect 3906 6822 3924 6840
rect 3906 6840 3924 6858
rect 3906 6858 3924 6876
rect 3906 6876 3924 6894
rect 3906 6894 3924 6912
rect 3906 6912 3924 6930
rect 3906 6930 3924 6948
rect 3906 6948 3924 6966
rect 3906 6966 3924 6984
rect 3906 6984 3924 7002
rect 3906 7002 3924 7020
rect 3906 7020 3924 7038
rect 3906 7038 3924 7056
rect 3906 7056 3924 7074
rect 3906 7074 3924 7092
rect 3906 7092 3924 7110
rect 3906 7110 3924 7128
rect 3906 7128 3924 7146
rect 3906 7146 3924 7164
rect 3906 7164 3924 7182
rect 3906 7182 3924 7200
rect 3906 7200 3924 7218
rect 3906 7218 3924 7236
rect 3906 7236 3924 7254
rect 3924 18 3942 36
rect 3924 36 3942 54
rect 3924 54 3942 72
rect 3924 72 3942 90
rect 3924 90 3942 108
rect 3924 108 3942 126
rect 3924 126 3942 144
rect 3924 144 3942 162
rect 3924 162 3942 180
rect 3924 180 3942 198
rect 3924 198 3942 216
rect 3924 216 3942 234
rect 3924 234 3942 252
rect 3924 252 3942 270
rect 3924 270 3942 288
rect 3924 288 3942 306
rect 3924 306 3942 324
rect 3924 324 3942 342
rect 3924 342 3942 360
rect 3924 360 3942 378
rect 3924 378 3942 396
rect 3924 396 3942 414
rect 3924 414 3942 432
rect 3924 432 3942 450
rect 3924 450 3942 468
rect 3924 468 3942 486
rect 3924 486 3942 504
rect 3924 504 3942 522
rect 3924 522 3942 540
rect 3924 540 3942 558
rect 3924 558 3942 576
rect 3924 576 3942 594
rect 3924 594 3942 612
rect 3924 612 3942 630
rect 3924 864 3942 882
rect 3924 882 3942 900
rect 3924 900 3942 918
rect 3924 918 3942 936
rect 3924 936 3942 954
rect 3924 954 3942 972
rect 3924 972 3942 990
rect 3924 990 3942 1008
rect 3924 1008 3942 1026
rect 3924 1026 3942 1044
rect 3924 1044 3942 1062
rect 3924 1062 3942 1080
rect 3924 1080 3942 1098
rect 3924 1098 3942 1116
rect 3924 1116 3942 1134
rect 3924 1134 3942 1152
rect 3924 1152 3942 1170
rect 3924 1170 3942 1188
rect 3924 1188 3942 1206
rect 3924 1206 3942 1224
rect 3924 1224 3942 1242
rect 3924 1242 3942 1260
rect 3924 1260 3942 1278
rect 3924 1278 3942 1296
rect 3924 1296 3942 1314
rect 3924 1314 3942 1332
rect 3924 1332 3942 1350
rect 3924 1350 3942 1368
rect 3924 1368 3942 1386
rect 3924 1386 3942 1404
rect 3924 1404 3942 1422
rect 3924 1422 3942 1440
rect 3924 1440 3942 1458
rect 3924 1458 3942 1476
rect 3924 1476 3942 1494
rect 3924 1494 3942 1512
rect 3924 1746 3942 1764
rect 3924 1764 3942 1782
rect 3924 1782 3942 1800
rect 3924 1800 3942 1818
rect 3924 1818 3942 1836
rect 3924 1836 3942 1854
rect 3924 1854 3942 1872
rect 3924 1872 3942 1890
rect 3924 1890 3942 1908
rect 3924 1908 3942 1926
rect 3924 1926 3942 1944
rect 3924 1944 3942 1962
rect 3924 1962 3942 1980
rect 3924 1980 3942 1998
rect 3924 1998 3942 2016
rect 3924 2016 3942 2034
rect 3924 2034 3942 2052
rect 3924 2052 3942 2070
rect 3924 2070 3942 2088
rect 3924 2088 3942 2106
rect 3924 2106 3942 2124
rect 3924 2124 3942 2142
rect 3924 2142 3942 2160
rect 3924 2160 3942 2178
rect 3924 2178 3942 2196
rect 3924 2196 3942 2214
rect 3924 2214 3942 2232
rect 3924 2232 3942 2250
rect 3924 2250 3942 2268
rect 3924 2268 3942 2286
rect 3924 2286 3942 2304
rect 3924 2304 3942 2322
rect 3924 2322 3942 2340
rect 3924 2340 3942 2358
rect 3924 2358 3942 2376
rect 3924 2376 3942 2394
rect 3924 2394 3942 2412
rect 3924 2412 3942 2430
rect 3924 2430 3942 2448
rect 3924 2448 3942 2466
rect 3924 2466 3942 2484
rect 3924 2484 3942 2502
rect 3924 2502 3942 2520
rect 3924 2520 3942 2538
rect 3924 2538 3942 2556
rect 3924 2556 3942 2574
rect 3924 2574 3942 2592
rect 3924 2592 3942 2610
rect 3924 2610 3942 2628
rect 3924 2628 3942 2646
rect 3924 2646 3942 2664
rect 3924 2664 3942 2682
rect 3924 2682 3942 2700
rect 3924 2700 3942 2718
rect 3924 2718 3942 2736
rect 3924 2736 3942 2754
rect 3924 2754 3942 2772
rect 3924 2772 3942 2790
rect 3924 2790 3942 2808
rect 3924 2808 3942 2826
rect 3924 2826 3942 2844
rect 3924 2844 3942 2862
rect 3924 2862 3942 2880
rect 3924 2880 3942 2898
rect 3924 2898 3942 2916
rect 3924 2916 3942 2934
rect 3924 2934 3942 2952
rect 3924 2952 3942 2970
rect 3924 2970 3942 2988
rect 3924 3222 3942 3240
rect 3924 3240 3942 3258
rect 3924 3258 3942 3276
rect 3924 3276 3942 3294
rect 3924 3294 3942 3312
rect 3924 3312 3942 3330
rect 3924 3330 3942 3348
rect 3924 3348 3942 3366
rect 3924 3366 3942 3384
rect 3924 3384 3942 3402
rect 3924 3402 3942 3420
rect 3924 3420 3942 3438
rect 3924 3438 3942 3456
rect 3924 3456 3942 3474
rect 3924 3474 3942 3492
rect 3924 3492 3942 3510
rect 3924 3510 3942 3528
rect 3924 3528 3942 3546
rect 3924 3546 3942 3564
rect 3924 3564 3942 3582
rect 3924 3582 3942 3600
rect 3924 3600 3942 3618
rect 3924 3618 3942 3636
rect 3924 3636 3942 3654
rect 3924 3654 3942 3672
rect 3924 3672 3942 3690
rect 3924 3690 3942 3708
rect 3924 3708 3942 3726
rect 3924 3726 3942 3744
rect 3924 3744 3942 3762
rect 3924 3762 3942 3780
rect 3924 3780 3942 3798
rect 3924 3798 3942 3816
rect 3924 3816 3942 3834
rect 3924 3834 3942 3852
rect 3924 3852 3942 3870
rect 3924 3870 3942 3888
rect 3924 3888 3942 3906
rect 3924 3906 3942 3924
rect 3924 3924 3942 3942
rect 3924 3942 3942 3960
rect 3924 3960 3942 3978
rect 3924 3978 3942 3996
rect 3924 3996 3942 4014
rect 3924 4014 3942 4032
rect 3924 4032 3942 4050
rect 3924 4050 3942 4068
rect 3924 4068 3942 4086
rect 3924 4086 3942 4104
rect 3924 4104 3942 4122
rect 3924 4122 3942 4140
rect 3924 4140 3942 4158
rect 3924 4158 3942 4176
rect 3924 4176 3942 4194
rect 3924 4194 3942 4212
rect 3924 4212 3942 4230
rect 3924 4230 3942 4248
rect 3924 4248 3942 4266
rect 3924 4266 3942 4284
rect 3924 4284 3942 4302
rect 3924 4302 3942 4320
rect 3924 4320 3942 4338
rect 3924 4338 3942 4356
rect 3924 4356 3942 4374
rect 3924 4374 3942 4392
rect 3924 4392 3942 4410
rect 3924 4410 3942 4428
rect 3924 4428 3942 4446
rect 3924 4446 3942 4464
rect 3924 4464 3942 4482
rect 3924 4482 3942 4500
rect 3924 4500 3942 4518
rect 3924 4518 3942 4536
rect 3924 4536 3942 4554
rect 3924 4554 3942 4572
rect 3924 4572 3942 4590
rect 3924 4590 3942 4608
rect 3924 4608 3942 4626
rect 3924 4626 3942 4644
rect 3924 4644 3942 4662
rect 3924 4662 3942 4680
rect 3924 4680 3942 4698
rect 3924 4698 3942 4716
rect 3924 4716 3942 4734
rect 3924 4734 3942 4752
rect 3924 4752 3942 4770
rect 3924 4770 3942 4788
rect 3924 4788 3942 4806
rect 3924 4806 3942 4824
rect 3924 4824 3942 4842
rect 3924 4842 3942 4860
rect 3924 4860 3942 4878
rect 3924 4878 3942 4896
rect 3924 4896 3942 4914
rect 3924 4914 3942 4932
rect 3924 4932 3942 4950
rect 3924 4950 3942 4968
rect 3924 4968 3942 4986
rect 3924 4986 3942 5004
rect 3924 5004 3942 5022
rect 3924 5022 3942 5040
rect 3924 5040 3942 5058
rect 3924 5058 3942 5076
rect 3924 5076 3942 5094
rect 3924 5094 3942 5112
rect 3924 5112 3942 5130
rect 3924 5130 3942 5148
rect 3924 5148 3942 5166
rect 3924 5166 3942 5184
rect 3924 5184 3942 5202
rect 3924 5202 3942 5220
rect 3924 5220 3942 5238
rect 3924 5238 3942 5256
rect 3924 5256 3942 5274
rect 3924 5274 3942 5292
rect 3924 5292 3942 5310
rect 3924 5310 3942 5328
rect 3924 5328 3942 5346
rect 3924 5346 3942 5364
rect 3924 5364 3942 5382
rect 3924 5382 3942 5400
rect 3924 5400 3942 5418
rect 3924 5418 3942 5436
rect 3924 5436 3942 5454
rect 3924 5454 3942 5472
rect 3924 5472 3942 5490
rect 3924 5490 3942 5508
rect 3924 5508 3942 5526
rect 3924 5526 3942 5544
rect 3924 5544 3942 5562
rect 3924 5562 3942 5580
rect 3924 5580 3942 5598
rect 3924 5598 3942 5616
rect 3924 5616 3942 5634
rect 3924 5634 3942 5652
rect 3924 5652 3942 5670
rect 3924 5670 3942 5688
rect 3924 5688 3942 5706
rect 3924 5706 3942 5724
rect 3924 5724 3942 5742
rect 3924 5742 3942 5760
rect 3924 5760 3942 5778
rect 3924 5778 3942 5796
rect 3924 5796 3942 5814
rect 3924 5814 3942 5832
rect 3924 5832 3942 5850
rect 3924 5850 3942 5868
rect 3924 5868 3942 5886
rect 3924 5886 3942 5904
rect 3924 5904 3942 5922
rect 3924 6642 3942 6660
rect 3924 6660 3942 6678
rect 3924 6678 3942 6696
rect 3924 6696 3942 6714
rect 3924 6714 3942 6732
rect 3924 6732 3942 6750
rect 3924 6750 3942 6768
rect 3924 6768 3942 6786
rect 3924 6786 3942 6804
rect 3924 6804 3942 6822
rect 3924 6822 3942 6840
rect 3924 6840 3942 6858
rect 3924 6858 3942 6876
rect 3924 6876 3942 6894
rect 3924 6894 3942 6912
rect 3924 6912 3942 6930
rect 3924 6930 3942 6948
rect 3924 6948 3942 6966
rect 3924 6966 3942 6984
rect 3924 6984 3942 7002
rect 3924 7002 3942 7020
rect 3924 7020 3942 7038
rect 3924 7038 3942 7056
rect 3924 7056 3942 7074
rect 3924 7074 3942 7092
rect 3924 7092 3942 7110
rect 3924 7110 3942 7128
rect 3924 7128 3942 7146
rect 3924 7146 3942 7164
rect 3924 7164 3942 7182
rect 3924 7182 3942 7200
rect 3924 7200 3942 7218
rect 3924 7218 3942 7236
rect 3924 7236 3942 7254
rect 3942 18 3960 36
rect 3942 36 3960 54
rect 3942 54 3960 72
rect 3942 72 3960 90
rect 3942 90 3960 108
rect 3942 108 3960 126
rect 3942 126 3960 144
rect 3942 144 3960 162
rect 3942 162 3960 180
rect 3942 180 3960 198
rect 3942 198 3960 216
rect 3942 216 3960 234
rect 3942 234 3960 252
rect 3942 252 3960 270
rect 3942 270 3960 288
rect 3942 288 3960 306
rect 3942 306 3960 324
rect 3942 324 3960 342
rect 3942 342 3960 360
rect 3942 360 3960 378
rect 3942 378 3960 396
rect 3942 396 3960 414
rect 3942 414 3960 432
rect 3942 432 3960 450
rect 3942 450 3960 468
rect 3942 468 3960 486
rect 3942 486 3960 504
rect 3942 504 3960 522
rect 3942 522 3960 540
rect 3942 540 3960 558
rect 3942 558 3960 576
rect 3942 576 3960 594
rect 3942 594 3960 612
rect 3942 612 3960 630
rect 3942 864 3960 882
rect 3942 882 3960 900
rect 3942 900 3960 918
rect 3942 918 3960 936
rect 3942 936 3960 954
rect 3942 954 3960 972
rect 3942 972 3960 990
rect 3942 990 3960 1008
rect 3942 1008 3960 1026
rect 3942 1026 3960 1044
rect 3942 1044 3960 1062
rect 3942 1062 3960 1080
rect 3942 1080 3960 1098
rect 3942 1098 3960 1116
rect 3942 1116 3960 1134
rect 3942 1134 3960 1152
rect 3942 1152 3960 1170
rect 3942 1170 3960 1188
rect 3942 1188 3960 1206
rect 3942 1206 3960 1224
rect 3942 1224 3960 1242
rect 3942 1242 3960 1260
rect 3942 1260 3960 1278
rect 3942 1278 3960 1296
rect 3942 1296 3960 1314
rect 3942 1314 3960 1332
rect 3942 1332 3960 1350
rect 3942 1350 3960 1368
rect 3942 1368 3960 1386
rect 3942 1386 3960 1404
rect 3942 1404 3960 1422
rect 3942 1422 3960 1440
rect 3942 1440 3960 1458
rect 3942 1458 3960 1476
rect 3942 1476 3960 1494
rect 3942 1494 3960 1512
rect 3942 1512 3960 1530
rect 3942 1764 3960 1782
rect 3942 1782 3960 1800
rect 3942 1800 3960 1818
rect 3942 1818 3960 1836
rect 3942 1836 3960 1854
rect 3942 1854 3960 1872
rect 3942 1872 3960 1890
rect 3942 1890 3960 1908
rect 3942 1908 3960 1926
rect 3942 1926 3960 1944
rect 3942 1944 3960 1962
rect 3942 1962 3960 1980
rect 3942 1980 3960 1998
rect 3942 1998 3960 2016
rect 3942 2016 3960 2034
rect 3942 2034 3960 2052
rect 3942 2052 3960 2070
rect 3942 2070 3960 2088
rect 3942 2088 3960 2106
rect 3942 2106 3960 2124
rect 3942 2124 3960 2142
rect 3942 2142 3960 2160
rect 3942 2160 3960 2178
rect 3942 2178 3960 2196
rect 3942 2196 3960 2214
rect 3942 2214 3960 2232
rect 3942 2232 3960 2250
rect 3942 2250 3960 2268
rect 3942 2268 3960 2286
rect 3942 2286 3960 2304
rect 3942 2304 3960 2322
rect 3942 2322 3960 2340
rect 3942 2340 3960 2358
rect 3942 2358 3960 2376
rect 3942 2376 3960 2394
rect 3942 2394 3960 2412
rect 3942 2412 3960 2430
rect 3942 2430 3960 2448
rect 3942 2448 3960 2466
rect 3942 2466 3960 2484
rect 3942 2484 3960 2502
rect 3942 2502 3960 2520
rect 3942 2520 3960 2538
rect 3942 2538 3960 2556
rect 3942 2556 3960 2574
rect 3942 2574 3960 2592
rect 3942 2592 3960 2610
rect 3942 2610 3960 2628
rect 3942 2628 3960 2646
rect 3942 2646 3960 2664
rect 3942 2664 3960 2682
rect 3942 2682 3960 2700
rect 3942 2700 3960 2718
rect 3942 2718 3960 2736
rect 3942 2736 3960 2754
rect 3942 2754 3960 2772
rect 3942 2772 3960 2790
rect 3942 2790 3960 2808
rect 3942 2808 3960 2826
rect 3942 2826 3960 2844
rect 3942 2844 3960 2862
rect 3942 2862 3960 2880
rect 3942 2880 3960 2898
rect 3942 2898 3960 2916
rect 3942 2916 3960 2934
rect 3942 2934 3960 2952
rect 3942 2952 3960 2970
rect 3942 2970 3960 2988
rect 3942 2988 3960 3006
rect 3942 3240 3960 3258
rect 3942 3258 3960 3276
rect 3942 3276 3960 3294
rect 3942 3294 3960 3312
rect 3942 3312 3960 3330
rect 3942 3330 3960 3348
rect 3942 3348 3960 3366
rect 3942 3366 3960 3384
rect 3942 3384 3960 3402
rect 3942 3402 3960 3420
rect 3942 3420 3960 3438
rect 3942 3438 3960 3456
rect 3942 3456 3960 3474
rect 3942 3474 3960 3492
rect 3942 3492 3960 3510
rect 3942 3510 3960 3528
rect 3942 3528 3960 3546
rect 3942 3546 3960 3564
rect 3942 3564 3960 3582
rect 3942 3582 3960 3600
rect 3942 3600 3960 3618
rect 3942 3618 3960 3636
rect 3942 3636 3960 3654
rect 3942 3654 3960 3672
rect 3942 3672 3960 3690
rect 3942 3690 3960 3708
rect 3942 3708 3960 3726
rect 3942 3726 3960 3744
rect 3942 3744 3960 3762
rect 3942 3762 3960 3780
rect 3942 3780 3960 3798
rect 3942 3798 3960 3816
rect 3942 3816 3960 3834
rect 3942 3834 3960 3852
rect 3942 3852 3960 3870
rect 3942 3870 3960 3888
rect 3942 3888 3960 3906
rect 3942 3906 3960 3924
rect 3942 3924 3960 3942
rect 3942 3942 3960 3960
rect 3942 3960 3960 3978
rect 3942 3978 3960 3996
rect 3942 3996 3960 4014
rect 3942 4014 3960 4032
rect 3942 4032 3960 4050
rect 3942 4050 3960 4068
rect 3942 4068 3960 4086
rect 3942 4086 3960 4104
rect 3942 4104 3960 4122
rect 3942 4122 3960 4140
rect 3942 4140 3960 4158
rect 3942 4158 3960 4176
rect 3942 4176 3960 4194
rect 3942 4194 3960 4212
rect 3942 4212 3960 4230
rect 3942 4230 3960 4248
rect 3942 4248 3960 4266
rect 3942 4266 3960 4284
rect 3942 4284 3960 4302
rect 3942 4302 3960 4320
rect 3942 4320 3960 4338
rect 3942 4338 3960 4356
rect 3942 4356 3960 4374
rect 3942 4374 3960 4392
rect 3942 4392 3960 4410
rect 3942 4410 3960 4428
rect 3942 4428 3960 4446
rect 3942 4446 3960 4464
rect 3942 4464 3960 4482
rect 3942 4482 3960 4500
rect 3942 4500 3960 4518
rect 3942 4518 3960 4536
rect 3942 4536 3960 4554
rect 3942 4554 3960 4572
rect 3942 4572 3960 4590
rect 3942 4590 3960 4608
rect 3942 4608 3960 4626
rect 3942 4626 3960 4644
rect 3942 4644 3960 4662
rect 3942 4662 3960 4680
rect 3942 4680 3960 4698
rect 3942 4698 3960 4716
rect 3942 4716 3960 4734
rect 3942 4734 3960 4752
rect 3942 4752 3960 4770
rect 3942 4770 3960 4788
rect 3942 4788 3960 4806
rect 3942 4806 3960 4824
rect 3942 4824 3960 4842
rect 3942 4842 3960 4860
rect 3942 4860 3960 4878
rect 3942 4878 3960 4896
rect 3942 4896 3960 4914
rect 3942 4914 3960 4932
rect 3942 4932 3960 4950
rect 3942 4950 3960 4968
rect 3942 4968 3960 4986
rect 3942 4986 3960 5004
rect 3942 5004 3960 5022
rect 3942 5022 3960 5040
rect 3942 5040 3960 5058
rect 3942 5058 3960 5076
rect 3942 5076 3960 5094
rect 3942 5094 3960 5112
rect 3942 5112 3960 5130
rect 3942 5130 3960 5148
rect 3942 5148 3960 5166
rect 3942 5166 3960 5184
rect 3942 5184 3960 5202
rect 3942 5202 3960 5220
rect 3942 5220 3960 5238
rect 3942 5238 3960 5256
rect 3942 5256 3960 5274
rect 3942 5274 3960 5292
rect 3942 5292 3960 5310
rect 3942 5310 3960 5328
rect 3942 5328 3960 5346
rect 3942 5346 3960 5364
rect 3942 5364 3960 5382
rect 3942 5382 3960 5400
rect 3942 5400 3960 5418
rect 3942 5418 3960 5436
rect 3942 5436 3960 5454
rect 3942 5454 3960 5472
rect 3942 5472 3960 5490
rect 3942 5490 3960 5508
rect 3942 5508 3960 5526
rect 3942 5526 3960 5544
rect 3942 5544 3960 5562
rect 3942 5562 3960 5580
rect 3942 5580 3960 5598
rect 3942 5598 3960 5616
rect 3942 5616 3960 5634
rect 3942 5634 3960 5652
rect 3942 5652 3960 5670
rect 3942 5670 3960 5688
rect 3942 5688 3960 5706
rect 3942 5706 3960 5724
rect 3942 5724 3960 5742
rect 3942 5742 3960 5760
rect 3942 5760 3960 5778
rect 3942 5778 3960 5796
rect 3942 5796 3960 5814
rect 3942 5814 3960 5832
rect 3942 5832 3960 5850
rect 3942 5850 3960 5868
rect 3942 5868 3960 5886
rect 3942 5886 3960 5904
rect 3942 5904 3960 5922
rect 3942 5922 3960 5940
rect 3942 5940 3960 5958
rect 3942 6642 3960 6660
rect 3942 6660 3960 6678
rect 3942 6678 3960 6696
rect 3942 6696 3960 6714
rect 3942 6714 3960 6732
rect 3942 6732 3960 6750
rect 3942 6750 3960 6768
rect 3942 6768 3960 6786
rect 3942 6786 3960 6804
rect 3942 6804 3960 6822
rect 3942 6822 3960 6840
rect 3942 6840 3960 6858
rect 3942 6858 3960 6876
rect 3942 6876 3960 6894
rect 3942 6894 3960 6912
rect 3942 6912 3960 6930
rect 3942 6930 3960 6948
rect 3942 6948 3960 6966
rect 3942 6966 3960 6984
rect 3942 6984 3960 7002
rect 3942 7002 3960 7020
rect 3942 7020 3960 7038
rect 3942 7038 3960 7056
rect 3942 7056 3960 7074
rect 3942 7074 3960 7092
rect 3942 7092 3960 7110
rect 3942 7110 3960 7128
rect 3942 7128 3960 7146
rect 3942 7146 3960 7164
rect 3942 7164 3960 7182
rect 3942 7182 3960 7200
rect 3942 7200 3960 7218
rect 3942 7218 3960 7236
rect 3942 7236 3960 7254
rect 3960 18 3978 36
rect 3960 36 3978 54
rect 3960 54 3978 72
rect 3960 72 3978 90
rect 3960 90 3978 108
rect 3960 108 3978 126
rect 3960 126 3978 144
rect 3960 144 3978 162
rect 3960 162 3978 180
rect 3960 180 3978 198
rect 3960 198 3978 216
rect 3960 216 3978 234
rect 3960 234 3978 252
rect 3960 252 3978 270
rect 3960 270 3978 288
rect 3960 288 3978 306
rect 3960 306 3978 324
rect 3960 324 3978 342
rect 3960 342 3978 360
rect 3960 360 3978 378
rect 3960 378 3978 396
rect 3960 396 3978 414
rect 3960 414 3978 432
rect 3960 432 3978 450
rect 3960 450 3978 468
rect 3960 468 3978 486
rect 3960 486 3978 504
rect 3960 504 3978 522
rect 3960 522 3978 540
rect 3960 540 3978 558
rect 3960 558 3978 576
rect 3960 576 3978 594
rect 3960 594 3978 612
rect 3960 612 3978 630
rect 3960 864 3978 882
rect 3960 882 3978 900
rect 3960 900 3978 918
rect 3960 918 3978 936
rect 3960 936 3978 954
rect 3960 954 3978 972
rect 3960 972 3978 990
rect 3960 990 3978 1008
rect 3960 1008 3978 1026
rect 3960 1026 3978 1044
rect 3960 1044 3978 1062
rect 3960 1062 3978 1080
rect 3960 1080 3978 1098
rect 3960 1098 3978 1116
rect 3960 1116 3978 1134
rect 3960 1134 3978 1152
rect 3960 1152 3978 1170
rect 3960 1170 3978 1188
rect 3960 1188 3978 1206
rect 3960 1206 3978 1224
rect 3960 1224 3978 1242
rect 3960 1242 3978 1260
rect 3960 1260 3978 1278
rect 3960 1278 3978 1296
rect 3960 1296 3978 1314
rect 3960 1314 3978 1332
rect 3960 1332 3978 1350
rect 3960 1350 3978 1368
rect 3960 1368 3978 1386
rect 3960 1386 3978 1404
rect 3960 1404 3978 1422
rect 3960 1422 3978 1440
rect 3960 1440 3978 1458
rect 3960 1458 3978 1476
rect 3960 1476 3978 1494
rect 3960 1494 3978 1512
rect 3960 1512 3978 1530
rect 3960 1530 3978 1548
rect 3960 1782 3978 1800
rect 3960 1800 3978 1818
rect 3960 1818 3978 1836
rect 3960 1836 3978 1854
rect 3960 1854 3978 1872
rect 3960 1872 3978 1890
rect 3960 1890 3978 1908
rect 3960 1908 3978 1926
rect 3960 1926 3978 1944
rect 3960 1944 3978 1962
rect 3960 1962 3978 1980
rect 3960 1980 3978 1998
rect 3960 1998 3978 2016
rect 3960 2016 3978 2034
rect 3960 2034 3978 2052
rect 3960 2052 3978 2070
rect 3960 2070 3978 2088
rect 3960 2088 3978 2106
rect 3960 2106 3978 2124
rect 3960 2124 3978 2142
rect 3960 2142 3978 2160
rect 3960 2160 3978 2178
rect 3960 2178 3978 2196
rect 3960 2196 3978 2214
rect 3960 2214 3978 2232
rect 3960 2232 3978 2250
rect 3960 2250 3978 2268
rect 3960 2268 3978 2286
rect 3960 2286 3978 2304
rect 3960 2304 3978 2322
rect 3960 2322 3978 2340
rect 3960 2340 3978 2358
rect 3960 2358 3978 2376
rect 3960 2376 3978 2394
rect 3960 2394 3978 2412
rect 3960 2412 3978 2430
rect 3960 2430 3978 2448
rect 3960 2448 3978 2466
rect 3960 2466 3978 2484
rect 3960 2484 3978 2502
rect 3960 2502 3978 2520
rect 3960 2520 3978 2538
rect 3960 2538 3978 2556
rect 3960 2556 3978 2574
rect 3960 2574 3978 2592
rect 3960 2592 3978 2610
rect 3960 2610 3978 2628
rect 3960 2628 3978 2646
rect 3960 2646 3978 2664
rect 3960 2664 3978 2682
rect 3960 2682 3978 2700
rect 3960 2700 3978 2718
rect 3960 2718 3978 2736
rect 3960 2736 3978 2754
rect 3960 2754 3978 2772
rect 3960 2772 3978 2790
rect 3960 2790 3978 2808
rect 3960 2808 3978 2826
rect 3960 2826 3978 2844
rect 3960 2844 3978 2862
rect 3960 2862 3978 2880
rect 3960 2880 3978 2898
rect 3960 2898 3978 2916
rect 3960 2916 3978 2934
rect 3960 2934 3978 2952
rect 3960 2952 3978 2970
rect 3960 2970 3978 2988
rect 3960 2988 3978 3006
rect 3960 3006 3978 3024
rect 3960 3024 3978 3042
rect 3960 3276 3978 3294
rect 3960 3294 3978 3312
rect 3960 3312 3978 3330
rect 3960 3330 3978 3348
rect 3960 3348 3978 3366
rect 3960 3366 3978 3384
rect 3960 3384 3978 3402
rect 3960 3402 3978 3420
rect 3960 3420 3978 3438
rect 3960 3438 3978 3456
rect 3960 3456 3978 3474
rect 3960 3474 3978 3492
rect 3960 3492 3978 3510
rect 3960 3510 3978 3528
rect 3960 3528 3978 3546
rect 3960 3546 3978 3564
rect 3960 3564 3978 3582
rect 3960 3582 3978 3600
rect 3960 3600 3978 3618
rect 3960 3618 3978 3636
rect 3960 3636 3978 3654
rect 3960 3654 3978 3672
rect 3960 3672 3978 3690
rect 3960 3690 3978 3708
rect 3960 3708 3978 3726
rect 3960 3726 3978 3744
rect 3960 3744 3978 3762
rect 3960 3762 3978 3780
rect 3960 3780 3978 3798
rect 3960 3798 3978 3816
rect 3960 3816 3978 3834
rect 3960 3834 3978 3852
rect 3960 3852 3978 3870
rect 3960 3870 3978 3888
rect 3960 3888 3978 3906
rect 3960 3906 3978 3924
rect 3960 3924 3978 3942
rect 3960 3942 3978 3960
rect 3960 3960 3978 3978
rect 3960 3978 3978 3996
rect 3960 3996 3978 4014
rect 3960 4014 3978 4032
rect 3960 4032 3978 4050
rect 3960 4050 3978 4068
rect 3960 4068 3978 4086
rect 3960 4086 3978 4104
rect 3960 4104 3978 4122
rect 3960 4122 3978 4140
rect 3960 4140 3978 4158
rect 3960 4158 3978 4176
rect 3960 4176 3978 4194
rect 3960 4194 3978 4212
rect 3960 4212 3978 4230
rect 3960 4230 3978 4248
rect 3960 4248 3978 4266
rect 3960 4266 3978 4284
rect 3960 4284 3978 4302
rect 3960 4302 3978 4320
rect 3960 4320 3978 4338
rect 3960 4338 3978 4356
rect 3960 4356 3978 4374
rect 3960 4374 3978 4392
rect 3960 4392 3978 4410
rect 3960 4410 3978 4428
rect 3960 4428 3978 4446
rect 3960 4446 3978 4464
rect 3960 4464 3978 4482
rect 3960 4482 3978 4500
rect 3960 4500 3978 4518
rect 3960 4518 3978 4536
rect 3960 4536 3978 4554
rect 3960 4554 3978 4572
rect 3960 4572 3978 4590
rect 3960 4590 3978 4608
rect 3960 4608 3978 4626
rect 3960 4626 3978 4644
rect 3960 4644 3978 4662
rect 3960 4662 3978 4680
rect 3960 4680 3978 4698
rect 3960 4698 3978 4716
rect 3960 4716 3978 4734
rect 3960 4734 3978 4752
rect 3960 4752 3978 4770
rect 3960 4770 3978 4788
rect 3960 4788 3978 4806
rect 3960 4806 3978 4824
rect 3960 4824 3978 4842
rect 3960 4842 3978 4860
rect 3960 4860 3978 4878
rect 3960 4878 3978 4896
rect 3960 4896 3978 4914
rect 3960 4914 3978 4932
rect 3960 4932 3978 4950
rect 3960 4950 3978 4968
rect 3960 4968 3978 4986
rect 3960 4986 3978 5004
rect 3960 5004 3978 5022
rect 3960 5022 3978 5040
rect 3960 5040 3978 5058
rect 3960 5058 3978 5076
rect 3960 5076 3978 5094
rect 3960 5094 3978 5112
rect 3960 5112 3978 5130
rect 3960 5130 3978 5148
rect 3960 5148 3978 5166
rect 3960 5166 3978 5184
rect 3960 5184 3978 5202
rect 3960 5202 3978 5220
rect 3960 5220 3978 5238
rect 3960 5238 3978 5256
rect 3960 5256 3978 5274
rect 3960 5274 3978 5292
rect 3960 5292 3978 5310
rect 3960 5310 3978 5328
rect 3960 5328 3978 5346
rect 3960 5346 3978 5364
rect 3960 5364 3978 5382
rect 3960 5382 3978 5400
rect 3960 5400 3978 5418
rect 3960 5418 3978 5436
rect 3960 5436 3978 5454
rect 3960 5454 3978 5472
rect 3960 5472 3978 5490
rect 3960 5490 3978 5508
rect 3960 5508 3978 5526
rect 3960 5526 3978 5544
rect 3960 5544 3978 5562
rect 3960 5562 3978 5580
rect 3960 5580 3978 5598
rect 3960 5598 3978 5616
rect 3960 5616 3978 5634
rect 3960 5634 3978 5652
rect 3960 5652 3978 5670
rect 3960 5670 3978 5688
rect 3960 5688 3978 5706
rect 3960 5706 3978 5724
rect 3960 5724 3978 5742
rect 3960 5742 3978 5760
rect 3960 5760 3978 5778
rect 3960 5778 3978 5796
rect 3960 5796 3978 5814
rect 3960 5814 3978 5832
rect 3960 5832 3978 5850
rect 3960 5850 3978 5868
rect 3960 5868 3978 5886
rect 3960 5886 3978 5904
rect 3960 5904 3978 5922
rect 3960 5922 3978 5940
rect 3960 5940 3978 5958
rect 3960 5958 3978 5976
rect 3960 5976 3978 5994
rect 3960 5994 3978 6012
rect 3960 6642 3978 6660
rect 3960 6660 3978 6678
rect 3960 6678 3978 6696
rect 3960 6696 3978 6714
rect 3960 6714 3978 6732
rect 3960 6732 3978 6750
rect 3960 6750 3978 6768
rect 3960 6768 3978 6786
rect 3960 6786 3978 6804
rect 3960 6804 3978 6822
rect 3960 6822 3978 6840
rect 3960 6840 3978 6858
rect 3960 6858 3978 6876
rect 3960 6876 3978 6894
rect 3960 6894 3978 6912
rect 3960 6912 3978 6930
rect 3960 6930 3978 6948
rect 3960 6948 3978 6966
rect 3960 6966 3978 6984
rect 3960 6984 3978 7002
rect 3960 7002 3978 7020
rect 3960 7020 3978 7038
rect 3960 7038 3978 7056
rect 3960 7056 3978 7074
rect 3960 7074 3978 7092
rect 3960 7092 3978 7110
rect 3960 7110 3978 7128
rect 3960 7128 3978 7146
rect 3960 7146 3978 7164
rect 3960 7164 3978 7182
rect 3960 7182 3978 7200
rect 3960 7200 3978 7218
rect 3960 7218 3978 7236
rect 3960 7236 3978 7254
rect 3978 18 3996 36
rect 3978 36 3996 54
rect 3978 54 3996 72
rect 3978 72 3996 90
rect 3978 90 3996 108
rect 3978 108 3996 126
rect 3978 126 3996 144
rect 3978 144 3996 162
rect 3978 162 3996 180
rect 3978 180 3996 198
rect 3978 198 3996 216
rect 3978 216 3996 234
rect 3978 234 3996 252
rect 3978 252 3996 270
rect 3978 270 3996 288
rect 3978 288 3996 306
rect 3978 306 3996 324
rect 3978 324 3996 342
rect 3978 342 3996 360
rect 3978 360 3996 378
rect 3978 378 3996 396
rect 3978 396 3996 414
rect 3978 414 3996 432
rect 3978 432 3996 450
rect 3978 450 3996 468
rect 3978 468 3996 486
rect 3978 486 3996 504
rect 3978 504 3996 522
rect 3978 522 3996 540
rect 3978 540 3996 558
rect 3978 558 3996 576
rect 3978 576 3996 594
rect 3978 594 3996 612
rect 3978 612 3996 630
rect 3978 630 3996 648
rect 3978 864 3996 882
rect 3978 882 3996 900
rect 3978 900 3996 918
rect 3978 918 3996 936
rect 3978 936 3996 954
rect 3978 954 3996 972
rect 3978 972 3996 990
rect 3978 990 3996 1008
rect 3978 1008 3996 1026
rect 3978 1026 3996 1044
rect 3978 1044 3996 1062
rect 3978 1062 3996 1080
rect 3978 1080 3996 1098
rect 3978 1098 3996 1116
rect 3978 1116 3996 1134
rect 3978 1134 3996 1152
rect 3978 1152 3996 1170
rect 3978 1170 3996 1188
rect 3978 1188 3996 1206
rect 3978 1206 3996 1224
rect 3978 1224 3996 1242
rect 3978 1242 3996 1260
rect 3978 1260 3996 1278
rect 3978 1278 3996 1296
rect 3978 1296 3996 1314
rect 3978 1314 3996 1332
rect 3978 1332 3996 1350
rect 3978 1350 3996 1368
rect 3978 1368 3996 1386
rect 3978 1386 3996 1404
rect 3978 1404 3996 1422
rect 3978 1422 3996 1440
rect 3978 1440 3996 1458
rect 3978 1458 3996 1476
rect 3978 1476 3996 1494
rect 3978 1494 3996 1512
rect 3978 1512 3996 1530
rect 3978 1530 3996 1548
rect 3978 1782 3996 1800
rect 3978 1800 3996 1818
rect 3978 1818 3996 1836
rect 3978 1836 3996 1854
rect 3978 1854 3996 1872
rect 3978 1872 3996 1890
rect 3978 1890 3996 1908
rect 3978 1908 3996 1926
rect 3978 1926 3996 1944
rect 3978 1944 3996 1962
rect 3978 1962 3996 1980
rect 3978 1980 3996 1998
rect 3978 1998 3996 2016
rect 3978 2016 3996 2034
rect 3978 2034 3996 2052
rect 3978 2052 3996 2070
rect 3978 2070 3996 2088
rect 3978 2088 3996 2106
rect 3978 2106 3996 2124
rect 3978 2124 3996 2142
rect 3978 2142 3996 2160
rect 3978 2160 3996 2178
rect 3978 2178 3996 2196
rect 3978 2196 3996 2214
rect 3978 2214 3996 2232
rect 3978 2232 3996 2250
rect 3978 2250 3996 2268
rect 3978 2268 3996 2286
rect 3978 2286 3996 2304
rect 3978 2304 3996 2322
rect 3978 2322 3996 2340
rect 3978 2340 3996 2358
rect 3978 2358 3996 2376
rect 3978 2376 3996 2394
rect 3978 2394 3996 2412
rect 3978 2412 3996 2430
rect 3978 2430 3996 2448
rect 3978 2448 3996 2466
rect 3978 2466 3996 2484
rect 3978 2484 3996 2502
rect 3978 2502 3996 2520
rect 3978 2520 3996 2538
rect 3978 2538 3996 2556
rect 3978 2556 3996 2574
rect 3978 2574 3996 2592
rect 3978 2592 3996 2610
rect 3978 2610 3996 2628
rect 3978 2628 3996 2646
rect 3978 2646 3996 2664
rect 3978 2664 3996 2682
rect 3978 2682 3996 2700
rect 3978 2700 3996 2718
rect 3978 2718 3996 2736
rect 3978 2736 3996 2754
rect 3978 2754 3996 2772
rect 3978 2772 3996 2790
rect 3978 2790 3996 2808
rect 3978 2808 3996 2826
rect 3978 2826 3996 2844
rect 3978 2844 3996 2862
rect 3978 2862 3996 2880
rect 3978 2880 3996 2898
rect 3978 2898 3996 2916
rect 3978 2916 3996 2934
rect 3978 2934 3996 2952
rect 3978 2952 3996 2970
rect 3978 2970 3996 2988
rect 3978 2988 3996 3006
rect 3978 3006 3996 3024
rect 3978 3024 3996 3042
rect 3978 3042 3996 3060
rect 3978 3294 3996 3312
rect 3978 3312 3996 3330
rect 3978 3330 3996 3348
rect 3978 3348 3996 3366
rect 3978 3366 3996 3384
rect 3978 3384 3996 3402
rect 3978 3402 3996 3420
rect 3978 3420 3996 3438
rect 3978 3438 3996 3456
rect 3978 3456 3996 3474
rect 3978 3474 3996 3492
rect 3978 3492 3996 3510
rect 3978 3510 3996 3528
rect 3978 3528 3996 3546
rect 3978 3546 3996 3564
rect 3978 3564 3996 3582
rect 3978 3582 3996 3600
rect 3978 3600 3996 3618
rect 3978 3618 3996 3636
rect 3978 3636 3996 3654
rect 3978 3654 3996 3672
rect 3978 3672 3996 3690
rect 3978 3690 3996 3708
rect 3978 3708 3996 3726
rect 3978 3726 3996 3744
rect 3978 3744 3996 3762
rect 3978 3762 3996 3780
rect 3978 3780 3996 3798
rect 3978 3798 3996 3816
rect 3978 3816 3996 3834
rect 3978 3834 3996 3852
rect 3978 3852 3996 3870
rect 3978 3870 3996 3888
rect 3978 3888 3996 3906
rect 3978 3906 3996 3924
rect 3978 3924 3996 3942
rect 3978 3942 3996 3960
rect 3978 3960 3996 3978
rect 3978 3978 3996 3996
rect 3978 3996 3996 4014
rect 3978 4014 3996 4032
rect 3978 4032 3996 4050
rect 3978 4050 3996 4068
rect 3978 4068 3996 4086
rect 3978 4086 3996 4104
rect 3978 4104 3996 4122
rect 3978 4122 3996 4140
rect 3978 4140 3996 4158
rect 3978 4158 3996 4176
rect 3978 4176 3996 4194
rect 3978 4194 3996 4212
rect 3978 4212 3996 4230
rect 3978 4230 3996 4248
rect 3978 4248 3996 4266
rect 3978 4266 3996 4284
rect 3978 4284 3996 4302
rect 3978 4302 3996 4320
rect 3978 4320 3996 4338
rect 3978 4338 3996 4356
rect 3978 4356 3996 4374
rect 3978 4374 3996 4392
rect 3978 4392 3996 4410
rect 3978 4410 3996 4428
rect 3978 4428 3996 4446
rect 3978 4446 3996 4464
rect 3978 4464 3996 4482
rect 3978 4482 3996 4500
rect 3978 4500 3996 4518
rect 3978 4518 3996 4536
rect 3978 4536 3996 4554
rect 3978 4554 3996 4572
rect 3978 4572 3996 4590
rect 3978 4590 3996 4608
rect 3978 4608 3996 4626
rect 3978 4626 3996 4644
rect 3978 4644 3996 4662
rect 3978 4662 3996 4680
rect 3978 4680 3996 4698
rect 3978 4698 3996 4716
rect 3978 4716 3996 4734
rect 3978 4734 3996 4752
rect 3978 4752 3996 4770
rect 3978 4770 3996 4788
rect 3978 4788 3996 4806
rect 3978 4806 3996 4824
rect 3978 4824 3996 4842
rect 3978 4842 3996 4860
rect 3978 4860 3996 4878
rect 3978 4878 3996 4896
rect 3978 4896 3996 4914
rect 3978 4914 3996 4932
rect 3978 4932 3996 4950
rect 3978 4950 3996 4968
rect 3978 4968 3996 4986
rect 3978 4986 3996 5004
rect 3978 5004 3996 5022
rect 3978 5022 3996 5040
rect 3978 5040 3996 5058
rect 3978 5058 3996 5076
rect 3978 5076 3996 5094
rect 3978 5094 3996 5112
rect 3978 5112 3996 5130
rect 3978 5130 3996 5148
rect 3978 5148 3996 5166
rect 3978 5166 3996 5184
rect 3978 5184 3996 5202
rect 3978 5202 3996 5220
rect 3978 5220 3996 5238
rect 3978 5238 3996 5256
rect 3978 5256 3996 5274
rect 3978 5274 3996 5292
rect 3978 5292 3996 5310
rect 3978 5310 3996 5328
rect 3978 5328 3996 5346
rect 3978 5346 3996 5364
rect 3978 5364 3996 5382
rect 3978 5382 3996 5400
rect 3978 5400 3996 5418
rect 3978 5418 3996 5436
rect 3978 5436 3996 5454
rect 3978 5454 3996 5472
rect 3978 5472 3996 5490
rect 3978 5490 3996 5508
rect 3978 5508 3996 5526
rect 3978 5526 3996 5544
rect 3978 5544 3996 5562
rect 3978 5562 3996 5580
rect 3978 5580 3996 5598
rect 3978 5598 3996 5616
rect 3978 5616 3996 5634
rect 3978 5634 3996 5652
rect 3978 5652 3996 5670
rect 3978 5670 3996 5688
rect 3978 5688 3996 5706
rect 3978 5706 3996 5724
rect 3978 5724 3996 5742
rect 3978 5742 3996 5760
rect 3978 5760 3996 5778
rect 3978 5778 3996 5796
rect 3978 5796 3996 5814
rect 3978 5814 3996 5832
rect 3978 5832 3996 5850
rect 3978 5850 3996 5868
rect 3978 5868 3996 5886
rect 3978 5886 3996 5904
rect 3978 5904 3996 5922
rect 3978 5922 3996 5940
rect 3978 5940 3996 5958
rect 3978 5958 3996 5976
rect 3978 5976 3996 5994
rect 3978 5994 3996 6012
rect 3978 6012 3996 6030
rect 3978 6030 3996 6048
rect 3978 6624 3996 6642
rect 3978 6642 3996 6660
rect 3978 6660 3996 6678
rect 3978 6678 3996 6696
rect 3978 6696 3996 6714
rect 3978 6714 3996 6732
rect 3978 6732 3996 6750
rect 3978 6750 3996 6768
rect 3978 6768 3996 6786
rect 3978 6786 3996 6804
rect 3978 6804 3996 6822
rect 3978 6822 3996 6840
rect 3978 6840 3996 6858
rect 3978 6858 3996 6876
rect 3978 6876 3996 6894
rect 3978 6894 3996 6912
rect 3978 6912 3996 6930
rect 3978 6930 3996 6948
rect 3978 6948 3996 6966
rect 3978 6966 3996 6984
rect 3978 6984 3996 7002
rect 3978 7002 3996 7020
rect 3978 7020 3996 7038
rect 3978 7038 3996 7056
rect 3978 7056 3996 7074
rect 3978 7074 3996 7092
rect 3978 7092 3996 7110
rect 3978 7110 3996 7128
rect 3978 7128 3996 7146
rect 3978 7146 3996 7164
rect 3978 7164 3996 7182
rect 3978 7182 3996 7200
rect 3978 7200 3996 7218
rect 3978 7218 3996 7236
rect 3978 7236 3996 7254
rect 3996 18 4014 36
rect 3996 36 4014 54
rect 3996 54 4014 72
rect 3996 72 4014 90
rect 3996 90 4014 108
rect 3996 108 4014 126
rect 3996 126 4014 144
rect 3996 144 4014 162
rect 3996 162 4014 180
rect 3996 180 4014 198
rect 3996 198 4014 216
rect 3996 216 4014 234
rect 3996 234 4014 252
rect 3996 252 4014 270
rect 3996 270 4014 288
rect 3996 288 4014 306
rect 3996 306 4014 324
rect 3996 324 4014 342
rect 3996 342 4014 360
rect 3996 360 4014 378
rect 3996 378 4014 396
rect 3996 396 4014 414
rect 3996 414 4014 432
rect 3996 432 4014 450
rect 3996 450 4014 468
rect 3996 468 4014 486
rect 3996 486 4014 504
rect 3996 504 4014 522
rect 3996 522 4014 540
rect 3996 540 4014 558
rect 3996 558 4014 576
rect 3996 576 4014 594
rect 3996 594 4014 612
rect 3996 612 4014 630
rect 3996 630 4014 648
rect 3996 864 4014 882
rect 3996 882 4014 900
rect 3996 900 4014 918
rect 3996 918 4014 936
rect 3996 936 4014 954
rect 3996 954 4014 972
rect 3996 972 4014 990
rect 3996 990 4014 1008
rect 3996 1008 4014 1026
rect 3996 1026 4014 1044
rect 3996 1044 4014 1062
rect 3996 1062 4014 1080
rect 3996 1080 4014 1098
rect 3996 1098 4014 1116
rect 3996 1116 4014 1134
rect 3996 1134 4014 1152
rect 3996 1152 4014 1170
rect 3996 1170 4014 1188
rect 3996 1188 4014 1206
rect 3996 1206 4014 1224
rect 3996 1224 4014 1242
rect 3996 1242 4014 1260
rect 3996 1260 4014 1278
rect 3996 1278 4014 1296
rect 3996 1296 4014 1314
rect 3996 1314 4014 1332
rect 3996 1332 4014 1350
rect 3996 1350 4014 1368
rect 3996 1368 4014 1386
rect 3996 1386 4014 1404
rect 3996 1404 4014 1422
rect 3996 1422 4014 1440
rect 3996 1440 4014 1458
rect 3996 1458 4014 1476
rect 3996 1476 4014 1494
rect 3996 1494 4014 1512
rect 3996 1512 4014 1530
rect 3996 1530 4014 1548
rect 3996 1548 4014 1566
rect 3996 1800 4014 1818
rect 3996 1818 4014 1836
rect 3996 1836 4014 1854
rect 3996 1854 4014 1872
rect 3996 1872 4014 1890
rect 3996 1890 4014 1908
rect 3996 1908 4014 1926
rect 3996 1926 4014 1944
rect 3996 1944 4014 1962
rect 3996 1962 4014 1980
rect 3996 1980 4014 1998
rect 3996 1998 4014 2016
rect 3996 2016 4014 2034
rect 3996 2034 4014 2052
rect 3996 2052 4014 2070
rect 3996 2070 4014 2088
rect 3996 2088 4014 2106
rect 3996 2106 4014 2124
rect 3996 2124 4014 2142
rect 3996 2142 4014 2160
rect 3996 2160 4014 2178
rect 3996 2178 4014 2196
rect 3996 2196 4014 2214
rect 3996 2214 4014 2232
rect 3996 2232 4014 2250
rect 3996 2250 4014 2268
rect 3996 2268 4014 2286
rect 3996 2286 4014 2304
rect 3996 2304 4014 2322
rect 3996 2322 4014 2340
rect 3996 2340 4014 2358
rect 3996 2358 4014 2376
rect 3996 2376 4014 2394
rect 3996 2394 4014 2412
rect 3996 2412 4014 2430
rect 3996 2430 4014 2448
rect 3996 2448 4014 2466
rect 3996 2466 4014 2484
rect 3996 2484 4014 2502
rect 3996 2502 4014 2520
rect 3996 2520 4014 2538
rect 3996 2538 4014 2556
rect 3996 2556 4014 2574
rect 3996 2574 4014 2592
rect 3996 2592 4014 2610
rect 3996 2610 4014 2628
rect 3996 2628 4014 2646
rect 3996 2646 4014 2664
rect 3996 2664 4014 2682
rect 3996 2682 4014 2700
rect 3996 2700 4014 2718
rect 3996 2718 4014 2736
rect 3996 2736 4014 2754
rect 3996 2754 4014 2772
rect 3996 2772 4014 2790
rect 3996 2790 4014 2808
rect 3996 2808 4014 2826
rect 3996 2826 4014 2844
rect 3996 2844 4014 2862
rect 3996 2862 4014 2880
rect 3996 2880 4014 2898
rect 3996 2898 4014 2916
rect 3996 2916 4014 2934
rect 3996 2934 4014 2952
rect 3996 2952 4014 2970
rect 3996 2970 4014 2988
rect 3996 2988 4014 3006
rect 3996 3006 4014 3024
rect 3996 3024 4014 3042
rect 3996 3042 4014 3060
rect 3996 3060 4014 3078
rect 3996 3078 4014 3096
rect 3996 3312 4014 3330
rect 3996 3330 4014 3348
rect 3996 3348 4014 3366
rect 3996 3366 4014 3384
rect 3996 3384 4014 3402
rect 3996 3402 4014 3420
rect 3996 3420 4014 3438
rect 3996 3438 4014 3456
rect 3996 3456 4014 3474
rect 3996 3474 4014 3492
rect 3996 3492 4014 3510
rect 3996 3510 4014 3528
rect 3996 3528 4014 3546
rect 3996 3546 4014 3564
rect 3996 3564 4014 3582
rect 3996 3582 4014 3600
rect 3996 3600 4014 3618
rect 3996 3618 4014 3636
rect 3996 3636 4014 3654
rect 3996 3654 4014 3672
rect 3996 3672 4014 3690
rect 3996 3690 4014 3708
rect 3996 3708 4014 3726
rect 3996 3726 4014 3744
rect 3996 3744 4014 3762
rect 3996 3762 4014 3780
rect 3996 3780 4014 3798
rect 3996 3798 4014 3816
rect 3996 3816 4014 3834
rect 3996 3834 4014 3852
rect 3996 3852 4014 3870
rect 3996 3870 4014 3888
rect 3996 3888 4014 3906
rect 3996 3906 4014 3924
rect 3996 3924 4014 3942
rect 3996 3942 4014 3960
rect 3996 3960 4014 3978
rect 3996 3978 4014 3996
rect 3996 3996 4014 4014
rect 3996 4014 4014 4032
rect 3996 4032 4014 4050
rect 3996 4050 4014 4068
rect 3996 4068 4014 4086
rect 3996 4086 4014 4104
rect 3996 4104 4014 4122
rect 3996 4122 4014 4140
rect 3996 4140 4014 4158
rect 3996 4158 4014 4176
rect 3996 4176 4014 4194
rect 3996 4194 4014 4212
rect 3996 4212 4014 4230
rect 3996 4230 4014 4248
rect 3996 4248 4014 4266
rect 3996 4266 4014 4284
rect 3996 4284 4014 4302
rect 3996 4302 4014 4320
rect 3996 4320 4014 4338
rect 3996 4338 4014 4356
rect 3996 4356 4014 4374
rect 3996 4374 4014 4392
rect 3996 4392 4014 4410
rect 3996 4410 4014 4428
rect 3996 4428 4014 4446
rect 3996 4446 4014 4464
rect 3996 4464 4014 4482
rect 3996 4482 4014 4500
rect 3996 4500 4014 4518
rect 3996 4518 4014 4536
rect 3996 4536 4014 4554
rect 3996 4554 4014 4572
rect 3996 4572 4014 4590
rect 3996 4590 4014 4608
rect 3996 4608 4014 4626
rect 3996 4626 4014 4644
rect 3996 4644 4014 4662
rect 3996 4662 4014 4680
rect 3996 4680 4014 4698
rect 3996 4698 4014 4716
rect 3996 4716 4014 4734
rect 3996 4734 4014 4752
rect 3996 4752 4014 4770
rect 3996 4770 4014 4788
rect 3996 4788 4014 4806
rect 3996 4806 4014 4824
rect 3996 4824 4014 4842
rect 3996 4842 4014 4860
rect 3996 4860 4014 4878
rect 3996 4878 4014 4896
rect 3996 4896 4014 4914
rect 3996 4914 4014 4932
rect 3996 4932 4014 4950
rect 3996 4950 4014 4968
rect 3996 4968 4014 4986
rect 3996 4986 4014 5004
rect 3996 5004 4014 5022
rect 3996 5022 4014 5040
rect 3996 5040 4014 5058
rect 3996 5058 4014 5076
rect 3996 5076 4014 5094
rect 3996 5094 4014 5112
rect 3996 5112 4014 5130
rect 3996 5130 4014 5148
rect 3996 5148 4014 5166
rect 3996 5166 4014 5184
rect 3996 5184 4014 5202
rect 3996 5202 4014 5220
rect 3996 5220 4014 5238
rect 3996 5238 4014 5256
rect 3996 5256 4014 5274
rect 3996 5274 4014 5292
rect 3996 5292 4014 5310
rect 3996 5310 4014 5328
rect 3996 5328 4014 5346
rect 3996 5346 4014 5364
rect 3996 5364 4014 5382
rect 3996 5382 4014 5400
rect 3996 5400 4014 5418
rect 3996 5418 4014 5436
rect 3996 5436 4014 5454
rect 3996 5454 4014 5472
rect 3996 5472 4014 5490
rect 3996 5490 4014 5508
rect 3996 5508 4014 5526
rect 3996 5526 4014 5544
rect 3996 5544 4014 5562
rect 3996 5562 4014 5580
rect 3996 5580 4014 5598
rect 3996 5598 4014 5616
rect 3996 5616 4014 5634
rect 3996 5634 4014 5652
rect 3996 5652 4014 5670
rect 3996 5670 4014 5688
rect 3996 5688 4014 5706
rect 3996 5706 4014 5724
rect 3996 5724 4014 5742
rect 3996 5742 4014 5760
rect 3996 5760 4014 5778
rect 3996 5778 4014 5796
rect 3996 5796 4014 5814
rect 3996 5814 4014 5832
rect 3996 5832 4014 5850
rect 3996 5850 4014 5868
rect 3996 5868 4014 5886
rect 3996 5886 4014 5904
rect 3996 5904 4014 5922
rect 3996 5922 4014 5940
rect 3996 5940 4014 5958
rect 3996 5958 4014 5976
rect 3996 5976 4014 5994
rect 3996 5994 4014 6012
rect 3996 6012 4014 6030
rect 3996 6030 4014 6048
rect 3996 6048 4014 6066
rect 3996 6066 4014 6084
rect 3996 6624 4014 6642
rect 3996 6642 4014 6660
rect 3996 6660 4014 6678
rect 3996 6678 4014 6696
rect 3996 6696 4014 6714
rect 3996 6714 4014 6732
rect 3996 6732 4014 6750
rect 3996 6750 4014 6768
rect 3996 6768 4014 6786
rect 3996 6786 4014 6804
rect 3996 6804 4014 6822
rect 3996 6822 4014 6840
rect 3996 6840 4014 6858
rect 3996 6858 4014 6876
rect 3996 6876 4014 6894
rect 3996 6894 4014 6912
rect 3996 6912 4014 6930
rect 3996 6930 4014 6948
rect 3996 6948 4014 6966
rect 3996 6966 4014 6984
rect 3996 6984 4014 7002
rect 3996 7002 4014 7020
rect 3996 7020 4014 7038
rect 3996 7038 4014 7056
rect 3996 7056 4014 7074
rect 3996 7074 4014 7092
rect 3996 7092 4014 7110
rect 3996 7110 4014 7128
rect 3996 7128 4014 7146
rect 3996 7146 4014 7164
rect 3996 7164 4014 7182
rect 3996 7182 4014 7200
rect 3996 7200 4014 7218
rect 3996 7218 4014 7236
rect 3996 7236 4014 7254
rect 4014 18 4032 36
rect 4014 36 4032 54
rect 4014 54 4032 72
rect 4014 72 4032 90
rect 4014 90 4032 108
rect 4014 108 4032 126
rect 4014 126 4032 144
rect 4014 144 4032 162
rect 4014 162 4032 180
rect 4014 180 4032 198
rect 4014 198 4032 216
rect 4014 216 4032 234
rect 4014 234 4032 252
rect 4014 252 4032 270
rect 4014 270 4032 288
rect 4014 288 4032 306
rect 4014 306 4032 324
rect 4014 324 4032 342
rect 4014 342 4032 360
rect 4014 360 4032 378
rect 4014 378 4032 396
rect 4014 396 4032 414
rect 4014 414 4032 432
rect 4014 432 4032 450
rect 4014 450 4032 468
rect 4014 468 4032 486
rect 4014 486 4032 504
rect 4014 504 4032 522
rect 4014 522 4032 540
rect 4014 540 4032 558
rect 4014 558 4032 576
rect 4014 576 4032 594
rect 4014 594 4032 612
rect 4014 612 4032 630
rect 4014 630 4032 648
rect 4014 864 4032 882
rect 4014 882 4032 900
rect 4014 900 4032 918
rect 4014 918 4032 936
rect 4014 936 4032 954
rect 4014 954 4032 972
rect 4014 972 4032 990
rect 4014 990 4032 1008
rect 4014 1008 4032 1026
rect 4014 1026 4032 1044
rect 4014 1044 4032 1062
rect 4014 1062 4032 1080
rect 4014 1080 4032 1098
rect 4014 1098 4032 1116
rect 4014 1116 4032 1134
rect 4014 1134 4032 1152
rect 4014 1152 4032 1170
rect 4014 1170 4032 1188
rect 4014 1188 4032 1206
rect 4014 1206 4032 1224
rect 4014 1224 4032 1242
rect 4014 1242 4032 1260
rect 4014 1260 4032 1278
rect 4014 1278 4032 1296
rect 4014 1296 4032 1314
rect 4014 1314 4032 1332
rect 4014 1332 4032 1350
rect 4014 1350 4032 1368
rect 4014 1368 4032 1386
rect 4014 1386 4032 1404
rect 4014 1404 4032 1422
rect 4014 1422 4032 1440
rect 4014 1440 4032 1458
rect 4014 1458 4032 1476
rect 4014 1476 4032 1494
rect 4014 1494 4032 1512
rect 4014 1512 4032 1530
rect 4014 1530 4032 1548
rect 4014 1548 4032 1566
rect 4014 1566 4032 1584
rect 4014 1818 4032 1836
rect 4014 1836 4032 1854
rect 4014 1854 4032 1872
rect 4014 1872 4032 1890
rect 4014 1890 4032 1908
rect 4014 1908 4032 1926
rect 4014 1926 4032 1944
rect 4014 1944 4032 1962
rect 4014 1962 4032 1980
rect 4014 1980 4032 1998
rect 4014 1998 4032 2016
rect 4014 2016 4032 2034
rect 4014 2034 4032 2052
rect 4014 2052 4032 2070
rect 4014 2070 4032 2088
rect 4014 2088 4032 2106
rect 4014 2106 4032 2124
rect 4014 2124 4032 2142
rect 4014 2142 4032 2160
rect 4014 2160 4032 2178
rect 4014 2178 4032 2196
rect 4014 2196 4032 2214
rect 4014 2214 4032 2232
rect 4014 2232 4032 2250
rect 4014 2250 4032 2268
rect 4014 2268 4032 2286
rect 4014 2286 4032 2304
rect 4014 2304 4032 2322
rect 4014 2322 4032 2340
rect 4014 2340 4032 2358
rect 4014 2358 4032 2376
rect 4014 2376 4032 2394
rect 4014 2394 4032 2412
rect 4014 2412 4032 2430
rect 4014 2430 4032 2448
rect 4014 2448 4032 2466
rect 4014 2466 4032 2484
rect 4014 2484 4032 2502
rect 4014 2502 4032 2520
rect 4014 2520 4032 2538
rect 4014 2538 4032 2556
rect 4014 2556 4032 2574
rect 4014 2574 4032 2592
rect 4014 2592 4032 2610
rect 4014 2610 4032 2628
rect 4014 2628 4032 2646
rect 4014 2646 4032 2664
rect 4014 2664 4032 2682
rect 4014 2682 4032 2700
rect 4014 2700 4032 2718
rect 4014 2718 4032 2736
rect 4014 2736 4032 2754
rect 4014 2754 4032 2772
rect 4014 2772 4032 2790
rect 4014 2790 4032 2808
rect 4014 2808 4032 2826
rect 4014 2826 4032 2844
rect 4014 2844 4032 2862
rect 4014 2862 4032 2880
rect 4014 2880 4032 2898
rect 4014 2898 4032 2916
rect 4014 2916 4032 2934
rect 4014 2934 4032 2952
rect 4014 2952 4032 2970
rect 4014 2970 4032 2988
rect 4014 2988 4032 3006
rect 4014 3006 4032 3024
rect 4014 3024 4032 3042
rect 4014 3042 4032 3060
rect 4014 3060 4032 3078
rect 4014 3078 4032 3096
rect 4014 3096 4032 3114
rect 4014 3348 4032 3366
rect 4014 3366 4032 3384
rect 4014 3384 4032 3402
rect 4014 3402 4032 3420
rect 4014 3420 4032 3438
rect 4014 3438 4032 3456
rect 4014 3456 4032 3474
rect 4014 3474 4032 3492
rect 4014 3492 4032 3510
rect 4014 3510 4032 3528
rect 4014 3528 4032 3546
rect 4014 3546 4032 3564
rect 4014 3564 4032 3582
rect 4014 3582 4032 3600
rect 4014 3600 4032 3618
rect 4014 3618 4032 3636
rect 4014 3636 4032 3654
rect 4014 3654 4032 3672
rect 4014 3672 4032 3690
rect 4014 3690 4032 3708
rect 4014 3708 4032 3726
rect 4014 3726 4032 3744
rect 4014 3744 4032 3762
rect 4014 3762 4032 3780
rect 4014 3780 4032 3798
rect 4014 3798 4032 3816
rect 4014 3816 4032 3834
rect 4014 3834 4032 3852
rect 4014 3852 4032 3870
rect 4014 3870 4032 3888
rect 4014 3888 4032 3906
rect 4014 3906 4032 3924
rect 4014 3924 4032 3942
rect 4014 3942 4032 3960
rect 4014 3960 4032 3978
rect 4014 3978 4032 3996
rect 4014 3996 4032 4014
rect 4014 4014 4032 4032
rect 4014 4032 4032 4050
rect 4014 4050 4032 4068
rect 4014 4068 4032 4086
rect 4014 4086 4032 4104
rect 4014 4104 4032 4122
rect 4014 4122 4032 4140
rect 4014 4140 4032 4158
rect 4014 4158 4032 4176
rect 4014 4176 4032 4194
rect 4014 4194 4032 4212
rect 4014 4212 4032 4230
rect 4014 4230 4032 4248
rect 4014 4248 4032 4266
rect 4014 4266 4032 4284
rect 4014 4284 4032 4302
rect 4014 4302 4032 4320
rect 4014 4320 4032 4338
rect 4014 4338 4032 4356
rect 4014 4356 4032 4374
rect 4014 4374 4032 4392
rect 4014 4392 4032 4410
rect 4014 4410 4032 4428
rect 4014 4428 4032 4446
rect 4014 4446 4032 4464
rect 4014 4464 4032 4482
rect 4014 4482 4032 4500
rect 4014 4500 4032 4518
rect 4014 4518 4032 4536
rect 4014 4536 4032 4554
rect 4014 4554 4032 4572
rect 4014 4572 4032 4590
rect 4014 4590 4032 4608
rect 4014 4608 4032 4626
rect 4014 4626 4032 4644
rect 4014 4644 4032 4662
rect 4014 4662 4032 4680
rect 4014 4680 4032 4698
rect 4014 4698 4032 4716
rect 4014 4716 4032 4734
rect 4014 4734 4032 4752
rect 4014 4752 4032 4770
rect 4014 4770 4032 4788
rect 4014 4788 4032 4806
rect 4014 4806 4032 4824
rect 4014 4824 4032 4842
rect 4014 4842 4032 4860
rect 4014 4860 4032 4878
rect 4014 4878 4032 4896
rect 4014 4896 4032 4914
rect 4014 4914 4032 4932
rect 4014 4932 4032 4950
rect 4014 4950 4032 4968
rect 4014 4968 4032 4986
rect 4014 4986 4032 5004
rect 4014 5004 4032 5022
rect 4014 5022 4032 5040
rect 4014 5040 4032 5058
rect 4014 5058 4032 5076
rect 4014 5076 4032 5094
rect 4014 5094 4032 5112
rect 4014 5112 4032 5130
rect 4014 5130 4032 5148
rect 4014 5148 4032 5166
rect 4014 5166 4032 5184
rect 4014 5184 4032 5202
rect 4014 5202 4032 5220
rect 4014 5220 4032 5238
rect 4014 5238 4032 5256
rect 4014 5256 4032 5274
rect 4014 5274 4032 5292
rect 4014 5292 4032 5310
rect 4014 5310 4032 5328
rect 4014 5328 4032 5346
rect 4014 5346 4032 5364
rect 4014 5364 4032 5382
rect 4014 5382 4032 5400
rect 4014 5400 4032 5418
rect 4014 5418 4032 5436
rect 4014 5436 4032 5454
rect 4014 5454 4032 5472
rect 4014 5472 4032 5490
rect 4014 5490 4032 5508
rect 4014 5508 4032 5526
rect 4014 5526 4032 5544
rect 4014 5544 4032 5562
rect 4014 5562 4032 5580
rect 4014 5580 4032 5598
rect 4014 5598 4032 5616
rect 4014 5616 4032 5634
rect 4014 5634 4032 5652
rect 4014 5652 4032 5670
rect 4014 5670 4032 5688
rect 4014 5688 4032 5706
rect 4014 5706 4032 5724
rect 4014 5724 4032 5742
rect 4014 5742 4032 5760
rect 4014 5760 4032 5778
rect 4014 5778 4032 5796
rect 4014 5796 4032 5814
rect 4014 5814 4032 5832
rect 4014 5832 4032 5850
rect 4014 5850 4032 5868
rect 4014 5868 4032 5886
rect 4014 5886 4032 5904
rect 4014 5904 4032 5922
rect 4014 5922 4032 5940
rect 4014 5940 4032 5958
rect 4014 5958 4032 5976
rect 4014 5976 4032 5994
rect 4014 5994 4032 6012
rect 4014 6012 4032 6030
rect 4014 6030 4032 6048
rect 4014 6048 4032 6066
rect 4014 6066 4032 6084
rect 4014 6084 4032 6102
rect 4014 6102 4032 6120
rect 4014 6624 4032 6642
rect 4014 6642 4032 6660
rect 4014 6660 4032 6678
rect 4014 6678 4032 6696
rect 4014 6696 4032 6714
rect 4014 6714 4032 6732
rect 4014 6732 4032 6750
rect 4014 6750 4032 6768
rect 4014 6768 4032 6786
rect 4014 6786 4032 6804
rect 4014 6804 4032 6822
rect 4014 6822 4032 6840
rect 4014 6840 4032 6858
rect 4014 6858 4032 6876
rect 4014 6876 4032 6894
rect 4014 6894 4032 6912
rect 4014 6912 4032 6930
rect 4014 6930 4032 6948
rect 4014 6948 4032 6966
rect 4014 6966 4032 6984
rect 4014 6984 4032 7002
rect 4014 7002 4032 7020
rect 4014 7020 4032 7038
rect 4014 7038 4032 7056
rect 4014 7056 4032 7074
rect 4014 7074 4032 7092
rect 4014 7092 4032 7110
rect 4014 7110 4032 7128
rect 4014 7128 4032 7146
rect 4014 7146 4032 7164
rect 4014 7164 4032 7182
rect 4014 7182 4032 7200
rect 4014 7200 4032 7218
rect 4014 7218 4032 7236
rect 4014 7236 4032 7254
rect 4032 18 4050 36
rect 4032 36 4050 54
rect 4032 54 4050 72
rect 4032 72 4050 90
rect 4032 90 4050 108
rect 4032 108 4050 126
rect 4032 126 4050 144
rect 4032 144 4050 162
rect 4032 162 4050 180
rect 4032 180 4050 198
rect 4032 198 4050 216
rect 4032 216 4050 234
rect 4032 234 4050 252
rect 4032 252 4050 270
rect 4032 270 4050 288
rect 4032 288 4050 306
rect 4032 306 4050 324
rect 4032 324 4050 342
rect 4032 342 4050 360
rect 4032 360 4050 378
rect 4032 378 4050 396
rect 4032 396 4050 414
rect 4032 414 4050 432
rect 4032 432 4050 450
rect 4032 450 4050 468
rect 4032 468 4050 486
rect 4032 486 4050 504
rect 4032 504 4050 522
rect 4032 522 4050 540
rect 4032 540 4050 558
rect 4032 558 4050 576
rect 4032 576 4050 594
rect 4032 594 4050 612
rect 4032 612 4050 630
rect 4032 630 4050 648
rect 4032 864 4050 882
rect 4032 882 4050 900
rect 4032 900 4050 918
rect 4032 918 4050 936
rect 4032 936 4050 954
rect 4032 954 4050 972
rect 4032 972 4050 990
rect 4032 990 4050 1008
rect 4032 1008 4050 1026
rect 4032 1026 4050 1044
rect 4032 1044 4050 1062
rect 4032 1062 4050 1080
rect 4032 1080 4050 1098
rect 4032 1098 4050 1116
rect 4032 1116 4050 1134
rect 4032 1134 4050 1152
rect 4032 1152 4050 1170
rect 4032 1170 4050 1188
rect 4032 1188 4050 1206
rect 4032 1206 4050 1224
rect 4032 1224 4050 1242
rect 4032 1242 4050 1260
rect 4032 1260 4050 1278
rect 4032 1278 4050 1296
rect 4032 1296 4050 1314
rect 4032 1314 4050 1332
rect 4032 1332 4050 1350
rect 4032 1350 4050 1368
rect 4032 1368 4050 1386
rect 4032 1386 4050 1404
rect 4032 1404 4050 1422
rect 4032 1422 4050 1440
rect 4032 1440 4050 1458
rect 4032 1458 4050 1476
rect 4032 1476 4050 1494
rect 4032 1494 4050 1512
rect 4032 1512 4050 1530
rect 4032 1530 4050 1548
rect 4032 1548 4050 1566
rect 4032 1566 4050 1584
rect 4032 1818 4050 1836
rect 4032 1836 4050 1854
rect 4032 1854 4050 1872
rect 4032 1872 4050 1890
rect 4032 1890 4050 1908
rect 4032 1908 4050 1926
rect 4032 1926 4050 1944
rect 4032 1944 4050 1962
rect 4032 1962 4050 1980
rect 4032 1980 4050 1998
rect 4032 1998 4050 2016
rect 4032 2016 4050 2034
rect 4032 2034 4050 2052
rect 4032 2052 4050 2070
rect 4032 2070 4050 2088
rect 4032 2088 4050 2106
rect 4032 2106 4050 2124
rect 4032 2124 4050 2142
rect 4032 2142 4050 2160
rect 4032 2160 4050 2178
rect 4032 2178 4050 2196
rect 4032 2196 4050 2214
rect 4032 2214 4050 2232
rect 4032 2232 4050 2250
rect 4032 2250 4050 2268
rect 4032 2268 4050 2286
rect 4032 2286 4050 2304
rect 4032 2304 4050 2322
rect 4032 2322 4050 2340
rect 4032 2340 4050 2358
rect 4032 2358 4050 2376
rect 4032 2376 4050 2394
rect 4032 2394 4050 2412
rect 4032 2412 4050 2430
rect 4032 2430 4050 2448
rect 4032 2448 4050 2466
rect 4032 2466 4050 2484
rect 4032 2484 4050 2502
rect 4032 2502 4050 2520
rect 4032 2520 4050 2538
rect 4032 2538 4050 2556
rect 4032 2556 4050 2574
rect 4032 2574 4050 2592
rect 4032 2592 4050 2610
rect 4032 2610 4050 2628
rect 4032 2628 4050 2646
rect 4032 2646 4050 2664
rect 4032 2664 4050 2682
rect 4032 2682 4050 2700
rect 4032 2700 4050 2718
rect 4032 2718 4050 2736
rect 4032 2736 4050 2754
rect 4032 2754 4050 2772
rect 4032 2772 4050 2790
rect 4032 2790 4050 2808
rect 4032 2808 4050 2826
rect 4032 2826 4050 2844
rect 4032 2844 4050 2862
rect 4032 2862 4050 2880
rect 4032 2880 4050 2898
rect 4032 2898 4050 2916
rect 4032 2916 4050 2934
rect 4032 2934 4050 2952
rect 4032 2952 4050 2970
rect 4032 2970 4050 2988
rect 4032 2988 4050 3006
rect 4032 3006 4050 3024
rect 4032 3024 4050 3042
rect 4032 3042 4050 3060
rect 4032 3060 4050 3078
rect 4032 3078 4050 3096
rect 4032 3096 4050 3114
rect 4032 3114 4050 3132
rect 4032 3132 4050 3150
rect 4032 3366 4050 3384
rect 4032 3384 4050 3402
rect 4032 3402 4050 3420
rect 4032 3420 4050 3438
rect 4032 3438 4050 3456
rect 4032 3456 4050 3474
rect 4032 3474 4050 3492
rect 4032 3492 4050 3510
rect 4032 3510 4050 3528
rect 4032 3528 4050 3546
rect 4032 3546 4050 3564
rect 4032 3564 4050 3582
rect 4032 3582 4050 3600
rect 4032 3600 4050 3618
rect 4032 3618 4050 3636
rect 4032 3636 4050 3654
rect 4032 3654 4050 3672
rect 4032 3672 4050 3690
rect 4032 3690 4050 3708
rect 4032 3708 4050 3726
rect 4032 3726 4050 3744
rect 4032 3744 4050 3762
rect 4032 3762 4050 3780
rect 4032 3780 4050 3798
rect 4032 3798 4050 3816
rect 4032 3816 4050 3834
rect 4032 3834 4050 3852
rect 4032 3852 4050 3870
rect 4032 3870 4050 3888
rect 4032 3888 4050 3906
rect 4032 3906 4050 3924
rect 4032 3924 4050 3942
rect 4032 3942 4050 3960
rect 4032 3960 4050 3978
rect 4032 3978 4050 3996
rect 4032 3996 4050 4014
rect 4032 4014 4050 4032
rect 4032 4032 4050 4050
rect 4032 4050 4050 4068
rect 4032 4068 4050 4086
rect 4032 4086 4050 4104
rect 4032 4104 4050 4122
rect 4032 4122 4050 4140
rect 4032 4140 4050 4158
rect 4032 4158 4050 4176
rect 4032 4176 4050 4194
rect 4032 4194 4050 4212
rect 4032 4212 4050 4230
rect 4032 4230 4050 4248
rect 4032 4248 4050 4266
rect 4032 4266 4050 4284
rect 4032 4284 4050 4302
rect 4032 4302 4050 4320
rect 4032 4320 4050 4338
rect 4032 4338 4050 4356
rect 4032 4356 4050 4374
rect 4032 4374 4050 4392
rect 4032 4392 4050 4410
rect 4032 4410 4050 4428
rect 4032 4428 4050 4446
rect 4032 4446 4050 4464
rect 4032 4464 4050 4482
rect 4032 4482 4050 4500
rect 4032 4500 4050 4518
rect 4032 4518 4050 4536
rect 4032 4536 4050 4554
rect 4032 4554 4050 4572
rect 4032 4572 4050 4590
rect 4032 4590 4050 4608
rect 4032 4608 4050 4626
rect 4032 4626 4050 4644
rect 4032 4644 4050 4662
rect 4032 4662 4050 4680
rect 4032 4680 4050 4698
rect 4032 4698 4050 4716
rect 4032 4716 4050 4734
rect 4032 4734 4050 4752
rect 4032 4752 4050 4770
rect 4032 4770 4050 4788
rect 4032 4788 4050 4806
rect 4032 4806 4050 4824
rect 4032 4824 4050 4842
rect 4032 4842 4050 4860
rect 4032 4860 4050 4878
rect 4032 4878 4050 4896
rect 4032 4896 4050 4914
rect 4032 4914 4050 4932
rect 4032 4932 4050 4950
rect 4032 4950 4050 4968
rect 4032 4968 4050 4986
rect 4032 4986 4050 5004
rect 4032 5004 4050 5022
rect 4032 5022 4050 5040
rect 4032 5040 4050 5058
rect 4032 5058 4050 5076
rect 4032 5076 4050 5094
rect 4032 5094 4050 5112
rect 4032 5112 4050 5130
rect 4032 5130 4050 5148
rect 4032 5148 4050 5166
rect 4032 5166 4050 5184
rect 4032 5184 4050 5202
rect 4032 5202 4050 5220
rect 4032 5220 4050 5238
rect 4032 5238 4050 5256
rect 4032 5256 4050 5274
rect 4032 5274 4050 5292
rect 4032 5292 4050 5310
rect 4032 5310 4050 5328
rect 4032 5328 4050 5346
rect 4032 5346 4050 5364
rect 4032 5364 4050 5382
rect 4032 5382 4050 5400
rect 4032 5400 4050 5418
rect 4032 5418 4050 5436
rect 4032 5436 4050 5454
rect 4032 5454 4050 5472
rect 4032 5472 4050 5490
rect 4032 5490 4050 5508
rect 4032 5508 4050 5526
rect 4032 5526 4050 5544
rect 4032 5544 4050 5562
rect 4032 5562 4050 5580
rect 4032 5580 4050 5598
rect 4032 5598 4050 5616
rect 4032 5616 4050 5634
rect 4032 5634 4050 5652
rect 4032 5652 4050 5670
rect 4032 5670 4050 5688
rect 4032 5688 4050 5706
rect 4032 5706 4050 5724
rect 4032 5724 4050 5742
rect 4032 5742 4050 5760
rect 4032 5760 4050 5778
rect 4032 5778 4050 5796
rect 4032 5796 4050 5814
rect 4032 5814 4050 5832
rect 4032 5832 4050 5850
rect 4032 5850 4050 5868
rect 4032 5868 4050 5886
rect 4032 5886 4050 5904
rect 4032 5904 4050 5922
rect 4032 5922 4050 5940
rect 4032 5940 4050 5958
rect 4032 5958 4050 5976
rect 4032 5976 4050 5994
rect 4032 5994 4050 6012
rect 4032 6012 4050 6030
rect 4032 6030 4050 6048
rect 4032 6048 4050 6066
rect 4032 6066 4050 6084
rect 4032 6084 4050 6102
rect 4032 6102 4050 6120
rect 4032 6120 4050 6138
rect 4032 6138 4050 6156
rect 4032 6624 4050 6642
rect 4032 6642 4050 6660
rect 4032 6660 4050 6678
rect 4032 6678 4050 6696
rect 4032 6696 4050 6714
rect 4032 6714 4050 6732
rect 4032 6732 4050 6750
rect 4032 6750 4050 6768
rect 4032 6768 4050 6786
rect 4032 6786 4050 6804
rect 4032 6804 4050 6822
rect 4032 6822 4050 6840
rect 4032 6840 4050 6858
rect 4032 6858 4050 6876
rect 4032 6876 4050 6894
rect 4032 6894 4050 6912
rect 4032 6912 4050 6930
rect 4032 6930 4050 6948
rect 4032 6948 4050 6966
rect 4032 6966 4050 6984
rect 4032 6984 4050 7002
rect 4032 7002 4050 7020
rect 4032 7020 4050 7038
rect 4032 7038 4050 7056
rect 4032 7056 4050 7074
rect 4032 7074 4050 7092
rect 4032 7092 4050 7110
rect 4032 7110 4050 7128
rect 4032 7128 4050 7146
rect 4032 7146 4050 7164
rect 4032 7164 4050 7182
rect 4032 7182 4050 7200
rect 4032 7200 4050 7218
rect 4032 7218 4050 7236
rect 4032 7236 4050 7254
rect 4050 18 4068 36
rect 4050 36 4068 54
rect 4050 54 4068 72
rect 4050 72 4068 90
rect 4050 90 4068 108
rect 4050 108 4068 126
rect 4050 126 4068 144
rect 4050 144 4068 162
rect 4050 162 4068 180
rect 4050 180 4068 198
rect 4050 198 4068 216
rect 4050 216 4068 234
rect 4050 234 4068 252
rect 4050 252 4068 270
rect 4050 270 4068 288
rect 4050 288 4068 306
rect 4050 306 4068 324
rect 4050 324 4068 342
rect 4050 342 4068 360
rect 4050 360 4068 378
rect 4050 378 4068 396
rect 4050 396 4068 414
rect 4050 414 4068 432
rect 4050 432 4068 450
rect 4050 450 4068 468
rect 4050 468 4068 486
rect 4050 486 4068 504
rect 4050 504 4068 522
rect 4050 522 4068 540
rect 4050 540 4068 558
rect 4050 558 4068 576
rect 4050 576 4068 594
rect 4050 594 4068 612
rect 4050 612 4068 630
rect 4050 630 4068 648
rect 4050 864 4068 882
rect 4050 882 4068 900
rect 4050 900 4068 918
rect 4050 918 4068 936
rect 4050 936 4068 954
rect 4050 954 4068 972
rect 4050 972 4068 990
rect 4050 990 4068 1008
rect 4050 1008 4068 1026
rect 4050 1026 4068 1044
rect 4050 1044 4068 1062
rect 4050 1062 4068 1080
rect 4050 1080 4068 1098
rect 4050 1098 4068 1116
rect 4050 1116 4068 1134
rect 4050 1134 4068 1152
rect 4050 1152 4068 1170
rect 4050 1170 4068 1188
rect 4050 1188 4068 1206
rect 4050 1206 4068 1224
rect 4050 1224 4068 1242
rect 4050 1242 4068 1260
rect 4050 1260 4068 1278
rect 4050 1278 4068 1296
rect 4050 1296 4068 1314
rect 4050 1314 4068 1332
rect 4050 1332 4068 1350
rect 4050 1350 4068 1368
rect 4050 1368 4068 1386
rect 4050 1386 4068 1404
rect 4050 1404 4068 1422
rect 4050 1422 4068 1440
rect 4050 1440 4068 1458
rect 4050 1458 4068 1476
rect 4050 1476 4068 1494
rect 4050 1494 4068 1512
rect 4050 1512 4068 1530
rect 4050 1530 4068 1548
rect 4050 1548 4068 1566
rect 4050 1566 4068 1584
rect 4050 1584 4068 1602
rect 4050 1836 4068 1854
rect 4050 1854 4068 1872
rect 4050 1872 4068 1890
rect 4050 1890 4068 1908
rect 4050 1908 4068 1926
rect 4050 1926 4068 1944
rect 4050 1944 4068 1962
rect 4050 1962 4068 1980
rect 4050 1980 4068 1998
rect 4050 1998 4068 2016
rect 4050 2016 4068 2034
rect 4050 2034 4068 2052
rect 4050 2052 4068 2070
rect 4050 2070 4068 2088
rect 4050 2088 4068 2106
rect 4050 2106 4068 2124
rect 4050 2124 4068 2142
rect 4050 2142 4068 2160
rect 4050 2160 4068 2178
rect 4050 2178 4068 2196
rect 4050 2196 4068 2214
rect 4050 2214 4068 2232
rect 4050 2232 4068 2250
rect 4050 2250 4068 2268
rect 4050 2268 4068 2286
rect 4050 2286 4068 2304
rect 4050 2304 4068 2322
rect 4050 2322 4068 2340
rect 4050 2340 4068 2358
rect 4050 2358 4068 2376
rect 4050 2376 4068 2394
rect 4050 2394 4068 2412
rect 4050 2412 4068 2430
rect 4050 2430 4068 2448
rect 4050 2448 4068 2466
rect 4050 2466 4068 2484
rect 4050 2484 4068 2502
rect 4050 2502 4068 2520
rect 4050 2520 4068 2538
rect 4050 2538 4068 2556
rect 4050 2556 4068 2574
rect 4050 2574 4068 2592
rect 4050 2592 4068 2610
rect 4050 2610 4068 2628
rect 4050 2628 4068 2646
rect 4050 2646 4068 2664
rect 4050 2664 4068 2682
rect 4050 2682 4068 2700
rect 4050 2700 4068 2718
rect 4050 2718 4068 2736
rect 4050 2736 4068 2754
rect 4050 2754 4068 2772
rect 4050 2772 4068 2790
rect 4050 2790 4068 2808
rect 4050 2808 4068 2826
rect 4050 2826 4068 2844
rect 4050 2844 4068 2862
rect 4050 2862 4068 2880
rect 4050 2880 4068 2898
rect 4050 2898 4068 2916
rect 4050 2916 4068 2934
rect 4050 2934 4068 2952
rect 4050 2952 4068 2970
rect 4050 2970 4068 2988
rect 4050 2988 4068 3006
rect 4050 3006 4068 3024
rect 4050 3024 4068 3042
rect 4050 3042 4068 3060
rect 4050 3060 4068 3078
rect 4050 3078 4068 3096
rect 4050 3096 4068 3114
rect 4050 3114 4068 3132
rect 4050 3132 4068 3150
rect 4050 3150 4068 3168
rect 4050 3402 4068 3420
rect 4050 3420 4068 3438
rect 4050 3438 4068 3456
rect 4050 3456 4068 3474
rect 4050 3474 4068 3492
rect 4050 3492 4068 3510
rect 4050 3510 4068 3528
rect 4050 3528 4068 3546
rect 4050 3546 4068 3564
rect 4050 3564 4068 3582
rect 4050 3582 4068 3600
rect 4050 3600 4068 3618
rect 4050 3618 4068 3636
rect 4050 3636 4068 3654
rect 4050 3654 4068 3672
rect 4050 3672 4068 3690
rect 4050 3690 4068 3708
rect 4050 3708 4068 3726
rect 4050 3726 4068 3744
rect 4050 3744 4068 3762
rect 4050 3762 4068 3780
rect 4050 3780 4068 3798
rect 4050 3798 4068 3816
rect 4050 3816 4068 3834
rect 4050 3834 4068 3852
rect 4050 3852 4068 3870
rect 4050 3870 4068 3888
rect 4050 3888 4068 3906
rect 4050 3906 4068 3924
rect 4050 3924 4068 3942
rect 4050 3942 4068 3960
rect 4050 3960 4068 3978
rect 4050 3978 4068 3996
rect 4050 3996 4068 4014
rect 4050 4014 4068 4032
rect 4050 4032 4068 4050
rect 4050 4050 4068 4068
rect 4050 4068 4068 4086
rect 4050 4086 4068 4104
rect 4050 4104 4068 4122
rect 4050 4122 4068 4140
rect 4050 4140 4068 4158
rect 4050 4158 4068 4176
rect 4050 4176 4068 4194
rect 4050 4194 4068 4212
rect 4050 4212 4068 4230
rect 4050 4230 4068 4248
rect 4050 4248 4068 4266
rect 4050 4266 4068 4284
rect 4050 4284 4068 4302
rect 4050 4302 4068 4320
rect 4050 4320 4068 4338
rect 4050 4338 4068 4356
rect 4050 4356 4068 4374
rect 4050 4374 4068 4392
rect 4050 4392 4068 4410
rect 4050 4410 4068 4428
rect 4050 4428 4068 4446
rect 4050 4446 4068 4464
rect 4050 4464 4068 4482
rect 4050 4482 4068 4500
rect 4050 4500 4068 4518
rect 4050 4518 4068 4536
rect 4050 4536 4068 4554
rect 4050 4554 4068 4572
rect 4050 4572 4068 4590
rect 4050 4590 4068 4608
rect 4050 4608 4068 4626
rect 4050 4626 4068 4644
rect 4050 4644 4068 4662
rect 4050 4662 4068 4680
rect 4050 4680 4068 4698
rect 4050 4698 4068 4716
rect 4050 4716 4068 4734
rect 4050 4734 4068 4752
rect 4050 4752 4068 4770
rect 4050 4770 4068 4788
rect 4050 4788 4068 4806
rect 4050 4806 4068 4824
rect 4050 4824 4068 4842
rect 4050 4842 4068 4860
rect 4050 4860 4068 4878
rect 4050 4878 4068 4896
rect 4050 4896 4068 4914
rect 4050 4914 4068 4932
rect 4050 4932 4068 4950
rect 4050 4950 4068 4968
rect 4050 4968 4068 4986
rect 4050 4986 4068 5004
rect 4050 5004 4068 5022
rect 4050 5022 4068 5040
rect 4050 5040 4068 5058
rect 4050 5058 4068 5076
rect 4050 5076 4068 5094
rect 4050 5094 4068 5112
rect 4050 5112 4068 5130
rect 4050 5130 4068 5148
rect 4050 5148 4068 5166
rect 4050 5166 4068 5184
rect 4050 5184 4068 5202
rect 4050 5202 4068 5220
rect 4050 5220 4068 5238
rect 4050 5238 4068 5256
rect 4050 5256 4068 5274
rect 4050 5274 4068 5292
rect 4050 5292 4068 5310
rect 4050 5310 4068 5328
rect 4050 5328 4068 5346
rect 4050 5346 4068 5364
rect 4050 5364 4068 5382
rect 4050 5382 4068 5400
rect 4050 5400 4068 5418
rect 4050 5418 4068 5436
rect 4050 5436 4068 5454
rect 4050 5454 4068 5472
rect 4050 5472 4068 5490
rect 4050 5490 4068 5508
rect 4050 5508 4068 5526
rect 4050 5526 4068 5544
rect 4050 5544 4068 5562
rect 4050 5562 4068 5580
rect 4050 5580 4068 5598
rect 4050 5598 4068 5616
rect 4050 5616 4068 5634
rect 4050 5634 4068 5652
rect 4050 5652 4068 5670
rect 4050 5670 4068 5688
rect 4050 5688 4068 5706
rect 4050 5706 4068 5724
rect 4050 5724 4068 5742
rect 4050 5742 4068 5760
rect 4050 5760 4068 5778
rect 4050 5778 4068 5796
rect 4050 5796 4068 5814
rect 4050 5814 4068 5832
rect 4050 5832 4068 5850
rect 4050 5850 4068 5868
rect 4050 5868 4068 5886
rect 4050 5886 4068 5904
rect 4050 5904 4068 5922
rect 4050 5922 4068 5940
rect 4050 5940 4068 5958
rect 4050 5958 4068 5976
rect 4050 5976 4068 5994
rect 4050 5994 4068 6012
rect 4050 6012 4068 6030
rect 4050 6030 4068 6048
rect 4050 6048 4068 6066
rect 4050 6066 4068 6084
rect 4050 6084 4068 6102
rect 4050 6102 4068 6120
rect 4050 6120 4068 6138
rect 4050 6138 4068 6156
rect 4050 6156 4068 6174
rect 4050 6174 4068 6192
rect 4050 6624 4068 6642
rect 4050 6642 4068 6660
rect 4050 6660 4068 6678
rect 4050 6678 4068 6696
rect 4050 6696 4068 6714
rect 4050 6714 4068 6732
rect 4050 6732 4068 6750
rect 4050 6750 4068 6768
rect 4050 6768 4068 6786
rect 4050 6786 4068 6804
rect 4050 6804 4068 6822
rect 4050 6822 4068 6840
rect 4050 6840 4068 6858
rect 4050 6858 4068 6876
rect 4050 6876 4068 6894
rect 4050 6894 4068 6912
rect 4050 6912 4068 6930
rect 4050 6930 4068 6948
rect 4050 6948 4068 6966
rect 4050 6966 4068 6984
rect 4050 6984 4068 7002
rect 4050 7002 4068 7020
rect 4050 7020 4068 7038
rect 4050 7038 4068 7056
rect 4050 7056 4068 7074
rect 4050 7074 4068 7092
rect 4050 7092 4068 7110
rect 4050 7110 4068 7128
rect 4050 7128 4068 7146
rect 4050 7146 4068 7164
rect 4050 7164 4068 7182
rect 4050 7182 4068 7200
rect 4050 7200 4068 7218
rect 4050 7218 4068 7236
rect 4050 7236 4068 7254
rect 4068 18 4086 36
rect 4068 36 4086 54
rect 4068 54 4086 72
rect 4068 72 4086 90
rect 4068 90 4086 108
rect 4068 108 4086 126
rect 4068 126 4086 144
rect 4068 144 4086 162
rect 4068 162 4086 180
rect 4068 180 4086 198
rect 4068 198 4086 216
rect 4068 216 4086 234
rect 4068 234 4086 252
rect 4068 252 4086 270
rect 4068 270 4086 288
rect 4068 288 4086 306
rect 4068 306 4086 324
rect 4068 324 4086 342
rect 4068 342 4086 360
rect 4068 360 4086 378
rect 4068 378 4086 396
rect 4068 396 4086 414
rect 4068 414 4086 432
rect 4068 432 4086 450
rect 4068 450 4086 468
rect 4068 468 4086 486
rect 4068 486 4086 504
rect 4068 504 4086 522
rect 4068 522 4086 540
rect 4068 540 4086 558
rect 4068 558 4086 576
rect 4068 576 4086 594
rect 4068 594 4086 612
rect 4068 612 4086 630
rect 4068 630 4086 648
rect 4068 864 4086 882
rect 4068 882 4086 900
rect 4068 900 4086 918
rect 4068 918 4086 936
rect 4068 936 4086 954
rect 4068 954 4086 972
rect 4068 972 4086 990
rect 4068 990 4086 1008
rect 4068 1008 4086 1026
rect 4068 1026 4086 1044
rect 4068 1044 4086 1062
rect 4068 1062 4086 1080
rect 4068 1080 4086 1098
rect 4068 1098 4086 1116
rect 4068 1116 4086 1134
rect 4068 1134 4086 1152
rect 4068 1152 4086 1170
rect 4068 1170 4086 1188
rect 4068 1188 4086 1206
rect 4068 1206 4086 1224
rect 4068 1224 4086 1242
rect 4068 1242 4086 1260
rect 4068 1260 4086 1278
rect 4068 1278 4086 1296
rect 4068 1296 4086 1314
rect 4068 1314 4086 1332
rect 4068 1332 4086 1350
rect 4068 1350 4086 1368
rect 4068 1368 4086 1386
rect 4068 1386 4086 1404
rect 4068 1404 4086 1422
rect 4068 1422 4086 1440
rect 4068 1440 4086 1458
rect 4068 1458 4086 1476
rect 4068 1476 4086 1494
rect 4068 1494 4086 1512
rect 4068 1512 4086 1530
rect 4068 1530 4086 1548
rect 4068 1548 4086 1566
rect 4068 1566 4086 1584
rect 4068 1584 4086 1602
rect 4068 1602 4086 1620
rect 4068 1854 4086 1872
rect 4068 1872 4086 1890
rect 4068 1890 4086 1908
rect 4068 1908 4086 1926
rect 4068 1926 4086 1944
rect 4068 1944 4086 1962
rect 4068 1962 4086 1980
rect 4068 1980 4086 1998
rect 4068 1998 4086 2016
rect 4068 2016 4086 2034
rect 4068 2034 4086 2052
rect 4068 2052 4086 2070
rect 4068 2070 4086 2088
rect 4068 2088 4086 2106
rect 4068 2106 4086 2124
rect 4068 2124 4086 2142
rect 4068 2142 4086 2160
rect 4068 2160 4086 2178
rect 4068 2178 4086 2196
rect 4068 2196 4086 2214
rect 4068 2214 4086 2232
rect 4068 2232 4086 2250
rect 4068 2250 4086 2268
rect 4068 2268 4086 2286
rect 4068 2286 4086 2304
rect 4068 2304 4086 2322
rect 4068 2322 4086 2340
rect 4068 2340 4086 2358
rect 4068 2358 4086 2376
rect 4068 2376 4086 2394
rect 4068 2394 4086 2412
rect 4068 2412 4086 2430
rect 4068 2430 4086 2448
rect 4068 2448 4086 2466
rect 4068 2466 4086 2484
rect 4068 2484 4086 2502
rect 4068 2502 4086 2520
rect 4068 2520 4086 2538
rect 4068 2538 4086 2556
rect 4068 2556 4086 2574
rect 4068 2574 4086 2592
rect 4068 2592 4086 2610
rect 4068 2610 4086 2628
rect 4068 2628 4086 2646
rect 4068 2646 4086 2664
rect 4068 2664 4086 2682
rect 4068 2682 4086 2700
rect 4068 2700 4086 2718
rect 4068 2718 4086 2736
rect 4068 2736 4086 2754
rect 4068 2754 4086 2772
rect 4068 2772 4086 2790
rect 4068 2790 4086 2808
rect 4068 2808 4086 2826
rect 4068 2826 4086 2844
rect 4068 2844 4086 2862
rect 4068 2862 4086 2880
rect 4068 2880 4086 2898
rect 4068 2898 4086 2916
rect 4068 2916 4086 2934
rect 4068 2934 4086 2952
rect 4068 2952 4086 2970
rect 4068 2970 4086 2988
rect 4068 2988 4086 3006
rect 4068 3006 4086 3024
rect 4068 3024 4086 3042
rect 4068 3042 4086 3060
rect 4068 3060 4086 3078
rect 4068 3078 4086 3096
rect 4068 3096 4086 3114
rect 4068 3114 4086 3132
rect 4068 3132 4086 3150
rect 4068 3150 4086 3168
rect 4068 3168 4086 3186
rect 4068 3186 4086 3204
rect 4068 3420 4086 3438
rect 4068 3438 4086 3456
rect 4068 3456 4086 3474
rect 4068 3474 4086 3492
rect 4068 3492 4086 3510
rect 4068 3510 4086 3528
rect 4068 3528 4086 3546
rect 4068 3546 4086 3564
rect 4068 3564 4086 3582
rect 4068 3582 4086 3600
rect 4068 3600 4086 3618
rect 4068 3618 4086 3636
rect 4068 3636 4086 3654
rect 4068 3654 4086 3672
rect 4068 3672 4086 3690
rect 4068 3690 4086 3708
rect 4068 3708 4086 3726
rect 4068 3726 4086 3744
rect 4068 3744 4086 3762
rect 4068 3762 4086 3780
rect 4068 3780 4086 3798
rect 4068 3798 4086 3816
rect 4068 3816 4086 3834
rect 4068 3834 4086 3852
rect 4068 3852 4086 3870
rect 4068 3870 4086 3888
rect 4068 3888 4086 3906
rect 4068 3906 4086 3924
rect 4068 3924 4086 3942
rect 4068 3942 4086 3960
rect 4068 3960 4086 3978
rect 4068 3978 4086 3996
rect 4068 3996 4086 4014
rect 4068 4014 4086 4032
rect 4068 4032 4086 4050
rect 4068 4050 4086 4068
rect 4068 4068 4086 4086
rect 4068 4086 4086 4104
rect 4068 4104 4086 4122
rect 4068 4122 4086 4140
rect 4068 4140 4086 4158
rect 4068 4158 4086 4176
rect 4068 4176 4086 4194
rect 4068 4194 4086 4212
rect 4068 4212 4086 4230
rect 4068 4230 4086 4248
rect 4068 4248 4086 4266
rect 4068 4266 4086 4284
rect 4068 4284 4086 4302
rect 4068 4302 4086 4320
rect 4068 4320 4086 4338
rect 4068 4338 4086 4356
rect 4068 4356 4086 4374
rect 4068 4374 4086 4392
rect 4068 4392 4086 4410
rect 4068 4410 4086 4428
rect 4068 4428 4086 4446
rect 4068 4446 4086 4464
rect 4068 4464 4086 4482
rect 4068 4482 4086 4500
rect 4068 4500 4086 4518
rect 4068 4518 4086 4536
rect 4068 4536 4086 4554
rect 4068 4554 4086 4572
rect 4068 4572 4086 4590
rect 4068 4590 4086 4608
rect 4068 4608 4086 4626
rect 4068 4626 4086 4644
rect 4068 4644 4086 4662
rect 4068 4662 4086 4680
rect 4068 4680 4086 4698
rect 4068 4698 4086 4716
rect 4068 4716 4086 4734
rect 4068 4734 4086 4752
rect 4068 4752 4086 4770
rect 4068 4770 4086 4788
rect 4068 4788 4086 4806
rect 4068 4806 4086 4824
rect 4068 4824 4086 4842
rect 4068 4842 4086 4860
rect 4068 4860 4086 4878
rect 4068 4878 4086 4896
rect 4068 4896 4086 4914
rect 4068 4914 4086 4932
rect 4068 4932 4086 4950
rect 4068 4950 4086 4968
rect 4068 4968 4086 4986
rect 4068 4986 4086 5004
rect 4068 5004 4086 5022
rect 4068 5022 4086 5040
rect 4068 5040 4086 5058
rect 4068 5058 4086 5076
rect 4068 5076 4086 5094
rect 4068 5094 4086 5112
rect 4068 5112 4086 5130
rect 4068 5130 4086 5148
rect 4068 5148 4086 5166
rect 4068 5166 4086 5184
rect 4068 5184 4086 5202
rect 4068 5202 4086 5220
rect 4068 5220 4086 5238
rect 4068 5238 4086 5256
rect 4068 5256 4086 5274
rect 4068 5274 4086 5292
rect 4068 5292 4086 5310
rect 4068 5310 4086 5328
rect 4068 5328 4086 5346
rect 4068 5346 4086 5364
rect 4068 5364 4086 5382
rect 4068 5382 4086 5400
rect 4068 5400 4086 5418
rect 4068 5418 4086 5436
rect 4068 5436 4086 5454
rect 4068 5454 4086 5472
rect 4068 5472 4086 5490
rect 4068 5490 4086 5508
rect 4068 5508 4086 5526
rect 4068 5526 4086 5544
rect 4068 5544 4086 5562
rect 4068 5562 4086 5580
rect 4068 5580 4086 5598
rect 4068 5598 4086 5616
rect 4068 5616 4086 5634
rect 4068 5634 4086 5652
rect 4068 5652 4086 5670
rect 4068 5670 4086 5688
rect 4068 5688 4086 5706
rect 4068 5706 4086 5724
rect 4068 5724 4086 5742
rect 4068 5742 4086 5760
rect 4068 5760 4086 5778
rect 4068 5778 4086 5796
rect 4068 5796 4086 5814
rect 4068 5814 4086 5832
rect 4068 5832 4086 5850
rect 4068 5850 4086 5868
rect 4068 5868 4086 5886
rect 4068 5886 4086 5904
rect 4068 5904 4086 5922
rect 4068 5922 4086 5940
rect 4068 5940 4086 5958
rect 4068 5958 4086 5976
rect 4068 5976 4086 5994
rect 4068 5994 4086 6012
rect 4068 6012 4086 6030
rect 4068 6030 4086 6048
rect 4068 6048 4086 6066
rect 4068 6066 4086 6084
rect 4068 6084 4086 6102
rect 4068 6102 4086 6120
rect 4068 6120 4086 6138
rect 4068 6138 4086 6156
rect 4068 6156 4086 6174
rect 4068 6174 4086 6192
rect 4068 6192 4086 6210
rect 4068 6210 4086 6228
rect 4068 6624 4086 6642
rect 4068 6642 4086 6660
rect 4068 6660 4086 6678
rect 4068 6678 4086 6696
rect 4068 6696 4086 6714
rect 4068 6714 4086 6732
rect 4068 6732 4086 6750
rect 4068 6750 4086 6768
rect 4068 6768 4086 6786
rect 4068 6786 4086 6804
rect 4068 6804 4086 6822
rect 4068 6822 4086 6840
rect 4068 6840 4086 6858
rect 4068 6858 4086 6876
rect 4068 6876 4086 6894
rect 4068 6894 4086 6912
rect 4068 6912 4086 6930
rect 4068 6930 4086 6948
rect 4068 6948 4086 6966
rect 4068 6966 4086 6984
rect 4068 6984 4086 7002
rect 4068 7002 4086 7020
rect 4068 7020 4086 7038
rect 4068 7038 4086 7056
rect 4068 7056 4086 7074
rect 4068 7074 4086 7092
rect 4068 7092 4086 7110
rect 4068 7110 4086 7128
rect 4068 7128 4086 7146
rect 4068 7146 4086 7164
rect 4068 7164 4086 7182
rect 4068 7182 4086 7200
rect 4068 7200 4086 7218
rect 4068 7218 4086 7236
rect 4068 7236 4086 7254
rect 4086 18 4104 36
rect 4086 36 4104 54
rect 4086 54 4104 72
rect 4086 72 4104 90
rect 4086 90 4104 108
rect 4086 108 4104 126
rect 4086 126 4104 144
rect 4086 144 4104 162
rect 4086 162 4104 180
rect 4086 180 4104 198
rect 4086 198 4104 216
rect 4086 216 4104 234
rect 4086 234 4104 252
rect 4086 252 4104 270
rect 4086 270 4104 288
rect 4086 288 4104 306
rect 4086 306 4104 324
rect 4086 324 4104 342
rect 4086 342 4104 360
rect 4086 360 4104 378
rect 4086 378 4104 396
rect 4086 396 4104 414
rect 4086 414 4104 432
rect 4086 432 4104 450
rect 4086 450 4104 468
rect 4086 468 4104 486
rect 4086 486 4104 504
rect 4086 504 4104 522
rect 4086 522 4104 540
rect 4086 540 4104 558
rect 4086 558 4104 576
rect 4086 576 4104 594
rect 4086 594 4104 612
rect 4086 612 4104 630
rect 4086 630 4104 648
rect 4086 864 4104 882
rect 4086 882 4104 900
rect 4086 900 4104 918
rect 4086 918 4104 936
rect 4086 936 4104 954
rect 4086 954 4104 972
rect 4086 972 4104 990
rect 4086 990 4104 1008
rect 4086 1008 4104 1026
rect 4086 1026 4104 1044
rect 4086 1044 4104 1062
rect 4086 1062 4104 1080
rect 4086 1080 4104 1098
rect 4086 1098 4104 1116
rect 4086 1116 4104 1134
rect 4086 1134 4104 1152
rect 4086 1152 4104 1170
rect 4086 1170 4104 1188
rect 4086 1188 4104 1206
rect 4086 1206 4104 1224
rect 4086 1224 4104 1242
rect 4086 1242 4104 1260
rect 4086 1260 4104 1278
rect 4086 1278 4104 1296
rect 4086 1296 4104 1314
rect 4086 1314 4104 1332
rect 4086 1332 4104 1350
rect 4086 1350 4104 1368
rect 4086 1368 4104 1386
rect 4086 1386 4104 1404
rect 4086 1404 4104 1422
rect 4086 1422 4104 1440
rect 4086 1440 4104 1458
rect 4086 1458 4104 1476
rect 4086 1476 4104 1494
rect 4086 1494 4104 1512
rect 4086 1512 4104 1530
rect 4086 1530 4104 1548
rect 4086 1548 4104 1566
rect 4086 1566 4104 1584
rect 4086 1584 4104 1602
rect 4086 1602 4104 1620
rect 4086 1854 4104 1872
rect 4086 1872 4104 1890
rect 4086 1890 4104 1908
rect 4086 1908 4104 1926
rect 4086 1926 4104 1944
rect 4086 1944 4104 1962
rect 4086 1962 4104 1980
rect 4086 1980 4104 1998
rect 4086 1998 4104 2016
rect 4086 2016 4104 2034
rect 4086 2034 4104 2052
rect 4086 2052 4104 2070
rect 4086 2070 4104 2088
rect 4086 2088 4104 2106
rect 4086 2106 4104 2124
rect 4086 2124 4104 2142
rect 4086 2142 4104 2160
rect 4086 2160 4104 2178
rect 4086 2178 4104 2196
rect 4086 2196 4104 2214
rect 4086 2214 4104 2232
rect 4086 2232 4104 2250
rect 4086 2250 4104 2268
rect 4086 2268 4104 2286
rect 4086 2286 4104 2304
rect 4086 2304 4104 2322
rect 4086 2322 4104 2340
rect 4086 2340 4104 2358
rect 4086 2358 4104 2376
rect 4086 2376 4104 2394
rect 4086 2394 4104 2412
rect 4086 2412 4104 2430
rect 4086 2430 4104 2448
rect 4086 2448 4104 2466
rect 4086 2466 4104 2484
rect 4086 2484 4104 2502
rect 4086 2502 4104 2520
rect 4086 2520 4104 2538
rect 4086 2538 4104 2556
rect 4086 2556 4104 2574
rect 4086 2574 4104 2592
rect 4086 2592 4104 2610
rect 4086 2610 4104 2628
rect 4086 2628 4104 2646
rect 4086 2646 4104 2664
rect 4086 2664 4104 2682
rect 4086 2682 4104 2700
rect 4086 2700 4104 2718
rect 4086 2718 4104 2736
rect 4086 2736 4104 2754
rect 4086 2754 4104 2772
rect 4086 2772 4104 2790
rect 4086 2790 4104 2808
rect 4086 2808 4104 2826
rect 4086 2826 4104 2844
rect 4086 2844 4104 2862
rect 4086 2862 4104 2880
rect 4086 2880 4104 2898
rect 4086 2898 4104 2916
rect 4086 2916 4104 2934
rect 4086 2934 4104 2952
rect 4086 2952 4104 2970
rect 4086 2970 4104 2988
rect 4086 2988 4104 3006
rect 4086 3006 4104 3024
rect 4086 3024 4104 3042
rect 4086 3042 4104 3060
rect 4086 3060 4104 3078
rect 4086 3078 4104 3096
rect 4086 3096 4104 3114
rect 4086 3114 4104 3132
rect 4086 3132 4104 3150
rect 4086 3150 4104 3168
rect 4086 3168 4104 3186
rect 4086 3186 4104 3204
rect 4086 3204 4104 3222
rect 4086 3438 4104 3456
rect 4086 3456 4104 3474
rect 4086 3474 4104 3492
rect 4086 3492 4104 3510
rect 4086 3510 4104 3528
rect 4086 3528 4104 3546
rect 4086 3546 4104 3564
rect 4086 3564 4104 3582
rect 4086 3582 4104 3600
rect 4086 3600 4104 3618
rect 4086 3618 4104 3636
rect 4086 3636 4104 3654
rect 4086 3654 4104 3672
rect 4086 3672 4104 3690
rect 4086 3690 4104 3708
rect 4086 3708 4104 3726
rect 4086 3726 4104 3744
rect 4086 3744 4104 3762
rect 4086 3762 4104 3780
rect 4086 3780 4104 3798
rect 4086 3798 4104 3816
rect 4086 3816 4104 3834
rect 4086 3834 4104 3852
rect 4086 3852 4104 3870
rect 4086 3870 4104 3888
rect 4086 3888 4104 3906
rect 4086 3906 4104 3924
rect 4086 3924 4104 3942
rect 4086 3942 4104 3960
rect 4086 3960 4104 3978
rect 4086 3978 4104 3996
rect 4086 3996 4104 4014
rect 4086 4014 4104 4032
rect 4086 4032 4104 4050
rect 4086 4050 4104 4068
rect 4086 4068 4104 4086
rect 4086 4086 4104 4104
rect 4086 4104 4104 4122
rect 4086 4122 4104 4140
rect 4086 4140 4104 4158
rect 4086 4158 4104 4176
rect 4086 4176 4104 4194
rect 4086 4194 4104 4212
rect 4086 4212 4104 4230
rect 4086 4230 4104 4248
rect 4086 4248 4104 4266
rect 4086 4266 4104 4284
rect 4086 4284 4104 4302
rect 4086 4302 4104 4320
rect 4086 4320 4104 4338
rect 4086 4338 4104 4356
rect 4086 4356 4104 4374
rect 4086 4374 4104 4392
rect 4086 4392 4104 4410
rect 4086 4410 4104 4428
rect 4086 4428 4104 4446
rect 4086 4446 4104 4464
rect 4086 4464 4104 4482
rect 4086 4482 4104 4500
rect 4086 4500 4104 4518
rect 4086 4518 4104 4536
rect 4086 4536 4104 4554
rect 4086 4554 4104 4572
rect 4086 4572 4104 4590
rect 4086 4590 4104 4608
rect 4086 4608 4104 4626
rect 4086 4626 4104 4644
rect 4086 4644 4104 4662
rect 4086 4662 4104 4680
rect 4086 4680 4104 4698
rect 4086 4698 4104 4716
rect 4086 4716 4104 4734
rect 4086 4734 4104 4752
rect 4086 4752 4104 4770
rect 4086 4770 4104 4788
rect 4086 4788 4104 4806
rect 4086 4806 4104 4824
rect 4086 4824 4104 4842
rect 4086 4842 4104 4860
rect 4086 4860 4104 4878
rect 4086 4878 4104 4896
rect 4086 4896 4104 4914
rect 4086 4914 4104 4932
rect 4086 4932 4104 4950
rect 4086 4950 4104 4968
rect 4086 4968 4104 4986
rect 4086 4986 4104 5004
rect 4086 5004 4104 5022
rect 4086 5022 4104 5040
rect 4086 5040 4104 5058
rect 4086 5058 4104 5076
rect 4086 5076 4104 5094
rect 4086 5094 4104 5112
rect 4086 5112 4104 5130
rect 4086 5130 4104 5148
rect 4086 5148 4104 5166
rect 4086 5166 4104 5184
rect 4086 5184 4104 5202
rect 4086 5202 4104 5220
rect 4086 5220 4104 5238
rect 4086 5238 4104 5256
rect 4086 5256 4104 5274
rect 4086 5274 4104 5292
rect 4086 5292 4104 5310
rect 4086 5310 4104 5328
rect 4086 5328 4104 5346
rect 4086 5346 4104 5364
rect 4086 5364 4104 5382
rect 4086 5382 4104 5400
rect 4086 5400 4104 5418
rect 4086 5418 4104 5436
rect 4086 5436 4104 5454
rect 4086 5454 4104 5472
rect 4086 5472 4104 5490
rect 4086 5490 4104 5508
rect 4086 5508 4104 5526
rect 4086 5526 4104 5544
rect 4086 5544 4104 5562
rect 4086 5562 4104 5580
rect 4086 5580 4104 5598
rect 4086 5598 4104 5616
rect 4086 5616 4104 5634
rect 4086 5634 4104 5652
rect 4086 5652 4104 5670
rect 4086 5670 4104 5688
rect 4086 5688 4104 5706
rect 4086 5706 4104 5724
rect 4086 5724 4104 5742
rect 4086 5742 4104 5760
rect 4086 5760 4104 5778
rect 4086 5778 4104 5796
rect 4086 5796 4104 5814
rect 4086 5814 4104 5832
rect 4086 5832 4104 5850
rect 4086 5850 4104 5868
rect 4086 5868 4104 5886
rect 4086 5886 4104 5904
rect 4086 5904 4104 5922
rect 4086 5922 4104 5940
rect 4086 5940 4104 5958
rect 4086 5958 4104 5976
rect 4086 5976 4104 5994
rect 4086 5994 4104 6012
rect 4086 6012 4104 6030
rect 4086 6030 4104 6048
rect 4086 6048 4104 6066
rect 4086 6066 4104 6084
rect 4086 6084 4104 6102
rect 4086 6102 4104 6120
rect 4086 6120 4104 6138
rect 4086 6138 4104 6156
rect 4086 6156 4104 6174
rect 4086 6174 4104 6192
rect 4086 6192 4104 6210
rect 4086 6210 4104 6228
rect 4086 6228 4104 6246
rect 4086 6246 4104 6264
rect 4086 6624 4104 6642
rect 4086 6642 4104 6660
rect 4086 6660 4104 6678
rect 4086 6678 4104 6696
rect 4086 6696 4104 6714
rect 4086 6714 4104 6732
rect 4086 6732 4104 6750
rect 4086 6750 4104 6768
rect 4086 6768 4104 6786
rect 4086 6786 4104 6804
rect 4086 6804 4104 6822
rect 4086 6822 4104 6840
rect 4086 6840 4104 6858
rect 4086 6858 4104 6876
rect 4086 6876 4104 6894
rect 4086 6894 4104 6912
rect 4086 6912 4104 6930
rect 4086 6930 4104 6948
rect 4086 6948 4104 6966
rect 4086 6966 4104 6984
rect 4086 6984 4104 7002
rect 4086 7002 4104 7020
rect 4086 7020 4104 7038
rect 4086 7038 4104 7056
rect 4086 7056 4104 7074
rect 4086 7074 4104 7092
rect 4086 7092 4104 7110
rect 4086 7110 4104 7128
rect 4086 7128 4104 7146
rect 4086 7146 4104 7164
rect 4086 7164 4104 7182
rect 4086 7182 4104 7200
rect 4086 7200 4104 7218
rect 4086 7218 4104 7236
rect 4086 7236 4104 7254
rect 4104 36 4122 54
rect 4104 54 4122 72
rect 4104 72 4122 90
rect 4104 90 4122 108
rect 4104 108 4122 126
rect 4104 126 4122 144
rect 4104 144 4122 162
rect 4104 162 4122 180
rect 4104 180 4122 198
rect 4104 198 4122 216
rect 4104 216 4122 234
rect 4104 234 4122 252
rect 4104 252 4122 270
rect 4104 270 4122 288
rect 4104 288 4122 306
rect 4104 306 4122 324
rect 4104 324 4122 342
rect 4104 342 4122 360
rect 4104 360 4122 378
rect 4104 378 4122 396
rect 4104 396 4122 414
rect 4104 414 4122 432
rect 4104 432 4122 450
rect 4104 450 4122 468
rect 4104 468 4122 486
rect 4104 486 4122 504
rect 4104 504 4122 522
rect 4104 522 4122 540
rect 4104 540 4122 558
rect 4104 558 4122 576
rect 4104 576 4122 594
rect 4104 594 4122 612
rect 4104 612 4122 630
rect 4104 630 4122 648
rect 4104 864 4122 882
rect 4104 882 4122 900
rect 4104 900 4122 918
rect 4104 918 4122 936
rect 4104 936 4122 954
rect 4104 954 4122 972
rect 4104 972 4122 990
rect 4104 990 4122 1008
rect 4104 1008 4122 1026
rect 4104 1026 4122 1044
rect 4104 1044 4122 1062
rect 4104 1062 4122 1080
rect 4104 1080 4122 1098
rect 4104 1098 4122 1116
rect 4104 1116 4122 1134
rect 4104 1134 4122 1152
rect 4104 1152 4122 1170
rect 4104 1170 4122 1188
rect 4104 1188 4122 1206
rect 4104 1206 4122 1224
rect 4104 1224 4122 1242
rect 4104 1242 4122 1260
rect 4104 1260 4122 1278
rect 4104 1278 4122 1296
rect 4104 1296 4122 1314
rect 4104 1314 4122 1332
rect 4104 1332 4122 1350
rect 4104 1350 4122 1368
rect 4104 1368 4122 1386
rect 4104 1386 4122 1404
rect 4104 1404 4122 1422
rect 4104 1422 4122 1440
rect 4104 1440 4122 1458
rect 4104 1458 4122 1476
rect 4104 1476 4122 1494
rect 4104 1494 4122 1512
rect 4104 1512 4122 1530
rect 4104 1530 4122 1548
rect 4104 1548 4122 1566
rect 4104 1566 4122 1584
rect 4104 1584 4122 1602
rect 4104 1602 4122 1620
rect 4104 1620 4122 1638
rect 4104 1872 4122 1890
rect 4104 1890 4122 1908
rect 4104 1908 4122 1926
rect 4104 1926 4122 1944
rect 4104 1944 4122 1962
rect 4104 1962 4122 1980
rect 4104 1980 4122 1998
rect 4104 1998 4122 2016
rect 4104 2016 4122 2034
rect 4104 2034 4122 2052
rect 4104 2052 4122 2070
rect 4104 2070 4122 2088
rect 4104 2088 4122 2106
rect 4104 2106 4122 2124
rect 4104 2124 4122 2142
rect 4104 2142 4122 2160
rect 4104 2160 4122 2178
rect 4104 2178 4122 2196
rect 4104 2196 4122 2214
rect 4104 2214 4122 2232
rect 4104 2232 4122 2250
rect 4104 2250 4122 2268
rect 4104 2268 4122 2286
rect 4104 2286 4122 2304
rect 4104 2304 4122 2322
rect 4104 2322 4122 2340
rect 4104 2340 4122 2358
rect 4104 2358 4122 2376
rect 4104 2376 4122 2394
rect 4104 2394 4122 2412
rect 4104 2412 4122 2430
rect 4104 2430 4122 2448
rect 4104 2448 4122 2466
rect 4104 2466 4122 2484
rect 4104 2484 4122 2502
rect 4104 2502 4122 2520
rect 4104 2520 4122 2538
rect 4104 2538 4122 2556
rect 4104 2556 4122 2574
rect 4104 2574 4122 2592
rect 4104 2592 4122 2610
rect 4104 2610 4122 2628
rect 4104 2628 4122 2646
rect 4104 2646 4122 2664
rect 4104 2664 4122 2682
rect 4104 2682 4122 2700
rect 4104 2700 4122 2718
rect 4104 2718 4122 2736
rect 4104 2736 4122 2754
rect 4104 2754 4122 2772
rect 4104 2772 4122 2790
rect 4104 2790 4122 2808
rect 4104 2808 4122 2826
rect 4104 2826 4122 2844
rect 4104 2844 4122 2862
rect 4104 2862 4122 2880
rect 4104 2880 4122 2898
rect 4104 2898 4122 2916
rect 4104 2916 4122 2934
rect 4104 2934 4122 2952
rect 4104 2952 4122 2970
rect 4104 2970 4122 2988
rect 4104 2988 4122 3006
rect 4104 3006 4122 3024
rect 4104 3024 4122 3042
rect 4104 3042 4122 3060
rect 4104 3060 4122 3078
rect 4104 3078 4122 3096
rect 4104 3096 4122 3114
rect 4104 3114 4122 3132
rect 4104 3132 4122 3150
rect 4104 3150 4122 3168
rect 4104 3168 4122 3186
rect 4104 3186 4122 3204
rect 4104 3204 4122 3222
rect 4104 3222 4122 3240
rect 4104 3240 4122 3258
rect 4104 3474 4122 3492
rect 4104 3492 4122 3510
rect 4104 3510 4122 3528
rect 4104 3528 4122 3546
rect 4104 3546 4122 3564
rect 4104 3564 4122 3582
rect 4104 3582 4122 3600
rect 4104 3600 4122 3618
rect 4104 3618 4122 3636
rect 4104 3636 4122 3654
rect 4104 3654 4122 3672
rect 4104 3672 4122 3690
rect 4104 3690 4122 3708
rect 4104 3708 4122 3726
rect 4104 3726 4122 3744
rect 4104 3744 4122 3762
rect 4104 3762 4122 3780
rect 4104 3780 4122 3798
rect 4104 3798 4122 3816
rect 4104 3816 4122 3834
rect 4104 3834 4122 3852
rect 4104 3852 4122 3870
rect 4104 3870 4122 3888
rect 4104 3888 4122 3906
rect 4104 3906 4122 3924
rect 4104 3924 4122 3942
rect 4104 3942 4122 3960
rect 4104 3960 4122 3978
rect 4104 3978 4122 3996
rect 4104 3996 4122 4014
rect 4104 4014 4122 4032
rect 4104 4032 4122 4050
rect 4104 4050 4122 4068
rect 4104 4068 4122 4086
rect 4104 4086 4122 4104
rect 4104 4104 4122 4122
rect 4104 4122 4122 4140
rect 4104 4140 4122 4158
rect 4104 4158 4122 4176
rect 4104 4176 4122 4194
rect 4104 4194 4122 4212
rect 4104 4212 4122 4230
rect 4104 4230 4122 4248
rect 4104 4248 4122 4266
rect 4104 4266 4122 4284
rect 4104 4284 4122 4302
rect 4104 4302 4122 4320
rect 4104 4320 4122 4338
rect 4104 4338 4122 4356
rect 4104 4356 4122 4374
rect 4104 4374 4122 4392
rect 4104 4392 4122 4410
rect 4104 4410 4122 4428
rect 4104 4428 4122 4446
rect 4104 4446 4122 4464
rect 4104 4464 4122 4482
rect 4104 4482 4122 4500
rect 4104 4500 4122 4518
rect 4104 4518 4122 4536
rect 4104 4536 4122 4554
rect 4104 4554 4122 4572
rect 4104 4572 4122 4590
rect 4104 4590 4122 4608
rect 4104 4608 4122 4626
rect 4104 4626 4122 4644
rect 4104 4644 4122 4662
rect 4104 4662 4122 4680
rect 4104 4680 4122 4698
rect 4104 4698 4122 4716
rect 4104 4716 4122 4734
rect 4104 4734 4122 4752
rect 4104 4752 4122 4770
rect 4104 4770 4122 4788
rect 4104 4788 4122 4806
rect 4104 4806 4122 4824
rect 4104 4824 4122 4842
rect 4104 4842 4122 4860
rect 4104 4860 4122 4878
rect 4104 4878 4122 4896
rect 4104 4896 4122 4914
rect 4104 4914 4122 4932
rect 4104 4932 4122 4950
rect 4104 4950 4122 4968
rect 4104 4968 4122 4986
rect 4104 4986 4122 5004
rect 4104 5004 4122 5022
rect 4104 5022 4122 5040
rect 4104 5040 4122 5058
rect 4104 5058 4122 5076
rect 4104 5076 4122 5094
rect 4104 5094 4122 5112
rect 4104 5112 4122 5130
rect 4104 5130 4122 5148
rect 4104 5148 4122 5166
rect 4104 5166 4122 5184
rect 4104 5184 4122 5202
rect 4104 5202 4122 5220
rect 4104 5220 4122 5238
rect 4104 5238 4122 5256
rect 4104 5256 4122 5274
rect 4104 5274 4122 5292
rect 4104 5292 4122 5310
rect 4104 5310 4122 5328
rect 4104 5328 4122 5346
rect 4104 5346 4122 5364
rect 4104 5364 4122 5382
rect 4104 5382 4122 5400
rect 4104 5400 4122 5418
rect 4104 5418 4122 5436
rect 4104 5436 4122 5454
rect 4104 5454 4122 5472
rect 4104 5472 4122 5490
rect 4104 5490 4122 5508
rect 4104 5508 4122 5526
rect 4104 5526 4122 5544
rect 4104 5544 4122 5562
rect 4104 5562 4122 5580
rect 4104 5580 4122 5598
rect 4104 5598 4122 5616
rect 4104 5616 4122 5634
rect 4104 5634 4122 5652
rect 4104 5652 4122 5670
rect 4104 5670 4122 5688
rect 4104 5688 4122 5706
rect 4104 5706 4122 5724
rect 4104 5724 4122 5742
rect 4104 5742 4122 5760
rect 4104 5760 4122 5778
rect 4104 5778 4122 5796
rect 4104 5796 4122 5814
rect 4104 5814 4122 5832
rect 4104 5832 4122 5850
rect 4104 5850 4122 5868
rect 4104 5868 4122 5886
rect 4104 5886 4122 5904
rect 4104 5904 4122 5922
rect 4104 5922 4122 5940
rect 4104 5940 4122 5958
rect 4104 5958 4122 5976
rect 4104 5976 4122 5994
rect 4104 5994 4122 6012
rect 4104 6012 4122 6030
rect 4104 6030 4122 6048
rect 4104 6048 4122 6066
rect 4104 6066 4122 6084
rect 4104 6084 4122 6102
rect 4104 6102 4122 6120
rect 4104 6120 4122 6138
rect 4104 6138 4122 6156
rect 4104 6156 4122 6174
rect 4104 6174 4122 6192
rect 4104 6192 4122 6210
rect 4104 6210 4122 6228
rect 4104 6228 4122 6246
rect 4104 6246 4122 6264
rect 4104 6264 4122 6282
rect 4104 6282 4122 6300
rect 4104 6642 4122 6660
rect 4104 6660 4122 6678
rect 4104 6678 4122 6696
rect 4104 6696 4122 6714
rect 4104 6714 4122 6732
rect 4104 6732 4122 6750
rect 4104 6750 4122 6768
rect 4104 6768 4122 6786
rect 4104 6786 4122 6804
rect 4104 6804 4122 6822
rect 4104 6822 4122 6840
rect 4104 6840 4122 6858
rect 4104 6858 4122 6876
rect 4104 6876 4122 6894
rect 4104 6894 4122 6912
rect 4104 6912 4122 6930
rect 4104 6930 4122 6948
rect 4104 6948 4122 6966
rect 4104 6966 4122 6984
rect 4104 6984 4122 7002
rect 4104 7002 4122 7020
rect 4104 7020 4122 7038
rect 4104 7038 4122 7056
rect 4104 7056 4122 7074
rect 4104 7074 4122 7092
rect 4104 7092 4122 7110
rect 4104 7110 4122 7128
rect 4104 7128 4122 7146
rect 4104 7146 4122 7164
rect 4104 7164 4122 7182
rect 4104 7182 4122 7200
rect 4104 7200 4122 7218
rect 4104 7218 4122 7236
rect 4122 36 4140 54
rect 4122 54 4140 72
rect 4122 72 4140 90
rect 4122 90 4140 108
rect 4122 108 4140 126
rect 4122 126 4140 144
rect 4122 144 4140 162
rect 4122 162 4140 180
rect 4122 180 4140 198
rect 4122 198 4140 216
rect 4122 216 4140 234
rect 4122 234 4140 252
rect 4122 252 4140 270
rect 4122 270 4140 288
rect 4122 288 4140 306
rect 4122 306 4140 324
rect 4122 324 4140 342
rect 4122 342 4140 360
rect 4122 360 4140 378
rect 4122 378 4140 396
rect 4122 396 4140 414
rect 4122 414 4140 432
rect 4122 432 4140 450
rect 4122 450 4140 468
rect 4122 468 4140 486
rect 4122 486 4140 504
rect 4122 504 4140 522
rect 4122 522 4140 540
rect 4122 540 4140 558
rect 4122 558 4140 576
rect 4122 576 4140 594
rect 4122 594 4140 612
rect 4122 612 4140 630
rect 4122 630 4140 648
rect 4122 648 4140 666
rect 4122 864 4140 882
rect 4122 882 4140 900
rect 4122 900 4140 918
rect 4122 918 4140 936
rect 4122 936 4140 954
rect 4122 954 4140 972
rect 4122 972 4140 990
rect 4122 990 4140 1008
rect 4122 1008 4140 1026
rect 4122 1026 4140 1044
rect 4122 1044 4140 1062
rect 4122 1062 4140 1080
rect 4122 1080 4140 1098
rect 4122 1098 4140 1116
rect 4122 1116 4140 1134
rect 4122 1134 4140 1152
rect 4122 1152 4140 1170
rect 4122 1170 4140 1188
rect 4122 1188 4140 1206
rect 4122 1206 4140 1224
rect 4122 1224 4140 1242
rect 4122 1242 4140 1260
rect 4122 1260 4140 1278
rect 4122 1278 4140 1296
rect 4122 1296 4140 1314
rect 4122 1314 4140 1332
rect 4122 1332 4140 1350
rect 4122 1350 4140 1368
rect 4122 1368 4140 1386
rect 4122 1386 4140 1404
rect 4122 1404 4140 1422
rect 4122 1422 4140 1440
rect 4122 1440 4140 1458
rect 4122 1458 4140 1476
rect 4122 1476 4140 1494
rect 4122 1494 4140 1512
rect 4122 1512 4140 1530
rect 4122 1530 4140 1548
rect 4122 1548 4140 1566
rect 4122 1566 4140 1584
rect 4122 1584 4140 1602
rect 4122 1602 4140 1620
rect 4122 1620 4140 1638
rect 4122 1638 4140 1656
rect 4122 1890 4140 1908
rect 4122 1908 4140 1926
rect 4122 1926 4140 1944
rect 4122 1944 4140 1962
rect 4122 1962 4140 1980
rect 4122 1980 4140 1998
rect 4122 1998 4140 2016
rect 4122 2016 4140 2034
rect 4122 2034 4140 2052
rect 4122 2052 4140 2070
rect 4122 2070 4140 2088
rect 4122 2088 4140 2106
rect 4122 2106 4140 2124
rect 4122 2124 4140 2142
rect 4122 2142 4140 2160
rect 4122 2160 4140 2178
rect 4122 2178 4140 2196
rect 4122 2196 4140 2214
rect 4122 2214 4140 2232
rect 4122 2232 4140 2250
rect 4122 2250 4140 2268
rect 4122 2268 4140 2286
rect 4122 2286 4140 2304
rect 4122 2304 4140 2322
rect 4122 2322 4140 2340
rect 4122 2340 4140 2358
rect 4122 2358 4140 2376
rect 4122 2376 4140 2394
rect 4122 2394 4140 2412
rect 4122 2412 4140 2430
rect 4122 2430 4140 2448
rect 4122 2448 4140 2466
rect 4122 2466 4140 2484
rect 4122 2484 4140 2502
rect 4122 2502 4140 2520
rect 4122 2520 4140 2538
rect 4122 2538 4140 2556
rect 4122 2556 4140 2574
rect 4122 2574 4140 2592
rect 4122 2592 4140 2610
rect 4122 2610 4140 2628
rect 4122 2628 4140 2646
rect 4122 2646 4140 2664
rect 4122 2664 4140 2682
rect 4122 2682 4140 2700
rect 4122 2700 4140 2718
rect 4122 2718 4140 2736
rect 4122 2736 4140 2754
rect 4122 2754 4140 2772
rect 4122 2772 4140 2790
rect 4122 2790 4140 2808
rect 4122 2808 4140 2826
rect 4122 2826 4140 2844
rect 4122 2844 4140 2862
rect 4122 2862 4140 2880
rect 4122 2880 4140 2898
rect 4122 2898 4140 2916
rect 4122 2916 4140 2934
rect 4122 2934 4140 2952
rect 4122 2952 4140 2970
rect 4122 2970 4140 2988
rect 4122 2988 4140 3006
rect 4122 3006 4140 3024
rect 4122 3024 4140 3042
rect 4122 3042 4140 3060
rect 4122 3060 4140 3078
rect 4122 3078 4140 3096
rect 4122 3096 4140 3114
rect 4122 3114 4140 3132
rect 4122 3132 4140 3150
rect 4122 3150 4140 3168
rect 4122 3168 4140 3186
rect 4122 3186 4140 3204
rect 4122 3204 4140 3222
rect 4122 3222 4140 3240
rect 4122 3240 4140 3258
rect 4122 3258 4140 3276
rect 4122 3492 4140 3510
rect 4122 3510 4140 3528
rect 4122 3528 4140 3546
rect 4122 3546 4140 3564
rect 4122 3564 4140 3582
rect 4122 3582 4140 3600
rect 4122 3600 4140 3618
rect 4122 3618 4140 3636
rect 4122 3636 4140 3654
rect 4122 3654 4140 3672
rect 4122 3672 4140 3690
rect 4122 3690 4140 3708
rect 4122 3708 4140 3726
rect 4122 3726 4140 3744
rect 4122 3744 4140 3762
rect 4122 3762 4140 3780
rect 4122 3780 4140 3798
rect 4122 3798 4140 3816
rect 4122 3816 4140 3834
rect 4122 3834 4140 3852
rect 4122 3852 4140 3870
rect 4122 3870 4140 3888
rect 4122 3888 4140 3906
rect 4122 3906 4140 3924
rect 4122 3924 4140 3942
rect 4122 3942 4140 3960
rect 4122 3960 4140 3978
rect 4122 3978 4140 3996
rect 4122 3996 4140 4014
rect 4122 4014 4140 4032
rect 4122 4032 4140 4050
rect 4122 4050 4140 4068
rect 4122 4068 4140 4086
rect 4122 4086 4140 4104
rect 4122 4104 4140 4122
rect 4122 4122 4140 4140
rect 4122 4140 4140 4158
rect 4122 4158 4140 4176
rect 4122 4176 4140 4194
rect 4122 4194 4140 4212
rect 4122 4212 4140 4230
rect 4122 4230 4140 4248
rect 4122 4248 4140 4266
rect 4122 4266 4140 4284
rect 4122 4284 4140 4302
rect 4122 4302 4140 4320
rect 4122 4320 4140 4338
rect 4122 4338 4140 4356
rect 4122 4356 4140 4374
rect 4122 4374 4140 4392
rect 4122 4392 4140 4410
rect 4122 4410 4140 4428
rect 4122 4428 4140 4446
rect 4122 4446 4140 4464
rect 4122 4464 4140 4482
rect 4122 4482 4140 4500
rect 4122 4500 4140 4518
rect 4122 4518 4140 4536
rect 4122 4536 4140 4554
rect 4122 4554 4140 4572
rect 4122 4572 4140 4590
rect 4122 4590 4140 4608
rect 4122 4608 4140 4626
rect 4122 4626 4140 4644
rect 4122 4644 4140 4662
rect 4122 4662 4140 4680
rect 4122 4680 4140 4698
rect 4122 4698 4140 4716
rect 4122 4716 4140 4734
rect 4122 4734 4140 4752
rect 4122 4752 4140 4770
rect 4122 4770 4140 4788
rect 4122 4788 4140 4806
rect 4122 4806 4140 4824
rect 4122 4824 4140 4842
rect 4122 4842 4140 4860
rect 4122 4860 4140 4878
rect 4122 4878 4140 4896
rect 4122 4896 4140 4914
rect 4122 4914 4140 4932
rect 4122 4932 4140 4950
rect 4122 4950 4140 4968
rect 4122 4968 4140 4986
rect 4122 4986 4140 5004
rect 4122 5004 4140 5022
rect 4122 5022 4140 5040
rect 4122 5040 4140 5058
rect 4122 5058 4140 5076
rect 4122 5076 4140 5094
rect 4122 5094 4140 5112
rect 4122 5112 4140 5130
rect 4122 5130 4140 5148
rect 4122 5148 4140 5166
rect 4122 5166 4140 5184
rect 4122 5184 4140 5202
rect 4122 5202 4140 5220
rect 4122 5220 4140 5238
rect 4122 5238 4140 5256
rect 4122 5256 4140 5274
rect 4122 5274 4140 5292
rect 4122 5292 4140 5310
rect 4122 5310 4140 5328
rect 4122 5328 4140 5346
rect 4122 5346 4140 5364
rect 4122 5364 4140 5382
rect 4122 5382 4140 5400
rect 4122 5400 4140 5418
rect 4122 5418 4140 5436
rect 4122 5436 4140 5454
rect 4122 5454 4140 5472
rect 4122 5472 4140 5490
rect 4122 5490 4140 5508
rect 4122 5508 4140 5526
rect 4122 5526 4140 5544
rect 4122 5544 4140 5562
rect 4122 5562 4140 5580
rect 4122 5580 4140 5598
rect 4122 5598 4140 5616
rect 4122 5616 4140 5634
rect 4122 5634 4140 5652
rect 4122 5652 4140 5670
rect 4122 5670 4140 5688
rect 4122 5688 4140 5706
rect 4122 5706 4140 5724
rect 4122 5724 4140 5742
rect 4122 5742 4140 5760
rect 4122 5760 4140 5778
rect 4122 5778 4140 5796
rect 4122 5796 4140 5814
rect 4122 5814 4140 5832
rect 4122 5832 4140 5850
rect 4122 5850 4140 5868
rect 4122 5868 4140 5886
rect 4122 5886 4140 5904
rect 4122 5904 4140 5922
rect 4122 5922 4140 5940
rect 4122 5940 4140 5958
rect 4122 5958 4140 5976
rect 4122 5976 4140 5994
rect 4122 5994 4140 6012
rect 4122 6012 4140 6030
rect 4122 6030 4140 6048
rect 4122 6048 4140 6066
rect 4122 6066 4140 6084
rect 4122 6084 4140 6102
rect 4122 6102 4140 6120
rect 4122 6120 4140 6138
rect 4122 6138 4140 6156
rect 4122 6156 4140 6174
rect 4122 6174 4140 6192
rect 4122 6192 4140 6210
rect 4122 6210 4140 6228
rect 4122 6228 4140 6246
rect 4122 6246 4140 6264
rect 4122 6264 4140 6282
rect 4122 6282 4140 6300
rect 4122 6300 4140 6318
rect 4122 6318 4140 6336
rect 4122 6678 4140 6696
rect 4122 6696 4140 6714
rect 4122 6714 4140 6732
rect 4122 6732 4140 6750
rect 4122 6750 4140 6768
rect 4122 6768 4140 6786
rect 4122 6786 4140 6804
rect 4122 6804 4140 6822
rect 4122 6822 4140 6840
rect 4122 6840 4140 6858
rect 4122 6858 4140 6876
rect 4122 6876 4140 6894
rect 4122 6894 4140 6912
rect 4122 6912 4140 6930
rect 4122 6930 4140 6948
rect 4122 6948 4140 6966
rect 4122 6966 4140 6984
rect 4122 6984 4140 7002
rect 4122 7002 4140 7020
rect 4122 7020 4140 7038
rect 4122 7038 4140 7056
rect 4122 7056 4140 7074
rect 4122 7074 4140 7092
rect 4122 7092 4140 7110
rect 4122 7110 4140 7128
rect 4122 7128 4140 7146
rect 4122 7146 4140 7164
rect 4122 7164 4140 7182
rect 4122 7182 4140 7200
rect 4122 7200 4140 7218
rect 4122 7218 4140 7236
rect 4140 36 4158 54
rect 4140 54 4158 72
rect 4140 72 4158 90
rect 4140 90 4158 108
rect 4140 108 4158 126
rect 4140 126 4158 144
rect 4140 144 4158 162
rect 4140 162 4158 180
rect 4140 180 4158 198
rect 4140 198 4158 216
rect 4140 216 4158 234
rect 4140 234 4158 252
rect 4140 252 4158 270
rect 4140 270 4158 288
rect 4140 288 4158 306
rect 4140 306 4158 324
rect 4140 324 4158 342
rect 4140 342 4158 360
rect 4140 360 4158 378
rect 4140 378 4158 396
rect 4140 396 4158 414
rect 4140 414 4158 432
rect 4140 432 4158 450
rect 4140 450 4158 468
rect 4140 468 4158 486
rect 4140 486 4158 504
rect 4140 504 4158 522
rect 4140 522 4158 540
rect 4140 540 4158 558
rect 4140 558 4158 576
rect 4140 576 4158 594
rect 4140 594 4158 612
rect 4140 612 4158 630
rect 4140 630 4158 648
rect 4140 648 4158 666
rect 4140 864 4158 882
rect 4140 882 4158 900
rect 4140 900 4158 918
rect 4140 918 4158 936
rect 4140 936 4158 954
rect 4140 954 4158 972
rect 4140 972 4158 990
rect 4140 990 4158 1008
rect 4140 1008 4158 1026
rect 4140 1026 4158 1044
rect 4140 1044 4158 1062
rect 4140 1062 4158 1080
rect 4140 1080 4158 1098
rect 4140 1098 4158 1116
rect 4140 1116 4158 1134
rect 4140 1134 4158 1152
rect 4140 1152 4158 1170
rect 4140 1170 4158 1188
rect 4140 1188 4158 1206
rect 4140 1206 4158 1224
rect 4140 1224 4158 1242
rect 4140 1242 4158 1260
rect 4140 1260 4158 1278
rect 4140 1278 4158 1296
rect 4140 1296 4158 1314
rect 4140 1314 4158 1332
rect 4140 1332 4158 1350
rect 4140 1350 4158 1368
rect 4140 1368 4158 1386
rect 4140 1386 4158 1404
rect 4140 1404 4158 1422
rect 4140 1422 4158 1440
rect 4140 1440 4158 1458
rect 4140 1458 4158 1476
rect 4140 1476 4158 1494
rect 4140 1494 4158 1512
rect 4140 1512 4158 1530
rect 4140 1530 4158 1548
rect 4140 1548 4158 1566
rect 4140 1566 4158 1584
rect 4140 1584 4158 1602
rect 4140 1602 4158 1620
rect 4140 1620 4158 1638
rect 4140 1638 4158 1656
rect 4140 1908 4158 1926
rect 4140 1926 4158 1944
rect 4140 1944 4158 1962
rect 4140 1962 4158 1980
rect 4140 1980 4158 1998
rect 4140 1998 4158 2016
rect 4140 2016 4158 2034
rect 4140 2034 4158 2052
rect 4140 2052 4158 2070
rect 4140 2070 4158 2088
rect 4140 2088 4158 2106
rect 4140 2106 4158 2124
rect 4140 2124 4158 2142
rect 4140 2142 4158 2160
rect 4140 2160 4158 2178
rect 4140 2178 4158 2196
rect 4140 2196 4158 2214
rect 4140 2214 4158 2232
rect 4140 2232 4158 2250
rect 4140 2250 4158 2268
rect 4140 2268 4158 2286
rect 4140 2286 4158 2304
rect 4140 2304 4158 2322
rect 4140 2322 4158 2340
rect 4140 2340 4158 2358
rect 4140 2358 4158 2376
rect 4140 2376 4158 2394
rect 4140 2394 4158 2412
rect 4140 2412 4158 2430
rect 4140 2430 4158 2448
rect 4140 2448 4158 2466
rect 4140 2466 4158 2484
rect 4140 2484 4158 2502
rect 4140 2502 4158 2520
rect 4140 2520 4158 2538
rect 4140 2538 4158 2556
rect 4140 2556 4158 2574
rect 4140 2574 4158 2592
rect 4140 2592 4158 2610
rect 4140 2610 4158 2628
rect 4140 2628 4158 2646
rect 4140 2646 4158 2664
rect 4140 2664 4158 2682
rect 4140 2682 4158 2700
rect 4140 2700 4158 2718
rect 4140 2718 4158 2736
rect 4140 2736 4158 2754
rect 4140 2754 4158 2772
rect 4140 2772 4158 2790
rect 4140 2790 4158 2808
rect 4140 2808 4158 2826
rect 4140 2826 4158 2844
rect 4140 2844 4158 2862
rect 4140 2862 4158 2880
rect 4140 2880 4158 2898
rect 4140 2898 4158 2916
rect 4140 2916 4158 2934
rect 4140 2934 4158 2952
rect 4140 2952 4158 2970
rect 4140 2970 4158 2988
rect 4140 2988 4158 3006
rect 4140 3006 4158 3024
rect 4140 3024 4158 3042
rect 4140 3042 4158 3060
rect 4140 3060 4158 3078
rect 4140 3078 4158 3096
rect 4140 3096 4158 3114
rect 4140 3114 4158 3132
rect 4140 3132 4158 3150
rect 4140 3150 4158 3168
rect 4140 3168 4158 3186
rect 4140 3186 4158 3204
rect 4140 3204 4158 3222
rect 4140 3222 4158 3240
rect 4140 3240 4158 3258
rect 4140 3258 4158 3276
rect 4140 3276 4158 3294
rect 4140 3510 4158 3528
rect 4140 3528 4158 3546
rect 4140 3546 4158 3564
rect 4140 3564 4158 3582
rect 4140 3582 4158 3600
rect 4140 3600 4158 3618
rect 4140 3618 4158 3636
rect 4140 3636 4158 3654
rect 4140 3654 4158 3672
rect 4140 3672 4158 3690
rect 4140 3690 4158 3708
rect 4140 3708 4158 3726
rect 4140 3726 4158 3744
rect 4140 3744 4158 3762
rect 4140 3762 4158 3780
rect 4140 3780 4158 3798
rect 4140 3798 4158 3816
rect 4140 3816 4158 3834
rect 4140 3834 4158 3852
rect 4140 3852 4158 3870
rect 4140 3870 4158 3888
rect 4140 3888 4158 3906
rect 4140 3906 4158 3924
rect 4140 3924 4158 3942
rect 4140 3942 4158 3960
rect 4140 3960 4158 3978
rect 4140 3978 4158 3996
rect 4140 3996 4158 4014
rect 4140 4014 4158 4032
rect 4140 4032 4158 4050
rect 4140 4050 4158 4068
rect 4140 4068 4158 4086
rect 4140 4086 4158 4104
rect 4140 4104 4158 4122
rect 4140 4122 4158 4140
rect 4140 4140 4158 4158
rect 4140 4158 4158 4176
rect 4140 4176 4158 4194
rect 4140 4194 4158 4212
rect 4140 4212 4158 4230
rect 4140 4230 4158 4248
rect 4140 4248 4158 4266
rect 4140 4266 4158 4284
rect 4140 4284 4158 4302
rect 4140 4302 4158 4320
rect 4140 4320 4158 4338
rect 4140 4338 4158 4356
rect 4140 4356 4158 4374
rect 4140 4374 4158 4392
rect 4140 4392 4158 4410
rect 4140 4410 4158 4428
rect 4140 4428 4158 4446
rect 4140 4446 4158 4464
rect 4140 4464 4158 4482
rect 4140 4482 4158 4500
rect 4140 4500 4158 4518
rect 4140 4518 4158 4536
rect 4140 4536 4158 4554
rect 4140 4554 4158 4572
rect 4140 4572 4158 4590
rect 4140 4590 4158 4608
rect 4140 4608 4158 4626
rect 4140 4626 4158 4644
rect 4140 4644 4158 4662
rect 4140 4662 4158 4680
rect 4140 4680 4158 4698
rect 4140 4698 4158 4716
rect 4140 4716 4158 4734
rect 4140 4734 4158 4752
rect 4140 4752 4158 4770
rect 4140 4770 4158 4788
rect 4140 4788 4158 4806
rect 4140 4806 4158 4824
rect 4140 4824 4158 4842
rect 4140 4842 4158 4860
rect 4140 4860 4158 4878
rect 4140 4878 4158 4896
rect 4140 4896 4158 4914
rect 4140 4914 4158 4932
rect 4140 4932 4158 4950
rect 4140 4950 4158 4968
rect 4140 4968 4158 4986
rect 4140 4986 4158 5004
rect 4140 5004 4158 5022
rect 4140 5022 4158 5040
rect 4140 5040 4158 5058
rect 4140 5058 4158 5076
rect 4140 5076 4158 5094
rect 4140 5094 4158 5112
rect 4140 5112 4158 5130
rect 4140 5130 4158 5148
rect 4140 5148 4158 5166
rect 4140 5166 4158 5184
rect 4140 5184 4158 5202
rect 4140 5202 4158 5220
rect 4140 5220 4158 5238
rect 4140 5238 4158 5256
rect 4140 5256 4158 5274
rect 4140 5274 4158 5292
rect 4140 5292 4158 5310
rect 4140 5310 4158 5328
rect 4140 5328 4158 5346
rect 4140 5346 4158 5364
rect 4140 5364 4158 5382
rect 4140 5382 4158 5400
rect 4140 5400 4158 5418
rect 4140 5418 4158 5436
rect 4140 5436 4158 5454
rect 4140 5454 4158 5472
rect 4140 5472 4158 5490
rect 4140 5490 4158 5508
rect 4140 5508 4158 5526
rect 4140 5526 4158 5544
rect 4140 5544 4158 5562
rect 4140 5562 4158 5580
rect 4140 5580 4158 5598
rect 4140 5598 4158 5616
rect 4140 5616 4158 5634
rect 4140 5634 4158 5652
rect 4140 5652 4158 5670
rect 4140 5670 4158 5688
rect 4140 5688 4158 5706
rect 4140 5706 4158 5724
rect 4140 5724 4158 5742
rect 4140 5742 4158 5760
rect 4140 5760 4158 5778
rect 4140 5778 4158 5796
rect 4140 5796 4158 5814
rect 4140 5814 4158 5832
rect 4140 5832 4158 5850
rect 4140 5850 4158 5868
rect 4140 5868 4158 5886
rect 4140 5886 4158 5904
rect 4140 5904 4158 5922
rect 4140 5922 4158 5940
rect 4140 5940 4158 5958
rect 4140 5958 4158 5976
rect 4140 5976 4158 5994
rect 4140 5994 4158 6012
rect 4140 6012 4158 6030
rect 4140 6030 4158 6048
rect 4140 6048 4158 6066
rect 4140 6066 4158 6084
rect 4140 6084 4158 6102
rect 4140 6102 4158 6120
rect 4140 6120 4158 6138
rect 4140 6138 4158 6156
rect 4140 6156 4158 6174
rect 4140 6174 4158 6192
rect 4140 6192 4158 6210
rect 4140 6210 4158 6228
rect 4140 6228 4158 6246
rect 4140 6246 4158 6264
rect 4140 6264 4158 6282
rect 4140 6282 4158 6300
rect 4140 6300 4158 6318
rect 4140 6318 4158 6336
rect 4140 6336 4158 6354
rect 4140 6354 4158 6372
rect 4140 6714 4158 6732
rect 4140 6732 4158 6750
rect 4140 6750 4158 6768
rect 4140 6768 4158 6786
rect 4140 6786 4158 6804
rect 4140 6804 4158 6822
rect 4140 6822 4158 6840
rect 4140 6840 4158 6858
rect 4140 6858 4158 6876
rect 4140 6876 4158 6894
rect 4140 6894 4158 6912
rect 4140 6912 4158 6930
rect 4140 6930 4158 6948
rect 4140 6948 4158 6966
rect 4140 6966 4158 6984
rect 4140 6984 4158 7002
rect 4140 7002 4158 7020
rect 4140 7020 4158 7038
rect 4140 7038 4158 7056
rect 4140 7056 4158 7074
rect 4140 7074 4158 7092
rect 4140 7092 4158 7110
rect 4140 7110 4158 7128
rect 4140 7128 4158 7146
rect 4140 7146 4158 7164
rect 4140 7164 4158 7182
rect 4140 7182 4158 7200
rect 4140 7200 4158 7218
rect 4140 7218 4158 7236
rect 4158 36 4176 54
rect 4158 54 4176 72
rect 4158 72 4176 90
rect 4158 90 4176 108
rect 4158 108 4176 126
rect 4158 126 4176 144
rect 4158 144 4176 162
rect 4158 162 4176 180
rect 4158 180 4176 198
rect 4158 198 4176 216
rect 4158 216 4176 234
rect 4158 234 4176 252
rect 4158 252 4176 270
rect 4158 270 4176 288
rect 4158 288 4176 306
rect 4158 306 4176 324
rect 4158 324 4176 342
rect 4158 342 4176 360
rect 4158 360 4176 378
rect 4158 378 4176 396
rect 4158 396 4176 414
rect 4158 414 4176 432
rect 4158 432 4176 450
rect 4158 450 4176 468
rect 4158 468 4176 486
rect 4158 486 4176 504
rect 4158 504 4176 522
rect 4158 522 4176 540
rect 4158 540 4176 558
rect 4158 558 4176 576
rect 4158 576 4176 594
rect 4158 594 4176 612
rect 4158 612 4176 630
rect 4158 630 4176 648
rect 4158 648 4176 666
rect 4158 864 4176 882
rect 4158 882 4176 900
rect 4158 900 4176 918
rect 4158 918 4176 936
rect 4158 936 4176 954
rect 4158 954 4176 972
rect 4158 972 4176 990
rect 4158 990 4176 1008
rect 4158 1008 4176 1026
rect 4158 1026 4176 1044
rect 4158 1044 4176 1062
rect 4158 1062 4176 1080
rect 4158 1080 4176 1098
rect 4158 1098 4176 1116
rect 4158 1116 4176 1134
rect 4158 1134 4176 1152
rect 4158 1152 4176 1170
rect 4158 1170 4176 1188
rect 4158 1188 4176 1206
rect 4158 1206 4176 1224
rect 4158 1224 4176 1242
rect 4158 1242 4176 1260
rect 4158 1260 4176 1278
rect 4158 1278 4176 1296
rect 4158 1296 4176 1314
rect 4158 1314 4176 1332
rect 4158 1332 4176 1350
rect 4158 1350 4176 1368
rect 4158 1368 4176 1386
rect 4158 1386 4176 1404
rect 4158 1404 4176 1422
rect 4158 1422 4176 1440
rect 4158 1440 4176 1458
rect 4158 1458 4176 1476
rect 4158 1476 4176 1494
rect 4158 1494 4176 1512
rect 4158 1512 4176 1530
rect 4158 1530 4176 1548
rect 4158 1548 4176 1566
rect 4158 1566 4176 1584
rect 4158 1584 4176 1602
rect 4158 1602 4176 1620
rect 4158 1620 4176 1638
rect 4158 1638 4176 1656
rect 4158 1656 4176 1674
rect 4158 1908 4176 1926
rect 4158 1926 4176 1944
rect 4158 1944 4176 1962
rect 4158 1962 4176 1980
rect 4158 1980 4176 1998
rect 4158 1998 4176 2016
rect 4158 2016 4176 2034
rect 4158 2034 4176 2052
rect 4158 2052 4176 2070
rect 4158 2070 4176 2088
rect 4158 2088 4176 2106
rect 4158 2106 4176 2124
rect 4158 2124 4176 2142
rect 4158 2142 4176 2160
rect 4158 2160 4176 2178
rect 4158 2178 4176 2196
rect 4158 2196 4176 2214
rect 4158 2214 4176 2232
rect 4158 2232 4176 2250
rect 4158 2250 4176 2268
rect 4158 2268 4176 2286
rect 4158 2286 4176 2304
rect 4158 2304 4176 2322
rect 4158 2322 4176 2340
rect 4158 2340 4176 2358
rect 4158 2358 4176 2376
rect 4158 2376 4176 2394
rect 4158 2394 4176 2412
rect 4158 2412 4176 2430
rect 4158 2430 4176 2448
rect 4158 2448 4176 2466
rect 4158 2466 4176 2484
rect 4158 2484 4176 2502
rect 4158 2502 4176 2520
rect 4158 2520 4176 2538
rect 4158 2538 4176 2556
rect 4158 2556 4176 2574
rect 4158 2574 4176 2592
rect 4158 2592 4176 2610
rect 4158 2610 4176 2628
rect 4158 2628 4176 2646
rect 4158 2646 4176 2664
rect 4158 2664 4176 2682
rect 4158 2682 4176 2700
rect 4158 2700 4176 2718
rect 4158 2718 4176 2736
rect 4158 2736 4176 2754
rect 4158 2754 4176 2772
rect 4158 2772 4176 2790
rect 4158 2790 4176 2808
rect 4158 2808 4176 2826
rect 4158 2826 4176 2844
rect 4158 2844 4176 2862
rect 4158 2862 4176 2880
rect 4158 2880 4176 2898
rect 4158 2898 4176 2916
rect 4158 2916 4176 2934
rect 4158 2934 4176 2952
rect 4158 2952 4176 2970
rect 4158 2970 4176 2988
rect 4158 2988 4176 3006
rect 4158 3006 4176 3024
rect 4158 3024 4176 3042
rect 4158 3042 4176 3060
rect 4158 3060 4176 3078
rect 4158 3078 4176 3096
rect 4158 3096 4176 3114
rect 4158 3114 4176 3132
rect 4158 3132 4176 3150
rect 4158 3150 4176 3168
rect 4158 3168 4176 3186
rect 4158 3186 4176 3204
rect 4158 3204 4176 3222
rect 4158 3222 4176 3240
rect 4158 3240 4176 3258
rect 4158 3258 4176 3276
rect 4158 3276 4176 3294
rect 4158 3294 4176 3312
rect 4158 3312 4176 3330
rect 4158 3546 4176 3564
rect 4158 3564 4176 3582
rect 4158 3582 4176 3600
rect 4158 3600 4176 3618
rect 4158 3618 4176 3636
rect 4158 3636 4176 3654
rect 4158 3654 4176 3672
rect 4158 3672 4176 3690
rect 4158 3690 4176 3708
rect 4158 3708 4176 3726
rect 4158 3726 4176 3744
rect 4158 3744 4176 3762
rect 4158 3762 4176 3780
rect 4158 3780 4176 3798
rect 4158 3798 4176 3816
rect 4158 3816 4176 3834
rect 4158 3834 4176 3852
rect 4158 3852 4176 3870
rect 4158 3870 4176 3888
rect 4158 3888 4176 3906
rect 4158 3906 4176 3924
rect 4158 3924 4176 3942
rect 4158 3942 4176 3960
rect 4158 3960 4176 3978
rect 4158 3978 4176 3996
rect 4158 3996 4176 4014
rect 4158 4014 4176 4032
rect 4158 4032 4176 4050
rect 4158 4050 4176 4068
rect 4158 4068 4176 4086
rect 4158 4086 4176 4104
rect 4158 4104 4176 4122
rect 4158 4122 4176 4140
rect 4158 4140 4176 4158
rect 4158 4158 4176 4176
rect 4158 4176 4176 4194
rect 4158 4194 4176 4212
rect 4158 4212 4176 4230
rect 4158 4230 4176 4248
rect 4158 4248 4176 4266
rect 4158 4266 4176 4284
rect 4158 4284 4176 4302
rect 4158 4302 4176 4320
rect 4158 4320 4176 4338
rect 4158 4338 4176 4356
rect 4158 4356 4176 4374
rect 4158 4374 4176 4392
rect 4158 4392 4176 4410
rect 4158 4410 4176 4428
rect 4158 4428 4176 4446
rect 4158 4446 4176 4464
rect 4158 4464 4176 4482
rect 4158 4482 4176 4500
rect 4158 4500 4176 4518
rect 4158 4518 4176 4536
rect 4158 4536 4176 4554
rect 4158 4554 4176 4572
rect 4158 4572 4176 4590
rect 4158 4590 4176 4608
rect 4158 4608 4176 4626
rect 4158 4626 4176 4644
rect 4158 4644 4176 4662
rect 4158 4662 4176 4680
rect 4158 4680 4176 4698
rect 4158 4698 4176 4716
rect 4158 4716 4176 4734
rect 4158 4734 4176 4752
rect 4158 4752 4176 4770
rect 4158 4770 4176 4788
rect 4158 4788 4176 4806
rect 4158 4806 4176 4824
rect 4158 4824 4176 4842
rect 4158 4842 4176 4860
rect 4158 4860 4176 4878
rect 4158 4878 4176 4896
rect 4158 4896 4176 4914
rect 4158 4914 4176 4932
rect 4158 4932 4176 4950
rect 4158 4950 4176 4968
rect 4158 4968 4176 4986
rect 4158 4986 4176 5004
rect 4158 5004 4176 5022
rect 4158 5022 4176 5040
rect 4158 5040 4176 5058
rect 4158 5058 4176 5076
rect 4158 5076 4176 5094
rect 4158 5094 4176 5112
rect 4158 5112 4176 5130
rect 4158 5130 4176 5148
rect 4158 5148 4176 5166
rect 4158 5166 4176 5184
rect 4158 5184 4176 5202
rect 4158 5202 4176 5220
rect 4158 5220 4176 5238
rect 4158 5238 4176 5256
rect 4158 5256 4176 5274
rect 4158 5274 4176 5292
rect 4158 5292 4176 5310
rect 4158 5310 4176 5328
rect 4158 5328 4176 5346
rect 4158 5346 4176 5364
rect 4158 5364 4176 5382
rect 4158 5382 4176 5400
rect 4158 5400 4176 5418
rect 4158 5418 4176 5436
rect 4158 5436 4176 5454
rect 4158 5454 4176 5472
rect 4158 5472 4176 5490
rect 4158 5490 4176 5508
rect 4158 5508 4176 5526
rect 4158 5526 4176 5544
rect 4158 5544 4176 5562
rect 4158 5562 4176 5580
rect 4158 5580 4176 5598
rect 4158 5598 4176 5616
rect 4158 5616 4176 5634
rect 4158 5634 4176 5652
rect 4158 5652 4176 5670
rect 4158 5670 4176 5688
rect 4158 5688 4176 5706
rect 4158 5706 4176 5724
rect 4158 5724 4176 5742
rect 4158 5742 4176 5760
rect 4158 5760 4176 5778
rect 4158 5778 4176 5796
rect 4158 5796 4176 5814
rect 4158 5814 4176 5832
rect 4158 5832 4176 5850
rect 4158 5850 4176 5868
rect 4158 5868 4176 5886
rect 4158 5886 4176 5904
rect 4158 5904 4176 5922
rect 4158 5922 4176 5940
rect 4158 5940 4176 5958
rect 4158 5958 4176 5976
rect 4158 5976 4176 5994
rect 4158 5994 4176 6012
rect 4158 6012 4176 6030
rect 4158 6030 4176 6048
rect 4158 6048 4176 6066
rect 4158 6066 4176 6084
rect 4158 6084 4176 6102
rect 4158 6102 4176 6120
rect 4158 6120 4176 6138
rect 4158 6138 4176 6156
rect 4158 6156 4176 6174
rect 4158 6174 4176 6192
rect 4158 6192 4176 6210
rect 4158 6210 4176 6228
rect 4158 6228 4176 6246
rect 4158 6246 4176 6264
rect 4158 6264 4176 6282
rect 4158 6282 4176 6300
rect 4158 6300 4176 6318
rect 4158 6318 4176 6336
rect 4158 6336 4176 6354
rect 4158 6354 4176 6372
rect 4158 6372 4176 6390
rect 4158 6390 4176 6408
rect 4158 6750 4176 6768
rect 4158 6768 4176 6786
rect 4158 6786 4176 6804
rect 4158 6804 4176 6822
rect 4158 6822 4176 6840
rect 4158 6840 4176 6858
rect 4158 6858 4176 6876
rect 4158 6876 4176 6894
rect 4158 6894 4176 6912
rect 4158 6912 4176 6930
rect 4158 6930 4176 6948
rect 4158 6948 4176 6966
rect 4158 6966 4176 6984
rect 4158 6984 4176 7002
rect 4158 7002 4176 7020
rect 4158 7020 4176 7038
rect 4158 7038 4176 7056
rect 4158 7056 4176 7074
rect 4158 7074 4176 7092
rect 4158 7092 4176 7110
rect 4158 7110 4176 7128
rect 4158 7128 4176 7146
rect 4158 7146 4176 7164
rect 4158 7164 4176 7182
rect 4158 7182 4176 7200
rect 4158 7200 4176 7218
rect 4158 7218 4176 7236
rect 4176 36 4194 54
rect 4176 54 4194 72
rect 4176 72 4194 90
rect 4176 90 4194 108
rect 4176 108 4194 126
rect 4176 126 4194 144
rect 4176 144 4194 162
rect 4176 162 4194 180
rect 4176 180 4194 198
rect 4176 198 4194 216
rect 4176 216 4194 234
rect 4176 234 4194 252
rect 4176 252 4194 270
rect 4176 270 4194 288
rect 4176 288 4194 306
rect 4176 306 4194 324
rect 4176 324 4194 342
rect 4176 342 4194 360
rect 4176 360 4194 378
rect 4176 378 4194 396
rect 4176 396 4194 414
rect 4176 414 4194 432
rect 4176 432 4194 450
rect 4176 450 4194 468
rect 4176 468 4194 486
rect 4176 486 4194 504
rect 4176 504 4194 522
rect 4176 522 4194 540
rect 4176 540 4194 558
rect 4176 558 4194 576
rect 4176 576 4194 594
rect 4176 594 4194 612
rect 4176 612 4194 630
rect 4176 630 4194 648
rect 4176 648 4194 666
rect 4176 864 4194 882
rect 4176 882 4194 900
rect 4176 900 4194 918
rect 4176 918 4194 936
rect 4176 936 4194 954
rect 4176 954 4194 972
rect 4176 972 4194 990
rect 4176 990 4194 1008
rect 4176 1008 4194 1026
rect 4176 1026 4194 1044
rect 4176 1044 4194 1062
rect 4176 1062 4194 1080
rect 4176 1080 4194 1098
rect 4176 1098 4194 1116
rect 4176 1116 4194 1134
rect 4176 1134 4194 1152
rect 4176 1152 4194 1170
rect 4176 1170 4194 1188
rect 4176 1188 4194 1206
rect 4176 1206 4194 1224
rect 4176 1224 4194 1242
rect 4176 1242 4194 1260
rect 4176 1260 4194 1278
rect 4176 1278 4194 1296
rect 4176 1296 4194 1314
rect 4176 1314 4194 1332
rect 4176 1332 4194 1350
rect 4176 1350 4194 1368
rect 4176 1368 4194 1386
rect 4176 1386 4194 1404
rect 4176 1404 4194 1422
rect 4176 1422 4194 1440
rect 4176 1440 4194 1458
rect 4176 1458 4194 1476
rect 4176 1476 4194 1494
rect 4176 1494 4194 1512
rect 4176 1512 4194 1530
rect 4176 1530 4194 1548
rect 4176 1548 4194 1566
rect 4176 1566 4194 1584
rect 4176 1584 4194 1602
rect 4176 1602 4194 1620
rect 4176 1620 4194 1638
rect 4176 1638 4194 1656
rect 4176 1656 4194 1674
rect 4176 1674 4194 1692
rect 4176 1926 4194 1944
rect 4176 1944 4194 1962
rect 4176 1962 4194 1980
rect 4176 1980 4194 1998
rect 4176 1998 4194 2016
rect 4176 2016 4194 2034
rect 4176 2034 4194 2052
rect 4176 2052 4194 2070
rect 4176 2070 4194 2088
rect 4176 2088 4194 2106
rect 4176 2106 4194 2124
rect 4176 2124 4194 2142
rect 4176 2142 4194 2160
rect 4176 2160 4194 2178
rect 4176 2178 4194 2196
rect 4176 2196 4194 2214
rect 4176 2214 4194 2232
rect 4176 2232 4194 2250
rect 4176 2250 4194 2268
rect 4176 2268 4194 2286
rect 4176 2286 4194 2304
rect 4176 2304 4194 2322
rect 4176 2322 4194 2340
rect 4176 2340 4194 2358
rect 4176 2358 4194 2376
rect 4176 2376 4194 2394
rect 4176 2394 4194 2412
rect 4176 2412 4194 2430
rect 4176 2430 4194 2448
rect 4176 2448 4194 2466
rect 4176 2466 4194 2484
rect 4176 2484 4194 2502
rect 4176 2502 4194 2520
rect 4176 2520 4194 2538
rect 4176 2538 4194 2556
rect 4176 2556 4194 2574
rect 4176 2574 4194 2592
rect 4176 2592 4194 2610
rect 4176 2610 4194 2628
rect 4176 2628 4194 2646
rect 4176 2646 4194 2664
rect 4176 2664 4194 2682
rect 4176 2682 4194 2700
rect 4176 2700 4194 2718
rect 4176 2718 4194 2736
rect 4176 2736 4194 2754
rect 4176 2754 4194 2772
rect 4176 2772 4194 2790
rect 4176 2790 4194 2808
rect 4176 2808 4194 2826
rect 4176 2826 4194 2844
rect 4176 2844 4194 2862
rect 4176 2862 4194 2880
rect 4176 2880 4194 2898
rect 4176 2898 4194 2916
rect 4176 2916 4194 2934
rect 4176 2934 4194 2952
rect 4176 2952 4194 2970
rect 4176 2970 4194 2988
rect 4176 2988 4194 3006
rect 4176 3006 4194 3024
rect 4176 3024 4194 3042
rect 4176 3042 4194 3060
rect 4176 3060 4194 3078
rect 4176 3078 4194 3096
rect 4176 3096 4194 3114
rect 4176 3114 4194 3132
rect 4176 3132 4194 3150
rect 4176 3150 4194 3168
rect 4176 3168 4194 3186
rect 4176 3186 4194 3204
rect 4176 3204 4194 3222
rect 4176 3222 4194 3240
rect 4176 3240 4194 3258
rect 4176 3258 4194 3276
rect 4176 3276 4194 3294
rect 4176 3294 4194 3312
rect 4176 3312 4194 3330
rect 4176 3330 4194 3348
rect 4176 3564 4194 3582
rect 4176 3582 4194 3600
rect 4176 3600 4194 3618
rect 4176 3618 4194 3636
rect 4176 3636 4194 3654
rect 4176 3654 4194 3672
rect 4176 3672 4194 3690
rect 4176 3690 4194 3708
rect 4176 3708 4194 3726
rect 4176 3726 4194 3744
rect 4176 3744 4194 3762
rect 4176 3762 4194 3780
rect 4176 3780 4194 3798
rect 4176 3798 4194 3816
rect 4176 3816 4194 3834
rect 4176 3834 4194 3852
rect 4176 3852 4194 3870
rect 4176 3870 4194 3888
rect 4176 3888 4194 3906
rect 4176 3906 4194 3924
rect 4176 3924 4194 3942
rect 4176 3942 4194 3960
rect 4176 3960 4194 3978
rect 4176 3978 4194 3996
rect 4176 3996 4194 4014
rect 4176 4014 4194 4032
rect 4176 4032 4194 4050
rect 4176 4050 4194 4068
rect 4176 4068 4194 4086
rect 4176 4086 4194 4104
rect 4176 4104 4194 4122
rect 4176 4122 4194 4140
rect 4176 4140 4194 4158
rect 4176 4158 4194 4176
rect 4176 4176 4194 4194
rect 4176 4194 4194 4212
rect 4176 4212 4194 4230
rect 4176 4230 4194 4248
rect 4176 4248 4194 4266
rect 4176 4266 4194 4284
rect 4176 4284 4194 4302
rect 4176 4302 4194 4320
rect 4176 4320 4194 4338
rect 4176 4338 4194 4356
rect 4176 4356 4194 4374
rect 4176 4374 4194 4392
rect 4176 4392 4194 4410
rect 4176 4410 4194 4428
rect 4176 4428 4194 4446
rect 4176 4446 4194 4464
rect 4176 4464 4194 4482
rect 4176 4482 4194 4500
rect 4176 4500 4194 4518
rect 4176 4518 4194 4536
rect 4176 4536 4194 4554
rect 4176 4554 4194 4572
rect 4176 4572 4194 4590
rect 4176 4590 4194 4608
rect 4176 4608 4194 4626
rect 4176 4626 4194 4644
rect 4176 4644 4194 4662
rect 4176 4662 4194 4680
rect 4176 4680 4194 4698
rect 4176 4698 4194 4716
rect 4176 4716 4194 4734
rect 4176 4734 4194 4752
rect 4176 4752 4194 4770
rect 4176 4770 4194 4788
rect 4176 4788 4194 4806
rect 4176 4806 4194 4824
rect 4176 4824 4194 4842
rect 4176 4842 4194 4860
rect 4176 4860 4194 4878
rect 4176 4878 4194 4896
rect 4176 4896 4194 4914
rect 4176 4914 4194 4932
rect 4176 4932 4194 4950
rect 4176 4950 4194 4968
rect 4176 4968 4194 4986
rect 4176 4986 4194 5004
rect 4176 5004 4194 5022
rect 4176 5022 4194 5040
rect 4176 5040 4194 5058
rect 4176 5058 4194 5076
rect 4176 5076 4194 5094
rect 4176 5094 4194 5112
rect 4176 5112 4194 5130
rect 4176 5130 4194 5148
rect 4176 5148 4194 5166
rect 4176 5166 4194 5184
rect 4176 5184 4194 5202
rect 4176 5202 4194 5220
rect 4176 5220 4194 5238
rect 4176 5238 4194 5256
rect 4176 5256 4194 5274
rect 4176 5274 4194 5292
rect 4176 5292 4194 5310
rect 4176 5310 4194 5328
rect 4176 5328 4194 5346
rect 4176 5346 4194 5364
rect 4176 5364 4194 5382
rect 4176 5382 4194 5400
rect 4176 5400 4194 5418
rect 4176 5418 4194 5436
rect 4176 5436 4194 5454
rect 4176 5454 4194 5472
rect 4176 5472 4194 5490
rect 4176 5490 4194 5508
rect 4176 5508 4194 5526
rect 4176 5526 4194 5544
rect 4176 5544 4194 5562
rect 4176 5562 4194 5580
rect 4176 5580 4194 5598
rect 4176 5598 4194 5616
rect 4176 5616 4194 5634
rect 4176 5634 4194 5652
rect 4176 5652 4194 5670
rect 4176 5670 4194 5688
rect 4176 5688 4194 5706
rect 4176 5706 4194 5724
rect 4176 5724 4194 5742
rect 4176 5742 4194 5760
rect 4176 5760 4194 5778
rect 4176 5778 4194 5796
rect 4176 5796 4194 5814
rect 4176 5814 4194 5832
rect 4176 5832 4194 5850
rect 4176 5850 4194 5868
rect 4176 5868 4194 5886
rect 4176 5886 4194 5904
rect 4176 5904 4194 5922
rect 4176 5922 4194 5940
rect 4176 5940 4194 5958
rect 4176 5958 4194 5976
rect 4176 5976 4194 5994
rect 4176 5994 4194 6012
rect 4176 6012 4194 6030
rect 4176 6030 4194 6048
rect 4176 6048 4194 6066
rect 4176 6066 4194 6084
rect 4176 6084 4194 6102
rect 4176 6102 4194 6120
rect 4176 6120 4194 6138
rect 4176 6138 4194 6156
rect 4176 6156 4194 6174
rect 4176 6174 4194 6192
rect 4176 6192 4194 6210
rect 4176 6210 4194 6228
rect 4176 6228 4194 6246
rect 4176 6246 4194 6264
rect 4176 6264 4194 6282
rect 4176 6282 4194 6300
rect 4176 6300 4194 6318
rect 4176 6318 4194 6336
rect 4176 6336 4194 6354
rect 4176 6354 4194 6372
rect 4176 6372 4194 6390
rect 4176 6390 4194 6408
rect 4176 6408 4194 6426
rect 4176 6426 4194 6444
rect 4176 6786 4194 6804
rect 4176 6804 4194 6822
rect 4176 6822 4194 6840
rect 4176 6840 4194 6858
rect 4176 6858 4194 6876
rect 4176 6876 4194 6894
rect 4176 6894 4194 6912
rect 4176 6912 4194 6930
rect 4176 6930 4194 6948
rect 4176 6948 4194 6966
rect 4176 6966 4194 6984
rect 4176 6984 4194 7002
rect 4176 7002 4194 7020
rect 4176 7020 4194 7038
rect 4176 7038 4194 7056
rect 4176 7056 4194 7074
rect 4176 7074 4194 7092
rect 4176 7092 4194 7110
rect 4176 7110 4194 7128
rect 4176 7128 4194 7146
rect 4176 7146 4194 7164
rect 4176 7164 4194 7182
rect 4176 7182 4194 7200
rect 4176 7200 4194 7218
rect 4176 7218 4194 7236
rect 4194 36 4212 54
rect 4194 54 4212 72
rect 4194 72 4212 90
rect 4194 90 4212 108
rect 4194 108 4212 126
rect 4194 126 4212 144
rect 4194 144 4212 162
rect 4194 162 4212 180
rect 4194 180 4212 198
rect 4194 198 4212 216
rect 4194 216 4212 234
rect 4194 234 4212 252
rect 4194 252 4212 270
rect 4194 270 4212 288
rect 4194 288 4212 306
rect 4194 306 4212 324
rect 4194 324 4212 342
rect 4194 342 4212 360
rect 4194 360 4212 378
rect 4194 378 4212 396
rect 4194 396 4212 414
rect 4194 414 4212 432
rect 4194 432 4212 450
rect 4194 450 4212 468
rect 4194 468 4212 486
rect 4194 486 4212 504
rect 4194 504 4212 522
rect 4194 522 4212 540
rect 4194 540 4212 558
rect 4194 558 4212 576
rect 4194 576 4212 594
rect 4194 594 4212 612
rect 4194 612 4212 630
rect 4194 630 4212 648
rect 4194 648 4212 666
rect 4194 864 4212 882
rect 4194 882 4212 900
rect 4194 900 4212 918
rect 4194 918 4212 936
rect 4194 936 4212 954
rect 4194 954 4212 972
rect 4194 972 4212 990
rect 4194 990 4212 1008
rect 4194 1008 4212 1026
rect 4194 1026 4212 1044
rect 4194 1044 4212 1062
rect 4194 1062 4212 1080
rect 4194 1080 4212 1098
rect 4194 1098 4212 1116
rect 4194 1116 4212 1134
rect 4194 1134 4212 1152
rect 4194 1152 4212 1170
rect 4194 1170 4212 1188
rect 4194 1188 4212 1206
rect 4194 1206 4212 1224
rect 4194 1224 4212 1242
rect 4194 1242 4212 1260
rect 4194 1260 4212 1278
rect 4194 1278 4212 1296
rect 4194 1296 4212 1314
rect 4194 1314 4212 1332
rect 4194 1332 4212 1350
rect 4194 1350 4212 1368
rect 4194 1368 4212 1386
rect 4194 1386 4212 1404
rect 4194 1404 4212 1422
rect 4194 1422 4212 1440
rect 4194 1440 4212 1458
rect 4194 1458 4212 1476
rect 4194 1476 4212 1494
rect 4194 1494 4212 1512
rect 4194 1512 4212 1530
rect 4194 1530 4212 1548
rect 4194 1548 4212 1566
rect 4194 1566 4212 1584
rect 4194 1584 4212 1602
rect 4194 1602 4212 1620
rect 4194 1620 4212 1638
rect 4194 1638 4212 1656
rect 4194 1656 4212 1674
rect 4194 1674 4212 1692
rect 4194 1944 4212 1962
rect 4194 1962 4212 1980
rect 4194 1980 4212 1998
rect 4194 1998 4212 2016
rect 4194 2016 4212 2034
rect 4194 2034 4212 2052
rect 4194 2052 4212 2070
rect 4194 2070 4212 2088
rect 4194 2088 4212 2106
rect 4194 2106 4212 2124
rect 4194 2124 4212 2142
rect 4194 2142 4212 2160
rect 4194 2160 4212 2178
rect 4194 2178 4212 2196
rect 4194 2196 4212 2214
rect 4194 2214 4212 2232
rect 4194 2232 4212 2250
rect 4194 2250 4212 2268
rect 4194 2268 4212 2286
rect 4194 2286 4212 2304
rect 4194 2304 4212 2322
rect 4194 2322 4212 2340
rect 4194 2340 4212 2358
rect 4194 2358 4212 2376
rect 4194 2376 4212 2394
rect 4194 2394 4212 2412
rect 4194 2412 4212 2430
rect 4194 2430 4212 2448
rect 4194 2448 4212 2466
rect 4194 2466 4212 2484
rect 4194 2484 4212 2502
rect 4194 2502 4212 2520
rect 4194 2520 4212 2538
rect 4194 2538 4212 2556
rect 4194 2556 4212 2574
rect 4194 2574 4212 2592
rect 4194 2592 4212 2610
rect 4194 2610 4212 2628
rect 4194 2628 4212 2646
rect 4194 2646 4212 2664
rect 4194 2664 4212 2682
rect 4194 2682 4212 2700
rect 4194 2700 4212 2718
rect 4194 2718 4212 2736
rect 4194 2736 4212 2754
rect 4194 2754 4212 2772
rect 4194 2772 4212 2790
rect 4194 2790 4212 2808
rect 4194 2808 4212 2826
rect 4194 2826 4212 2844
rect 4194 2844 4212 2862
rect 4194 2862 4212 2880
rect 4194 2880 4212 2898
rect 4194 2898 4212 2916
rect 4194 2916 4212 2934
rect 4194 2934 4212 2952
rect 4194 2952 4212 2970
rect 4194 2970 4212 2988
rect 4194 2988 4212 3006
rect 4194 3006 4212 3024
rect 4194 3024 4212 3042
rect 4194 3042 4212 3060
rect 4194 3060 4212 3078
rect 4194 3078 4212 3096
rect 4194 3096 4212 3114
rect 4194 3114 4212 3132
rect 4194 3132 4212 3150
rect 4194 3150 4212 3168
rect 4194 3168 4212 3186
rect 4194 3186 4212 3204
rect 4194 3204 4212 3222
rect 4194 3222 4212 3240
rect 4194 3240 4212 3258
rect 4194 3258 4212 3276
rect 4194 3276 4212 3294
rect 4194 3294 4212 3312
rect 4194 3312 4212 3330
rect 4194 3330 4212 3348
rect 4194 3348 4212 3366
rect 4194 3366 4212 3384
rect 4194 3600 4212 3618
rect 4194 3618 4212 3636
rect 4194 3636 4212 3654
rect 4194 3654 4212 3672
rect 4194 3672 4212 3690
rect 4194 3690 4212 3708
rect 4194 3708 4212 3726
rect 4194 3726 4212 3744
rect 4194 3744 4212 3762
rect 4194 3762 4212 3780
rect 4194 3780 4212 3798
rect 4194 3798 4212 3816
rect 4194 3816 4212 3834
rect 4194 3834 4212 3852
rect 4194 3852 4212 3870
rect 4194 3870 4212 3888
rect 4194 3888 4212 3906
rect 4194 3906 4212 3924
rect 4194 3924 4212 3942
rect 4194 3942 4212 3960
rect 4194 3960 4212 3978
rect 4194 3978 4212 3996
rect 4194 3996 4212 4014
rect 4194 4014 4212 4032
rect 4194 4032 4212 4050
rect 4194 4050 4212 4068
rect 4194 4068 4212 4086
rect 4194 4086 4212 4104
rect 4194 4104 4212 4122
rect 4194 4122 4212 4140
rect 4194 4140 4212 4158
rect 4194 4158 4212 4176
rect 4194 4176 4212 4194
rect 4194 4194 4212 4212
rect 4194 4212 4212 4230
rect 4194 4230 4212 4248
rect 4194 4248 4212 4266
rect 4194 4266 4212 4284
rect 4194 4284 4212 4302
rect 4194 4302 4212 4320
rect 4194 4320 4212 4338
rect 4194 4338 4212 4356
rect 4194 4356 4212 4374
rect 4194 4374 4212 4392
rect 4194 4392 4212 4410
rect 4194 4410 4212 4428
rect 4194 4428 4212 4446
rect 4194 4446 4212 4464
rect 4194 4464 4212 4482
rect 4194 4482 4212 4500
rect 4194 4500 4212 4518
rect 4194 4518 4212 4536
rect 4194 4536 4212 4554
rect 4194 4554 4212 4572
rect 4194 4572 4212 4590
rect 4194 4590 4212 4608
rect 4194 4608 4212 4626
rect 4194 4626 4212 4644
rect 4194 4644 4212 4662
rect 4194 4662 4212 4680
rect 4194 4680 4212 4698
rect 4194 4698 4212 4716
rect 4194 4716 4212 4734
rect 4194 4734 4212 4752
rect 4194 4752 4212 4770
rect 4194 4770 4212 4788
rect 4194 4788 4212 4806
rect 4194 4806 4212 4824
rect 4194 4824 4212 4842
rect 4194 4842 4212 4860
rect 4194 4860 4212 4878
rect 4194 4878 4212 4896
rect 4194 4896 4212 4914
rect 4194 4914 4212 4932
rect 4194 4932 4212 4950
rect 4194 4950 4212 4968
rect 4194 4968 4212 4986
rect 4194 4986 4212 5004
rect 4194 5004 4212 5022
rect 4194 5022 4212 5040
rect 4194 5040 4212 5058
rect 4194 5058 4212 5076
rect 4194 5076 4212 5094
rect 4194 5094 4212 5112
rect 4194 5112 4212 5130
rect 4194 5130 4212 5148
rect 4194 5148 4212 5166
rect 4194 5166 4212 5184
rect 4194 5184 4212 5202
rect 4194 5202 4212 5220
rect 4194 5220 4212 5238
rect 4194 5238 4212 5256
rect 4194 5256 4212 5274
rect 4194 5274 4212 5292
rect 4194 5292 4212 5310
rect 4194 5310 4212 5328
rect 4194 5328 4212 5346
rect 4194 5346 4212 5364
rect 4194 5364 4212 5382
rect 4194 5382 4212 5400
rect 4194 5400 4212 5418
rect 4194 5418 4212 5436
rect 4194 5436 4212 5454
rect 4194 5454 4212 5472
rect 4194 5472 4212 5490
rect 4194 5490 4212 5508
rect 4194 5508 4212 5526
rect 4194 5526 4212 5544
rect 4194 5544 4212 5562
rect 4194 5562 4212 5580
rect 4194 5580 4212 5598
rect 4194 5598 4212 5616
rect 4194 5616 4212 5634
rect 4194 5634 4212 5652
rect 4194 5652 4212 5670
rect 4194 5670 4212 5688
rect 4194 5688 4212 5706
rect 4194 5706 4212 5724
rect 4194 5724 4212 5742
rect 4194 5742 4212 5760
rect 4194 5760 4212 5778
rect 4194 5778 4212 5796
rect 4194 5796 4212 5814
rect 4194 5814 4212 5832
rect 4194 5832 4212 5850
rect 4194 5850 4212 5868
rect 4194 5868 4212 5886
rect 4194 5886 4212 5904
rect 4194 5904 4212 5922
rect 4194 5922 4212 5940
rect 4194 5940 4212 5958
rect 4194 5958 4212 5976
rect 4194 5976 4212 5994
rect 4194 5994 4212 6012
rect 4194 6012 4212 6030
rect 4194 6030 4212 6048
rect 4194 6048 4212 6066
rect 4194 6066 4212 6084
rect 4194 6084 4212 6102
rect 4194 6102 4212 6120
rect 4194 6120 4212 6138
rect 4194 6138 4212 6156
rect 4194 6156 4212 6174
rect 4194 6174 4212 6192
rect 4194 6192 4212 6210
rect 4194 6210 4212 6228
rect 4194 6228 4212 6246
rect 4194 6246 4212 6264
rect 4194 6264 4212 6282
rect 4194 6282 4212 6300
rect 4194 6300 4212 6318
rect 4194 6318 4212 6336
rect 4194 6336 4212 6354
rect 4194 6354 4212 6372
rect 4194 6372 4212 6390
rect 4194 6390 4212 6408
rect 4194 6408 4212 6426
rect 4194 6426 4212 6444
rect 4194 6444 4212 6462
rect 4194 6462 4212 6480
rect 4194 6822 4212 6840
rect 4194 6840 4212 6858
rect 4194 6858 4212 6876
rect 4194 6876 4212 6894
rect 4194 6894 4212 6912
rect 4194 6912 4212 6930
rect 4194 6930 4212 6948
rect 4194 6948 4212 6966
rect 4194 6966 4212 6984
rect 4194 6984 4212 7002
rect 4194 7002 4212 7020
rect 4194 7020 4212 7038
rect 4194 7038 4212 7056
rect 4194 7056 4212 7074
rect 4194 7074 4212 7092
rect 4194 7092 4212 7110
rect 4194 7110 4212 7128
rect 4194 7128 4212 7146
rect 4194 7146 4212 7164
rect 4194 7164 4212 7182
rect 4194 7182 4212 7200
rect 4194 7200 4212 7218
rect 4194 7218 4212 7236
rect 4212 36 4230 54
rect 4212 54 4230 72
rect 4212 72 4230 90
rect 4212 90 4230 108
rect 4212 108 4230 126
rect 4212 126 4230 144
rect 4212 144 4230 162
rect 4212 162 4230 180
rect 4212 180 4230 198
rect 4212 198 4230 216
rect 4212 216 4230 234
rect 4212 234 4230 252
rect 4212 252 4230 270
rect 4212 270 4230 288
rect 4212 288 4230 306
rect 4212 306 4230 324
rect 4212 324 4230 342
rect 4212 342 4230 360
rect 4212 360 4230 378
rect 4212 378 4230 396
rect 4212 396 4230 414
rect 4212 414 4230 432
rect 4212 432 4230 450
rect 4212 450 4230 468
rect 4212 468 4230 486
rect 4212 486 4230 504
rect 4212 504 4230 522
rect 4212 522 4230 540
rect 4212 540 4230 558
rect 4212 558 4230 576
rect 4212 576 4230 594
rect 4212 594 4230 612
rect 4212 612 4230 630
rect 4212 630 4230 648
rect 4212 648 4230 666
rect 4212 864 4230 882
rect 4212 882 4230 900
rect 4212 900 4230 918
rect 4212 918 4230 936
rect 4212 936 4230 954
rect 4212 954 4230 972
rect 4212 972 4230 990
rect 4212 990 4230 1008
rect 4212 1008 4230 1026
rect 4212 1026 4230 1044
rect 4212 1044 4230 1062
rect 4212 1062 4230 1080
rect 4212 1080 4230 1098
rect 4212 1098 4230 1116
rect 4212 1116 4230 1134
rect 4212 1134 4230 1152
rect 4212 1152 4230 1170
rect 4212 1170 4230 1188
rect 4212 1188 4230 1206
rect 4212 1206 4230 1224
rect 4212 1224 4230 1242
rect 4212 1242 4230 1260
rect 4212 1260 4230 1278
rect 4212 1278 4230 1296
rect 4212 1296 4230 1314
rect 4212 1314 4230 1332
rect 4212 1332 4230 1350
rect 4212 1350 4230 1368
rect 4212 1368 4230 1386
rect 4212 1386 4230 1404
rect 4212 1404 4230 1422
rect 4212 1422 4230 1440
rect 4212 1440 4230 1458
rect 4212 1458 4230 1476
rect 4212 1476 4230 1494
rect 4212 1494 4230 1512
rect 4212 1512 4230 1530
rect 4212 1530 4230 1548
rect 4212 1548 4230 1566
rect 4212 1566 4230 1584
rect 4212 1584 4230 1602
rect 4212 1602 4230 1620
rect 4212 1620 4230 1638
rect 4212 1638 4230 1656
rect 4212 1656 4230 1674
rect 4212 1674 4230 1692
rect 4212 1692 4230 1710
rect 4212 1944 4230 1962
rect 4212 1962 4230 1980
rect 4212 1980 4230 1998
rect 4212 1998 4230 2016
rect 4212 2016 4230 2034
rect 4212 2034 4230 2052
rect 4212 2052 4230 2070
rect 4212 2070 4230 2088
rect 4212 2088 4230 2106
rect 4212 2106 4230 2124
rect 4212 2124 4230 2142
rect 4212 2142 4230 2160
rect 4212 2160 4230 2178
rect 4212 2178 4230 2196
rect 4212 2196 4230 2214
rect 4212 2214 4230 2232
rect 4212 2232 4230 2250
rect 4212 2250 4230 2268
rect 4212 2268 4230 2286
rect 4212 2286 4230 2304
rect 4212 2304 4230 2322
rect 4212 2322 4230 2340
rect 4212 2340 4230 2358
rect 4212 2358 4230 2376
rect 4212 2376 4230 2394
rect 4212 2394 4230 2412
rect 4212 2412 4230 2430
rect 4212 2430 4230 2448
rect 4212 2448 4230 2466
rect 4212 2466 4230 2484
rect 4212 2484 4230 2502
rect 4212 2502 4230 2520
rect 4212 2520 4230 2538
rect 4212 2538 4230 2556
rect 4212 2556 4230 2574
rect 4212 2574 4230 2592
rect 4212 2592 4230 2610
rect 4212 2610 4230 2628
rect 4212 2628 4230 2646
rect 4212 2646 4230 2664
rect 4212 2664 4230 2682
rect 4212 2682 4230 2700
rect 4212 2700 4230 2718
rect 4212 2718 4230 2736
rect 4212 2736 4230 2754
rect 4212 2754 4230 2772
rect 4212 2772 4230 2790
rect 4212 2790 4230 2808
rect 4212 2808 4230 2826
rect 4212 2826 4230 2844
rect 4212 2844 4230 2862
rect 4212 2862 4230 2880
rect 4212 2880 4230 2898
rect 4212 2898 4230 2916
rect 4212 2916 4230 2934
rect 4212 2934 4230 2952
rect 4212 2952 4230 2970
rect 4212 2970 4230 2988
rect 4212 2988 4230 3006
rect 4212 3006 4230 3024
rect 4212 3024 4230 3042
rect 4212 3042 4230 3060
rect 4212 3060 4230 3078
rect 4212 3078 4230 3096
rect 4212 3096 4230 3114
rect 4212 3114 4230 3132
rect 4212 3132 4230 3150
rect 4212 3150 4230 3168
rect 4212 3168 4230 3186
rect 4212 3186 4230 3204
rect 4212 3204 4230 3222
rect 4212 3222 4230 3240
rect 4212 3240 4230 3258
rect 4212 3258 4230 3276
rect 4212 3276 4230 3294
rect 4212 3294 4230 3312
rect 4212 3312 4230 3330
rect 4212 3330 4230 3348
rect 4212 3348 4230 3366
rect 4212 3366 4230 3384
rect 4212 3384 4230 3402
rect 4212 3618 4230 3636
rect 4212 3636 4230 3654
rect 4212 3654 4230 3672
rect 4212 3672 4230 3690
rect 4212 3690 4230 3708
rect 4212 3708 4230 3726
rect 4212 3726 4230 3744
rect 4212 3744 4230 3762
rect 4212 3762 4230 3780
rect 4212 3780 4230 3798
rect 4212 3798 4230 3816
rect 4212 3816 4230 3834
rect 4212 3834 4230 3852
rect 4212 3852 4230 3870
rect 4212 3870 4230 3888
rect 4212 3888 4230 3906
rect 4212 3906 4230 3924
rect 4212 3924 4230 3942
rect 4212 3942 4230 3960
rect 4212 3960 4230 3978
rect 4212 3978 4230 3996
rect 4212 3996 4230 4014
rect 4212 4014 4230 4032
rect 4212 4032 4230 4050
rect 4212 4050 4230 4068
rect 4212 4068 4230 4086
rect 4212 4086 4230 4104
rect 4212 4104 4230 4122
rect 4212 4122 4230 4140
rect 4212 4140 4230 4158
rect 4212 4158 4230 4176
rect 4212 4176 4230 4194
rect 4212 4194 4230 4212
rect 4212 4212 4230 4230
rect 4212 4230 4230 4248
rect 4212 4248 4230 4266
rect 4212 4266 4230 4284
rect 4212 4284 4230 4302
rect 4212 4302 4230 4320
rect 4212 4320 4230 4338
rect 4212 4338 4230 4356
rect 4212 4356 4230 4374
rect 4212 4374 4230 4392
rect 4212 4392 4230 4410
rect 4212 4410 4230 4428
rect 4212 4428 4230 4446
rect 4212 4446 4230 4464
rect 4212 4464 4230 4482
rect 4212 4482 4230 4500
rect 4212 4500 4230 4518
rect 4212 4518 4230 4536
rect 4212 4536 4230 4554
rect 4212 4554 4230 4572
rect 4212 4572 4230 4590
rect 4212 4590 4230 4608
rect 4212 4608 4230 4626
rect 4212 4626 4230 4644
rect 4212 4644 4230 4662
rect 4212 4662 4230 4680
rect 4212 4680 4230 4698
rect 4212 4698 4230 4716
rect 4212 4716 4230 4734
rect 4212 4734 4230 4752
rect 4212 4752 4230 4770
rect 4212 4770 4230 4788
rect 4212 4788 4230 4806
rect 4212 4806 4230 4824
rect 4212 4824 4230 4842
rect 4212 4842 4230 4860
rect 4212 4860 4230 4878
rect 4212 4878 4230 4896
rect 4212 4896 4230 4914
rect 4212 4914 4230 4932
rect 4212 4932 4230 4950
rect 4212 4950 4230 4968
rect 4212 4968 4230 4986
rect 4212 4986 4230 5004
rect 4212 5004 4230 5022
rect 4212 5022 4230 5040
rect 4212 5040 4230 5058
rect 4212 5058 4230 5076
rect 4212 5076 4230 5094
rect 4212 5094 4230 5112
rect 4212 5112 4230 5130
rect 4212 5130 4230 5148
rect 4212 5148 4230 5166
rect 4212 5166 4230 5184
rect 4212 5184 4230 5202
rect 4212 5202 4230 5220
rect 4212 5220 4230 5238
rect 4212 5238 4230 5256
rect 4212 5256 4230 5274
rect 4212 5274 4230 5292
rect 4212 5292 4230 5310
rect 4212 5310 4230 5328
rect 4212 5328 4230 5346
rect 4212 5346 4230 5364
rect 4212 5364 4230 5382
rect 4212 5382 4230 5400
rect 4212 5400 4230 5418
rect 4212 5418 4230 5436
rect 4212 5436 4230 5454
rect 4212 5454 4230 5472
rect 4212 5472 4230 5490
rect 4212 5490 4230 5508
rect 4212 5508 4230 5526
rect 4212 5526 4230 5544
rect 4212 5544 4230 5562
rect 4212 5562 4230 5580
rect 4212 5580 4230 5598
rect 4212 5598 4230 5616
rect 4212 5616 4230 5634
rect 4212 5634 4230 5652
rect 4212 5652 4230 5670
rect 4212 5670 4230 5688
rect 4212 5688 4230 5706
rect 4212 5706 4230 5724
rect 4212 5724 4230 5742
rect 4212 5742 4230 5760
rect 4212 5760 4230 5778
rect 4212 5778 4230 5796
rect 4212 5796 4230 5814
rect 4212 5814 4230 5832
rect 4212 5832 4230 5850
rect 4212 5850 4230 5868
rect 4212 5868 4230 5886
rect 4212 5886 4230 5904
rect 4212 5904 4230 5922
rect 4212 5922 4230 5940
rect 4212 5940 4230 5958
rect 4212 5958 4230 5976
rect 4212 5976 4230 5994
rect 4212 5994 4230 6012
rect 4212 6012 4230 6030
rect 4212 6030 4230 6048
rect 4212 6048 4230 6066
rect 4212 6066 4230 6084
rect 4212 6084 4230 6102
rect 4212 6102 4230 6120
rect 4212 6120 4230 6138
rect 4212 6138 4230 6156
rect 4212 6156 4230 6174
rect 4212 6174 4230 6192
rect 4212 6192 4230 6210
rect 4212 6210 4230 6228
rect 4212 6228 4230 6246
rect 4212 6246 4230 6264
rect 4212 6264 4230 6282
rect 4212 6282 4230 6300
rect 4212 6300 4230 6318
rect 4212 6318 4230 6336
rect 4212 6336 4230 6354
rect 4212 6354 4230 6372
rect 4212 6372 4230 6390
rect 4212 6390 4230 6408
rect 4212 6408 4230 6426
rect 4212 6426 4230 6444
rect 4212 6444 4230 6462
rect 4212 6462 4230 6480
rect 4212 6480 4230 6498
rect 4212 6498 4230 6516
rect 4212 6840 4230 6858
rect 4212 6858 4230 6876
rect 4212 6876 4230 6894
rect 4212 6894 4230 6912
rect 4212 6912 4230 6930
rect 4212 6930 4230 6948
rect 4212 6948 4230 6966
rect 4212 6966 4230 6984
rect 4212 6984 4230 7002
rect 4212 7002 4230 7020
rect 4212 7020 4230 7038
rect 4212 7038 4230 7056
rect 4212 7056 4230 7074
rect 4212 7074 4230 7092
rect 4212 7092 4230 7110
rect 4212 7110 4230 7128
rect 4212 7128 4230 7146
rect 4212 7146 4230 7164
rect 4212 7164 4230 7182
rect 4212 7182 4230 7200
rect 4212 7200 4230 7218
rect 4212 7218 4230 7236
rect 4230 54 4248 72
rect 4230 72 4248 90
rect 4230 90 4248 108
rect 4230 108 4248 126
rect 4230 126 4248 144
rect 4230 144 4248 162
rect 4230 162 4248 180
rect 4230 180 4248 198
rect 4230 198 4248 216
rect 4230 216 4248 234
rect 4230 234 4248 252
rect 4230 252 4248 270
rect 4230 270 4248 288
rect 4230 288 4248 306
rect 4230 306 4248 324
rect 4230 324 4248 342
rect 4230 342 4248 360
rect 4230 360 4248 378
rect 4230 378 4248 396
rect 4230 396 4248 414
rect 4230 414 4248 432
rect 4230 432 4248 450
rect 4230 450 4248 468
rect 4230 468 4248 486
rect 4230 486 4248 504
rect 4230 504 4248 522
rect 4230 522 4248 540
rect 4230 540 4248 558
rect 4230 558 4248 576
rect 4230 576 4248 594
rect 4230 594 4248 612
rect 4230 612 4248 630
rect 4230 630 4248 648
rect 4230 648 4248 666
rect 4230 666 4248 684
rect 4230 864 4248 882
rect 4230 882 4248 900
rect 4230 900 4248 918
rect 4230 918 4248 936
rect 4230 936 4248 954
rect 4230 954 4248 972
rect 4230 972 4248 990
rect 4230 990 4248 1008
rect 4230 1008 4248 1026
rect 4230 1026 4248 1044
rect 4230 1044 4248 1062
rect 4230 1062 4248 1080
rect 4230 1080 4248 1098
rect 4230 1098 4248 1116
rect 4230 1116 4248 1134
rect 4230 1134 4248 1152
rect 4230 1152 4248 1170
rect 4230 1170 4248 1188
rect 4230 1188 4248 1206
rect 4230 1206 4248 1224
rect 4230 1224 4248 1242
rect 4230 1242 4248 1260
rect 4230 1260 4248 1278
rect 4230 1278 4248 1296
rect 4230 1296 4248 1314
rect 4230 1314 4248 1332
rect 4230 1332 4248 1350
rect 4230 1350 4248 1368
rect 4230 1368 4248 1386
rect 4230 1386 4248 1404
rect 4230 1404 4248 1422
rect 4230 1422 4248 1440
rect 4230 1440 4248 1458
rect 4230 1458 4248 1476
rect 4230 1476 4248 1494
rect 4230 1494 4248 1512
rect 4230 1512 4248 1530
rect 4230 1530 4248 1548
rect 4230 1548 4248 1566
rect 4230 1566 4248 1584
rect 4230 1584 4248 1602
rect 4230 1602 4248 1620
rect 4230 1620 4248 1638
rect 4230 1638 4248 1656
rect 4230 1656 4248 1674
rect 4230 1674 4248 1692
rect 4230 1692 4248 1710
rect 4230 1710 4248 1728
rect 4230 1962 4248 1980
rect 4230 1980 4248 1998
rect 4230 1998 4248 2016
rect 4230 2016 4248 2034
rect 4230 2034 4248 2052
rect 4230 2052 4248 2070
rect 4230 2070 4248 2088
rect 4230 2088 4248 2106
rect 4230 2106 4248 2124
rect 4230 2124 4248 2142
rect 4230 2142 4248 2160
rect 4230 2160 4248 2178
rect 4230 2178 4248 2196
rect 4230 2196 4248 2214
rect 4230 2214 4248 2232
rect 4230 2232 4248 2250
rect 4230 2250 4248 2268
rect 4230 2268 4248 2286
rect 4230 2286 4248 2304
rect 4230 2304 4248 2322
rect 4230 2322 4248 2340
rect 4230 2340 4248 2358
rect 4230 2358 4248 2376
rect 4230 2376 4248 2394
rect 4230 2394 4248 2412
rect 4230 2412 4248 2430
rect 4230 2430 4248 2448
rect 4230 2448 4248 2466
rect 4230 2466 4248 2484
rect 4230 2484 4248 2502
rect 4230 2502 4248 2520
rect 4230 2520 4248 2538
rect 4230 2538 4248 2556
rect 4230 2556 4248 2574
rect 4230 2574 4248 2592
rect 4230 2592 4248 2610
rect 4230 2610 4248 2628
rect 4230 2628 4248 2646
rect 4230 2646 4248 2664
rect 4230 2664 4248 2682
rect 4230 2682 4248 2700
rect 4230 2700 4248 2718
rect 4230 2718 4248 2736
rect 4230 2736 4248 2754
rect 4230 2754 4248 2772
rect 4230 2772 4248 2790
rect 4230 2790 4248 2808
rect 4230 2808 4248 2826
rect 4230 2826 4248 2844
rect 4230 2844 4248 2862
rect 4230 2862 4248 2880
rect 4230 2880 4248 2898
rect 4230 2898 4248 2916
rect 4230 2916 4248 2934
rect 4230 2934 4248 2952
rect 4230 2952 4248 2970
rect 4230 2970 4248 2988
rect 4230 2988 4248 3006
rect 4230 3006 4248 3024
rect 4230 3024 4248 3042
rect 4230 3042 4248 3060
rect 4230 3060 4248 3078
rect 4230 3078 4248 3096
rect 4230 3096 4248 3114
rect 4230 3114 4248 3132
rect 4230 3132 4248 3150
rect 4230 3150 4248 3168
rect 4230 3168 4248 3186
rect 4230 3186 4248 3204
rect 4230 3204 4248 3222
rect 4230 3222 4248 3240
rect 4230 3240 4248 3258
rect 4230 3258 4248 3276
rect 4230 3276 4248 3294
rect 4230 3294 4248 3312
rect 4230 3312 4248 3330
rect 4230 3330 4248 3348
rect 4230 3348 4248 3366
rect 4230 3366 4248 3384
rect 4230 3384 4248 3402
rect 4230 3402 4248 3420
rect 4230 3420 4248 3438
rect 4230 3636 4248 3654
rect 4230 3654 4248 3672
rect 4230 3672 4248 3690
rect 4230 3690 4248 3708
rect 4230 3708 4248 3726
rect 4230 3726 4248 3744
rect 4230 3744 4248 3762
rect 4230 3762 4248 3780
rect 4230 3780 4248 3798
rect 4230 3798 4248 3816
rect 4230 3816 4248 3834
rect 4230 3834 4248 3852
rect 4230 3852 4248 3870
rect 4230 3870 4248 3888
rect 4230 3888 4248 3906
rect 4230 3906 4248 3924
rect 4230 3924 4248 3942
rect 4230 3942 4248 3960
rect 4230 3960 4248 3978
rect 4230 3978 4248 3996
rect 4230 3996 4248 4014
rect 4230 4014 4248 4032
rect 4230 4032 4248 4050
rect 4230 4050 4248 4068
rect 4230 4068 4248 4086
rect 4230 4086 4248 4104
rect 4230 4104 4248 4122
rect 4230 4122 4248 4140
rect 4230 4140 4248 4158
rect 4230 4158 4248 4176
rect 4230 4176 4248 4194
rect 4230 4194 4248 4212
rect 4230 4212 4248 4230
rect 4230 4230 4248 4248
rect 4230 4248 4248 4266
rect 4230 4266 4248 4284
rect 4230 4284 4248 4302
rect 4230 4302 4248 4320
rect 4230 4320 4248 4338
rect 4230 4338 4248 4356
rect 4230 4356 4248 4374
rect 4230 4374 4248 4392
rect 4230 4392 4248 4410
rect 4230 4410 4248 4428
rect 4230 4428 4248 4446
rect 4230 4446 4248 4464
rect 4230 4464 4248 4482
rect 4230 4482 4248 4500
rect 4230 4500 4248 4518
rect 4230 4518 4248 4536
rect 4230 4536 4248 4554
rect 4230 4554 4248 4572
rect 4230 4572 4248 4590
rect 4230 4590 4248 4608
rect 4230 4608 4248 4626
rect 4230 4626 4248 4644
rect 4230 4644 4248 4662
rect 4230 4662 4248 4680
rect 4230 4680 4248 4698
rect 4230 4698 4248 4716
rect 4230 4716 4248 4734
rect 4230 4734 4248 4752
rect 4230 4752 4248 4770
rect 4230 4770 4248 4788
rect 4230 4788 4248 4806
rect 4230 4806 4248 4824
rect 4230 4824 4248 4842
rect 4230 4842 4248 4860
rect 4230 4860 4248 4878
rect 4230 4878 4248 4896
rect 4230 4896 4248 4914
rect 4230 4914 4248 4932
rect 4230 4932 4248 4950
rect 4230 4950 4248 4968
rect 4230 4968 4248 4986
rect 4230 4986 4248 5004
rect 4230 5004 4248 5022
rect 4230 5022 4248 5040
rect 4230 5040 4248 5058
rect 4230 5058 4248 5076
rect 4230 5076 4248 5094
rect 4230 5094 4248 5112
rect 4230 5112 4248 5130
rect 4230 5130 4248 5148
rect 4230 5148 4248 5166
rect 4230 5166 4248 5184
rect 4230 5184 4248 5202
rect 4230 5202 4248 5220
rect 4230 5220 4248 5238
rect 4230 5238 4248 5256
rect 4230 5256 4248 5274
rect 4230 5274 4248 5292
rect 4230 5292 4248 5310
rect 4230 5310 4248 5328
rect 4230 5328 4248 5346
rect 4230 5346 4248 5364
rect 4230 5364 4248 5382
rect 4230 5382 4248 5400
rect 4230 5400 4248 5418
rect 4230 5418 4248 5436
rect 4230 5436 4248 5454
rect 4230 5454 4248 5472
rect 4230 5472 4248 5490
rect 4230 5490 4248 5508
rect 4230 5508 4248 5526
rect 4230 5526 4248 5544
rect 4230 5544 4248 5562
rect 4230 5562 4248 5580
rect 4230 5580 4248 5598
rect 4230 5598 4248 5616
rect 4230 5616 4248 5634
rect 4230 5634 4248 5652
rect 4230 5652 4248 5670
rect 4230 5670 4248 5688
rect 4230 5688 4248 5706
rect 4230 5706 4248 5724
rect 4230 5724 4248 5742
rect 4230 5742 4248 5760
rect 4230 5760 4248 5778
rect 4230 5778 4248 5796
rect 4230 5796 4248 5814
rect 4230 5814 4248 5832
rect 4230 5832 4248 5850
rect 4230 5850 4248 5868
rect 4230 5868 4248 5886
rect 4230 5886 4248 5904
rect 4230 5904 4248 5922
rect 4230 5922 4248 5940
rect 4230 5940 4248 5958
rect 4230 5958 4248 5976
rect 4230 5976 4248 5994
rect 4230 5994 4248 6012
rect 4230 6012 4248 6030
rect 4230 6030 4248 6048
rect 4230 6048 4248 6066
rect 4230 6066 4248 6084
rect 4230 6084 4248 6102
rect 4230 6102 4248 6120
rect 4230 6120 4248 6138
rect 4230 6138 4248 6156
rect 4230 6156 4248 6174
rect 4230 6174 4248 6192
rect 4230 6192 4248 6210
rect 4230 6210 4248 6228
rect 4230 6228 4248 6246
rect 4230 6246 4248 6264
rect 4230 6264 4248 6282
rect 4230 6282 4248 6300
rect 4230 6300 4248 6318
rect 4230 6318 4248 6336
rect 4230 6336 4248 6354
rect 4230 6354 4248 6372
rect 4230 6372 4248 6390
rect 4230 6390 4248 6408
rect 4230 6408 4248 6426
rect 4230 6426 4248 6444
rect 4230 6444 4248 6462
rect 4230 6462 4248 6480
rect 4230 6480 4248 6498
rect 4230 6498 4248 6516
rect 4230 6516 4248 6534
rect 4230 6534 4248 6552
rect 4230 6876 4248 6894
rect 4230 6894 4248 6912
rect 4230 6912 4248 6930
rect 4230 6930 4248 6948
rect 4230 6948 4248 6966
rect 4230 6966 4248 6984
rect 4230 6984 4248 7002
rect 4230 7002 4248 7020
rect 4230 7020 4248 7038
rect 4230 7038 4248 7056
rect 4230 7056 4248 7074
rect 4230 7074 4248 7092
rect 4230 7092 4248 7110
rect 4230 7110 4248 7128
rect 4230 7128 4248 7146
rect 4230 7146 4248 7164
rect 4230 7164 4248 7182
rect 4230 7182 4248 7200
rect 4230 7200 4248 7218
rect 4230 7218 4248 7236
rect 4248 54 4266 72
rect 4248 72 4266 90
rect 4248 90 4266 108
rect 4248 108 4266 126
rect 4248 126 4266 144
rect 4248 144 4266 162
rect 4248 162 4266 180
rect 4248 180 4266 198
rect 4248 198 4266 216
rect 4248 216 4266 234
rect 4248 234 4266 252
rect 4248 252 4266 270
rect 4248 270 4266 288
rect 4248 288 4266 306
rect 4248 306 4266 324
rect 4248 324 4266 342
rect 4248 342 4266 360
rect 4248 360 4266 378
rect 4248 378 4266 396
rect 4248 396 4266 414
rect 4248 414 4266 432
rect 4248 432 4266 450
rect 4248 450 4266 468
rect 4248 468 4266 486
rect 4248 486 4266 504
rect 4248 504 4266 522
rect 4248 522 4266 540
rect 4248 540 4266 558
rect 4248 558 4266 576
rect 4248 576 4266 594
rect 4248 594 4266 612
rect 4248 612 4266 630
rect 4248 630 4266 648
rect 4248 648 4266 666
rect 4248 666 4266 684
rect 4248 864 4266 882
rect 4248 882 4266 900
rect 4248 900 4266 918
rect 4248 918 4266 936
rect 4248 936 4266 954
rect 4248 954 4266 972
rect 4248 972 4266 990
rect 4248 990 4266 1008
rect 4248 1008 4266 1026
rect 4248 1026 4266 1044
rect 4248 1044 4266 1062
rect 4248 1062 4266 1080
rect 4248 1080 4266 1098
rect 4248 1098 4266 1116
rect 4248 1116 4266 1134
rect 4248 1134 4266 1152
rect 4248 1152 4266 1170
rect 4248 1170 4266 1188
rect 4248 1188 4266 1206
rect 4248 1206 4266 1224
rect 4248 1224 4266 1242
rect 4248 1242 4266 1260
rect 4248 1260 4266 1278
rect 4248 1278 4266 1296
rect 4248 1296 4266 1314
rect 4248 1314 4266 1332
rect 4248 1332 4266 1350
rect 4248 1350 4266 1368
rect 4248 1368 4266 1386
rect 4248 1386 4266 1404
rect 4248 1404 4266 1422
rect 4248 1422 4266 1440
rect 4248 1440 4266 1458
rect 4248 1458 4266 1476
rect 4248 1476 4266 1494
rect 4248 1494 4266 1512
rect 4248 1512 4266 1530
rect 4248 1530 4266 1548
rect 4248 1548 4266 1566
rect 4248 1566 4266 1584
rect 4248 1584 4266 1602
rect 4248 1602 4266 1620
rect 4248 1620 4266 1638
rect 4248 1638 4266 1656
rect 4248 1656 4266 1674
rect 4248 1674 4266 1692
rect 4248 1692 4266 1710
rect 4248 1710 4266 1728
rect 4248 1980 4266 1998
rect 4248 1998 4266 2016
rect 4248 2016 4266 2034
rect 4248 2034 4266 2052
rect 4248 2052 4266 2070
rect 4248 2070 4266 2088
rect 4248 2088 4266 2106
rect 4248 2106 4266 2124
rect 4248 2124 4266 2142
rect 4248 2142 4266 2160
rect 4248 2160 4266 2178
rect 4248 2178 4266 2196
rect 4248 2196 4266 2214
rect 4248 2214 4266 2232
rect 4248 2232 4266 2250
rect 4248 2250 4266 2268
rect 4248 2268 4266 2286
rect 4248 2286 4266 2304
rect 4248 2304 4266 2322
rect 4248 2322 4266 2340
rect 4248 2340 4266 2358
rect 4248 2358 4266 2376
rect 4248 2376 4266 2394
rect 4248 2394 4266 2412
rect 4248 2412 4266 2430
rect 4248 2430 4266 2448
rect 4248 2448 4266 2466
rect 4248 2466 4266 2484
rect 4248 2484 4266 2502
rect 4248 2502 4266 2520
rect 4248 2520 4266 2538
rect 4248 2538 4266 2556
rect 4248 2556 4266 2574
rect 4248 2574 4266 2592
rect 4248 2592 4266 2610
rect 4248 2610 4266 2628
rect 4248 2628 4266 2646
rect 4248 2646 4266 2664
rect 4248 2664 4266 2682
rect 4248 2682 4266 2700
rect 4248 2700 4266 2718
rect 4248 2718 4266 2736
rect 4248 2736 4266 2754
rect 4248 2754 4266 2772
rect 4248 2772 4266 2790
rect 4248 2790 4266 2808
rect 4248 2808 4266 2826
rect 4248 2826 4266 2844
rect 4248 2844 4266 2862
rect 4248 2862 4266 2880
rect 4248 2880 4266 2898
rect 4248 2898 4266 2916
rect 4248 2916 4266 2934
rect 4248 2934 4266 2952
rect 4248 2952 4266 2970
rect 4248 2970 4266 2988
rect 4248 2988 4266 3006
rect 4248 3006 4266 3024
rect 4248 3024 4266 3042
rect 4248 3042 4266 3060
rect 4248 3060 4266 3078
rect 4248 3078 4266 3096
rect 4248 3096 4266 3114
rect 4248 3114 4266 3132
rect 4248 3132 4266 3150
rect 4248 3150 4266 3168
rect 4248 3168 4266 3186
rect 4248 3186 4266 3204
rect 4248 3204 4266 3222
rect 4248 3222 4266 3240
rect 4248 3240 4266 3258
rect 4248 3258 4266 3276
rect 4248 3276 4266 3294
rect 4248 3294 4266 3312
rect 4248 3312 4266 3330
rect 4248 3330 4266 3348
rect 4248 3348 4266 3366
rect 4248 3366 4266 3384
rect 4248 3384 4266 3402
rect 4248 3402 4266 3420
rect 4248 3420 4266 3438
rect 4248 3438 4266 3456
rect 4248 3672 4266 3690
rect 4248 3690 4266 3708
rect 4248 3708 4266 3726
rect 4248 3726 4266 3744
rect 4248 3744 4266 3762
rect 4248 3762 4266 3780
rect 4248 3780 4266 3798
rect 4248 3798 4266 3816
rect 4248 3816 4266 3834
rect 4248 3834 4266 3852
rect 4248 3852 4266 3870
rect 4248 3870 4266 3888
rect 4248 3888 4266 3906
rect 4248 3906 4266 3924
rect 4248 3924 4266 3942
rect 4248 3942 4266 3960
rect 4248 3960 4266 3978
rect 4248 3978 4266 3996
rect 4248 3996 4266 4014
rect 4248 4014 4266 4032
rect 4248 4032 4266 4050
rect 4248 4050 4266 4068
rect 4248 4068 4266 4086
rect 4248 4086 4266 4104
rect 4248 4104 4266 4122
rect 4248 4122 4266 4140
rect 4248 4140 4266 4158
rect 4248 4158 4266 4176
rect 4248 4176 4266 4194
rect 4248 4194 4266 4212
rect 4248 4212 4266 4230
rect 4248 4230 4266 4248
rect 4248 4248 4266 4266
rect 4248 4266 4266 4284
rect 4248 4284 4266 4302
rect 4248 4302 4266 4320
rect 4248 4320 4266 4338
rect 4248 4338 4266 4356
rect 4248 4356 4266 4374
rect 4248 4374 4266 4392
rect 4248 4392 4266 4410
rect 4248 4410 4266 4428
rect 4248 4428 4266 4446
rect 4248 4446 4266 4464
rect 4248 4464 4266 4482
rect 4248 4482 4266 4500
rect 4248 4500 4266 4518
rect 4248 4518 4266 4536
rect 4248 4536 4266 4554
rect 4248 4554 4266 4572
rect 4248 4572 4266 4590
rect 4248 4590 4266 4608
rect 4248 4608 4266 4626
rect 4248 4626 4266 4644
rect 4248 4644 4266 4662
rect 4248 4662 4266 4680
rect 4248 4680 4266 4698
rect 4248 4698 4266 4716
rect 4248 4716 4266 4734
rect 4248 4734 4266 4752
rect 4248 4752 4266 4770
rect 4248 4770 4266 4788
rect 4248 4788 4266 4806
rect 4248 4806 4266 4824
rect 4248 4824 4266 4842
rect 4248 4842 4266 4860
rect 4248 4860 4266 4878
rect 4248 4878 4266 4896
rect 4248 4896 4266 4914
rect 4248 4914 4266 4932
rect 4248 4932 4266 4950
rect 4248 4950 4266 4968
rect 4248 4968 4266 4986
rect 4248 4986 4266 5004
rect 4248 5004 4266 5022
rect 4248 5022 4266 5040
rect 4248 5040 4266 5058
rect 4248 5058 4266 5076
rect 4248 5076 4266 5094
rect 4248 5094 4266 5112
rect 4248 5112 4266 5130
rect 4248 5130 4266 5148
rect 4248 5148 4266 5166
rect 4248 5166 4266 5184
rect 4248 5184 4266 5202
rect 4248 5202 4266 5220
rect 4248 5220 4266 5238
rect 4248 5238 4266 5256
rect 4248 5256 4266 5274
rect 4248 5274 4266 5292
rect 4248 5292 4266 5310
rect 4248 5310 4266 5328
rect 4248 5328 4266 5346
rect 4248 5346 4266 5364
rect 4248 5364 4266 5382
rect 4248 5382 4266 5400
rect 4248 5400 4266 5418
rect 4248 5418 4266 5436
rect 4248 5436 4266 5454
rect 4248 5454 4266 5472
rect 4248 5472 4266 5490
rect 4248 5490 4266 5508
rect 4248 5508 4266 5526
rect 4248 5526 4266 5544
rect 4248 5544 4266 5562
rect 4248 5562 4266 5580
rect 4248 5580 4266 5598
rect 4248 5598 4266 5616
rect 4248 5616 4266 5634
rect 4248 5634 4266 5652
rect 4248 5652 4266 5670
rect 4248 5670 4266 5688
rect 4248 5688 4266 5706
rect 4248 5706 4266 5724
rect 4248 5724 4266 5742
rect 4248 5742 4266 5760
rect 4248 5760 4266 5778
rect 4248 5778 4266 5796
rect 4248 5796 4266 5814
rect 4248 5814 4266 5832
rect 4248 5832 4266 5850
rect 4248 5850 4266 5868
rect 4248 5868 4266 5886
rect 4248 5886 4266 5904
rect 4248 5904 4266 5922
rect 4248 5922 4266 5940
rect 4248 5940 4266 5958
rect 4248 5958 4266 5976
rect 4248 5976 4266 5994
rect 4248 5994 4266 6012
rect 4248 6012 4266 6030
rect 4248 6030 4266 6048
rect 4248 6048 4266 6066
rect 4248 6066 4266 6084
rect 4248 6084 4266 6102
rect 4248 6102 4266 6120
rect 4248 6120 4266 6138
rect 4248 6138 4266 6156
rect 4248 6156 4266 6174
rect 4248 6174 4266 6192
rect 4248 6192 4266 6210
rect 4248 6210 4266 6228
rect 4248 6228 4266 6246
rect 4248 6246 4266 6264
rect 4248 6264 4266 6282
rect 4248 6282 4266 6300
rect 4248 6300 4266 6318
rect 4248 6318 4266 6336
rect 4248 6336 4266 6354
rect 4248 6354 4266 6372
rect 4248 6372 4266 6390
rect 4248 6390 4266 6408
rect 4248 6408 4266 6426
rect 4248 6426 4266 6444
rect 4248 6444 4266 6462
rect 4248 6462 4266 6480
rect 4248 6480 4266 6498
rect 4248 6498 4266 6516
rect 4248 6516 4266 6534
rect 4248 6534 4266 6552
rect 4248 6552 4266 6570
rect 4248 6570 4266 6588
rect 4248 6912 4266 6930
rect 4248 6930 4266 6948
rect 4248 6948 4266 6966
rect 4248 6966 4266 6984
rect 4248 6984 4266 7002
rect 4248 7002 4266 7020
rect 4248 7020 4266 7038
rect 4248 7038 4266 7056
rect 4248 7056 4266 7074
rect 4248 7074 4266 7092
rect 4248 7092 4266 7110
rect 4248 7110 4266 7128
rect 4248 7128 4266 7146
rect 4248 7146 4266 7164
rect 4248 7164 4266 7182
rect 4248 7182 4266 7200
rect 4248 7200 4266 7218
rect 4248 7218 4266 7236
rect 4266 54 4284 72
rect 4266 72 4284 90
rect 4266 90 4284 108
rect 4266 108 4284 126
rect 4266 126 4284 144
rect 4266 144 4284 162
rect 4266 162 4284 180
rect 4266 180 4284 198
rect 4266 198 4284 216
rect 4266 216 4284 234
rect 4266 234 4284 252
rect 4266 252 4284 270
rect 4266 270 4284 288
rect 4266 288 4284 306
rect 4266 306 4284 324
rect 4266 324 4284 342
rect 4266 342 4284 360
rect 4266 360 4284 378
rect 4266 378 4284 396
rect 4266 396 4284 414
rect 4266 414 4284 432
rect 4266 432 4284 450
rect 4266 450 4284 468
rect 4266 468 4284 486
rect 4266 486 4284 504
rect 4266 504 4284 522
rect 4266 522 4284 540
rect 4266 540 4284 558
rect 4266 558 4284 576
rect 4266 576 4284 594
rect 4266 594 4284 612
rect 4266 612 4284 630
rect 4266 630 4284 648
rect 4266 648 4284 666
rect 4266 666 4284 684
rect 4266 864 4284 882
rect 4266 882 4284 900
rect 4266 900 4284 918
rect 4266 918 4284 936
rect 4266 936 4284 954
rect 4266 954 4284 972
rect 4266 972 4284 990
rect 4266 990 4284 1008
rect 4266 1008 4284 1026
rect 4266 1026 4284 1044
rect 4266 1044 4284 1062
rect 4266 1062 4284 1080
rect 4266 1080 4284 1098
rect 4266 1098 4284 1116
rect 4266 1116 4284 1134
rect 4266 1134 4284 1152
rect 4266 1152 4284 1170
rect 4266 1170 4284 1188
rect 4266 1188 4284 1206
rect 4266 1206 4284 1224
rect 4266 1224 4284 1242
rect 4266 1242 4284 1260
rect 4266 1260 4284 1278
rect 4266 1278 4284 1296
rect 4266 1296 4284 1314
rect 4266 1314 4284 1332
rect 4266 1332 4284 1350
rect 4266 1350 4284 1368
rect 4266 1368 4284 1386
rect 4266 1386 4284 1404
rect 4266 1404 4284 1422
rect 4266 1422 4284 1440
rect 4266 1440 4284 1458
rect 4266 1458 4284 1476
rect 4266 1476 4284 1494
rect 4266 1494 4284 1512
rect 4266 1512 4284 1530
rect 4266 1530 4284 1548
rect 4266 1548 4284 1566
rect 4266 1566 4284 1584
rect 4266 1584 4284 1602
rect 4266 1602 4284 1620
rect 4266 1620 4284 1638
rect 4266 1638 4284 1656
rect 4266 1656 4284 1674
rect 4266 1674 4284 1692
rect 4266 1692 4284 1710
rect 4266 1710 4284 1728
rect 4266 1728 4284 1746
rect 4266 1980 4284 1998
rect 4266 1998 4284 2016
rect 4266 2016 4284 2034
rect 4266 2034 4284 2052
rect 4266 2052 4284 2070
rect 4266 2070 4284 2088
rect 4266 2088 4284 2106
rect 4266 2106 4284 2124
rect 4266 2124 4284 2142
rect 4266 2142 4284 2160
rect 4266 2160 4284 2178
rect 4266 2178 4284 2196
rect 4266 2196 4284 2214
rect 4266 2214 4284 2232
rect 4266 2232 4284 2250
rect 4266 2250 4284 2268
rect 4266 2268 4284 2286
rect 4266 2286 4284 2304
rect 4266 2304 4284 2322
rect 4266 2322 4284 2340
rect 4266 2340 4284 2358
rect 4266 2358 4284 2376
rect 4266 2376 4284 2394
rect 4266 2394 4284 2412
rect 4266 2412 4284 2430
rect 4266 2430 4284 2448
rect 4266 2448 4284 2466
rect 4266 2466 4284 2484
rect 4266 2484 4284 2502
rect 4266 2502 4284 2520
rect 4266 2520 4284 2538
rect 4266 2538 4284 2556
rect 4266 2556 4284 2574
rect 4266 2574 4284 2592
rect 4266 2592 4284 2610
rect 4266 2610 4284 2628
rect 4266 2628 4284 2646
rect 4266 2646 4284 2664
rect 4266 2664 4284 2682
rect 4266 2682 4284 2700
rect 4266 2700 4284 2718
rect 4266 2718 4284 2736
rect 4266 2736 4284 2754
rect 4266 2754 4284 2772
rect 4266 2772 4284 2790
rect 4266 2790 4284 2808
rect 4266 2808 4284 2826
rect 4266 2826 4284 2844
rect 4266 2844 4284 2862
rect 4266 2862 4284 2880
rect 4266 2880 4284 2898
rect 4266 2898 4284 2916
rect 4266 2916 4284 2934
rect 4266 2934 4284 2952
rect 4266 2952 4284 2970
rect 4266 2970 4284 2988
rect 4266 2988 4284 3006
rect 4266 3006 4284 3024
rect 4266 3024 4284 3042
rect 4266 3042 4284 3060
rect 4266 3060 4284 3078
rect 4266 3078 4284 3096
rect 4266 3096 4284 3114
rect 4266 3114 4284 3132
rect 4266 3132 4284 3150
rect 4266 3150 4284 3168
rect 4266 3168 4284 3186
rect 4266 3186 4284 3204
rect 4266 3204 4284 3222
rect 4266 3222 4284 3240
rect 4266 3240 4284 3258
rect 4266 3258 4284 3276
rect 4266 3276 4284 3294
rect 4266 3294 4284 3312
rect 4266 3312 4284 3330
rect 4266 3330 4284 3348
rect 4266 3348 4284 3366
rect 4266 3366 4284 3384
rect 4266 3384 4284 3402
rect 4266 3402 4284 3420
rect 4266 3420 4284 3438
rect 4266 3438 4284 3456
rect 4266 3456 4284 3474
rect 4266 3690 4284 3708
rect 4266 3708 4284 3726
rect 4266 3726 4284 3744
rect 4266 3744 4284 3762
rect 4266 3762 4284 3780
rect 4266 3780 4284 3798
rect 4266 3798 4284 3816
rect 4266 3816 4284 3834
rect 4266 3834 4284 3852
rect 4266 3852 4284 3870
rect 4266 3870 4284 3888
rect 4266 3888 4284 3906
rect 4266 3906 4284 3924
rect 4266 3924 4284 3942
rect 4266 3942 4284 3960
rect 4266 3960 4284 3978
rect 4266 3978 4284 3996
rect 4266 3996 4284 4014
rect 4266 4014 4284 4032
rect 4266 4032 4284 4050
rect 4266 4050 4284 4068
rect 4266 4068 4284 4086
rect 4266 4086 4284 4104
rect 4266 4104 4284 4122
rect 4266 4122 4284 4140
rect 4266 4140 4284 4158
rect 4266 4158 4284 4176
rect 4266 4176 4284 4194
rect 4266 4194 4284 4212
rect 4266 4212 4284 4230
rect 4266 4230 4284 4248
rect 4266 4248 4284 4266
rect 4266 4266 4284 4284
rect 4266 4284 4284 4302
rect 4266 4302 4284 4320
rect 4266 4320 4284 4338
rect 4266 4338 4284 4356
rect 4266 4356 4284 4374
rect 4266 4374 4284 4392
rect 4266 4392 4284 4410
rect 4266 4410 4284 4428
rect 4266 4428 4284 4446
rect 4266 4446 4284 4464
rect 4266 4464 4284 4482
rect 4266 4482 4284 4500
rect 4266 4500 4284 4518
rect 4266 4518 4284 4536
rect 4266 4536 4284 4554
rect 4266 4554 4284 4572
rect 4266 4572 4284 4590
rect 4266 4590 4284 4608
rect 4266 4608 4284 4626
rect 4266 4626 4284 4644
rect 4266 4644 4284 4662
rect 4266 4662 4284 4680
rect 4266 4680 4284 4698
rect 4266 4698 4284 4716
rect 4266 4716 4284 4734
rect 4266 4734 4284 4752
rect 4266 4752 4284 4770
rect 4266 4770 4284 4788
rect 4266 4788 4284 4806
rect 4266 4806 4284 4824
rect 4266 4824 4284 4842
rect 4266 4842 4284 4860
rect 4266 4860 4284 4878
rect 4266 4878 4284 4896
rect 4266 4896 4284 4914
rect 4266 4914 4284 4932
rect 4266 4932 4284 4950
rect 4266 4950 4284 4968
rect 4266 4968 4284 4986
rect 4266 4986 4284 5004
rect 4266 5004 4284 5022
rect 4266 5022 4284 5040
rect 4266 5040 4284 5058
rect 4266 5058 4284 5076
rect 4266 5076 4284 5094
rect 4266 5094 4284 5112
rect 4266 5112 4284 5130
rect 4266 5130 4284 5148
rect 4266 5148 4284 5166
rect 4266 5166 4284 5184
rect 4266 5184 4284 5202
rect 4266 5202 4284 5220
rect 4266 5220 4284 5238
rect 4266 5238 4284 5256
rect 4266 5256 4284 5274
rect 4266 5274 4284 5292
rect 4266 5292 4284 5310
rect 4266 5310 4284 5328
rect 4266 5328 4284 5346
rect 4266 5346 4284 5364
rect 4266 5364 4284 5382
rect 4266 5382 4284 5400
rect 4266 5400 4284 5418
rect 4266 5418 4284 5436
rect 4266 5436 4284 5454
rect 4266 5454 4284 5472
rect 4266 5472 4284 5490
rect 4266 5490 4284 5508
rect 4266 5508 4284 5526
rect 4266 5526 4284 5544
rect 4266 5544 4284 5562
rect 4266 5562 4284 5580
rect 4266 5580 4284 5598
rect 4266 5598 4284 5616
rect 4266 5616 4284 5634
rect 4266 5634 4284 5652
rect 4266 5652 4284 5670
rect 4266 5670 4284 5688
rect 4266 5688 4284 5706
rect 4266 5706 4284 5724
rect 4266 5724 4284 5742
rect 4266 5742 4284 5760
rect 4266 5760 4284 5778
rect 4266 5778 4284 5796
rect 4266 5796 4284 5814
rect 4266 5814 4284 5832
rect 4266 5832 4284 5850
rect 4266 5850 4284 5868
rect 4266 5868 4284 5886
rect 4266 5886 4284 5904
rect 4266 5904 4284 5922
rect 4266 5922 4284 5940
rect 4266 5940 4284 5958
rect 4266 5958 4284 5976
rect 4266 5976 4284 5994
rect 4266 5994 4284 6012
rect 4266 6012 4284 6030
rect 4266 6030 4284 6048
rect 4266 6048 4284 6066
rect 4266 6066 4284 6084
rect 4266 6084 4284 6102
rect 4266 6102 4284 6120
rect 4266 6120 4284 6138
rect 4266 6138 4284 6156
rect 4266 6156 4284 6174
rect 4266 6174 4284 6192
rect 4266 6192 4284 6210
rect 4266 6210 4284 6228
rect 4266 6228 4284 6246
rect 4266 6246 4284 6264
rect 4266 6264 4284 6282
rect 4266 6282 4284 6300
rect 4266 6300 4284 6318
rect 4266 6318 4284 6336
rect 4266 6336 4284 6354
rect 4266 6354 4284 6372
rect 4266 6372 4284 6390
rect 4266 6390 4284 6408
rect 4266 6408 4284 6426
rect 4266 6426 4284 6444
rect 4266 6444 4284 6462
rect 4266 6462 4284 6480
rect 4266 6480 4284 6498
rect 4266 6498 4284 6516
rect 4266 6516 4284 6534
rect 4266 6534 4284 6552
rect 4266 6552 4284 6570
rect 4266 6570 4284 6588
rect 4266 6588 4284 6606
rect 4266 6606 4284 6624
rect 4266 6948 4284 6966
rect 4266 6966 4284 6984
rect 4266 6984 4284 7002
rect 4266 7002 4284 7020
rect 4266 7020 4284 7038
rect 4266 7038 4284 7056
rect 4266 7056 4284 7074
rect 4266 7074 4284 7092
rect 4266 7092 4284 7110
rect 4266 7110 4284 7128
rect 4266 7128 4284 7146
rect 4266 7146 4284 7164
rect 4266 7164 4284 7182
rect 4266 7182 4284 7200
rect 4266 7200 4284 7218
rect 4266 7218 4284 7236
rect 4284 54 4302 72
rect 4284 72 4302 90
rect 4284 90 4302 108
rect 4284 108 4302 126
rect 4284 126 4302 144
rect 4284 144 4302 162
rect 4284 162 4302 180
rect 4284 180 4302 198
rect 4284 198 4302 216
rect 4284 216 4302 234
rect 4284 234 4302 252
rect 4284 252 4302 270
rect 4284 270 4302 288
rect 4284 288 4302 306
rect 4284 306 4302 324
rect 4284 324 4302 342
rect 4284 342 4302 360
rect 4284 360 4302 378
rect 4284 378 4302 396
rect 4284 396 4302 414
rect 4284 414 4302 432
rect 4284 432 4302 450
rect 4284 450 4302 468
rect 4284 468 4302 486
rect 4284 486 4302 504
rect 4284 504 4302 522
rect 4284 522 4302 540
rect 4284 540 4302 558
rect 4284 558 4302 576
rect 4284 576 4302 594
rect 4284 594 4302 612
rect 4284 612 4302 630
rect 4284 630 4302 648
rect 4284 648 4302 666
rect 4284 666 4302 684
rect 4284 864 4302 882
rect 4284 882 4302 900
rect 4284 900 4302 918
rect 4284 918 4302 936
rect 4284 936 4302 954
rect 4284 954 4302 972
rect 4284 972 4302 990
rect 4284 990 4302 1008
rect 4284 1008 4302 1026
rect 4284 1026 4302 1044
rect 4284 1044 4302 1062
rect 4284 1062 4302 1080
rect 4284 1080 4302 1098
rect 4284 1098 4302 1116
rect 4284 1116 4302 1134
rect 4284 1134 4302 1152
rect 4284 1152 4302 1170
rect 4284 1170 4302 1188
rect 4284 1188 4302 1206
rect 4284 1206 4302 1224
rect 4284 1224 4302 1242
rect 4284 1242 4302 1260
rect 4284 1260 4302 1278
rect 4284 1278 4302 1296
rect 4284 1296 4302 1314
rect 4284 1314 4302 1332
rect 4284 1332 4302 1350
rect 4284 1350 4302 1368
rect 4284 1368 4302 1386
rect 4284 1386 4302 1404
rect 4284 1404 4302 1422
rect 4284 1422 4302 1440
rect 4284 1440 4302 1458
rect 4284 1458 4302 1476
rect 4284 1476 4302 1494
rect 4284 1494 4302 1512
rect 4284 1512 4302 1530
rect 4284 1530 4302 1548
rect 4284 1548 4302 1566
rect 4284 1566 4302 1584
rect 4284 1584 4302 1602
rect 4284 1602 4302 1620
rect 4284 1620 4302 1638
rect 4284 1638 4302 1656
rect 4284 1656 4302 1674
rect 4284 1674 4302 1692
rect 4284 1692 4302 1710
rect 4284 1710 4302 1728
rect 4284 1728 4302 1746
rect 4284 1746 4302 1764
rect 4284 1998 4302 2016
rect 4284 2016 4302 2034
rect 4284 2034 4302 2052
rect 4284 2052 4302 2070
rect 4284 2070 4302 2088
rect 4284 2088 4302 2106
rect 4284 2106 4302 2124
rect 4284 2124 4302 2142
rect 4284 2142 4302 2160
rect 4284 2160 4302 2178
rect 4284 2178 4302 2196
rect 4284 2196 4302 2214
rect 4284 2214 4302 2232
rect 4284 2232 4302 2250
rect 4284 2250 4302 2268
rect 4284 2268 4302 2286
rect 4284 2286 4302 2304
rect 4284 2304 4302 2322
rect 4284 2322 4302 2340
rect 4284 2340 4302 2358
rect 4284 2358 4302 2376
rect 4284 2376 4302 2394
rect 4284 2394 4302 2412
rect 4284 2412 4302 2430
rect 4284 2430 4302 2448
rect 4284 2448 4302 2466
rect 4284 2466 4302 2484
rect 4284 2484 4302 2502
rect 4284 2502 4302 2520
rect 4284 2520 4302 2538
rect 4284 2538 4302 2556
rect 4284 2556 4302 2574
rect 4284 2574 4302 2592
rect 4284 2592 4302 2610
rect 4284 2610 4302 2628
rect 4284 2628 4302 2646
rect 4284 2646 4302 2664
rect 4284 2664 4302 2682
rect 4284 2682 4302 2700
rect 4284 2700 4302 2718
rect 4284 2718 4302 2736
rect 4284 2736 4302 2754
rect 4284 2754 4302 2772
rect 4284 2772 4302 2790
rect 4284 2790 4302 2808
rect 4284 2808 4302 2826
rect 4284 2826 4302 2844
rect 4284 2844 4302 2862
rect 4284 2862 4302 2880
rect 4284 2880 4302 2898
rect 4284 2898 4302 2916
rect 4284 2916 4302 2934
rect 4284 2934 4302 2952
rect 4284 2952 4302 2970
rect 4284 2970 4302 2988
rect 4284 2988 4302 3006
rect 4284 3006 4302 3024
rect 4284 3024 4302 3042
rect 4284 3042 4302 3060
rect 4284 3060 4302 3078
rect 4284 3078 4302 3096
rect 4284 3096 4302 3114
rect 4284 3114 4302 3132
rect 4284 3132 4302 3150
rect 4284 3150 4302 3168
rect 4284 3168 4302 3186
rect 4284 3186 4302 3204
rect 4284 3204 4302 3222
rect 4284 3222 4302 3240
rect 4284 3240 4302 3258
rect 4284 3258 4302 3276
rect 4284 3276 4302 3294
rect 4284 3294 4302 3312
rect 4284 3312 4302 3330
rect 4284 3330 4302 3348
rect 4284 3348 4302 3366
rect 4284 3366 4302 3384
rect 4284 3384 4302 3402
rect 4284 3402 4302 3420
rect 4284 3420 4302 3438
rect 4284 3438 4302 3456
rect 4284 3456 4302 3474
rect 4284 3474 4302 3492
rect 4284 3492 4302 3510
rect 4284 3708 4302 3726
rect 4284 3726 4302 3744
rect 4284 3744 4302 3762
rect 4284 3762 4302 3780
rect 4284 3780 4302 3798
rect 4284 3798 4302 3816
rect 4284 3816 4302 3834
rect 4284 3834 4302 3852
rect 4284 3852 4302 3870
rect 4284 3870 4302 3888
rect 4284 3888 4302 3906
rect 4284 3906 4302 3924
rect 4284 3924 4302 3942
rect 4284 3942 4302 3960
rect 4284 3960 4302 3978
rect 4284 3978 4302 3996
rect 4284 3996 4302 4014
rect 4284 4014 4302 4032
rect 4284 4032 4302 4050
rect 4284 4050 4302 4068
rect 4284 4068 4302 4086
rect 4284 4086 4302 4104
rect 4284 4104 4302 4122
rect 4284 4122 4302 4140
rect 4284 4140 4302 4158
rect 4284 4158 4302 4176
rect 4284 4176 4302 4194
rect 4284 4194 4302 4212
rect 4284 4212 4302 4230
rect 4284 4230 4302 4248
rect 4284 4248 4302 4266
rect 4284 4266 4302 4284
rect 4284 4284 4302 4302
rect 4284 4302 4302 4320
rect 4284 4320 4302 4338
rect 4284 4338 4302 4356
rect 4284 4356 4302 4374
rect 4284 4374 4302 4392
rect 4284 4392 4302 4410
rect 4284 4410 4302 4428
rect 4284 4428 4302 4446
rect 4284 4446 4302 4464
rect 4284 4464 4302 4482
rect 4284 4482 4302 4500
rect 4284 4500 4302 4518
rect 4284 4518 4302 4536
rect 4284 4536 4302 4554
rect 4284 4554 4302 4572
rect 4284 4572 4302 4590
rect 4284 4590 4302 4608
rect 4284 4608 4302 4626
rect 4284 4626 4302 4644
rect 4284 4644 4302 4662
rect 4284 4662 4302 4680
rect 4284 4680 4302 4698
rect 4284 4698 4302 4716
rect 4284 4716 4302 4734
rect 4284 4734 4302 4752
rect 4284 4752 4302 4770
rect 4284 4770 4302 4788
rect 4284 4788 4302 4806
rect 4284 4806 4302 4824
rect 4284 4824 4302 4842
rect 4284 4842 4302 4860
rect 4284 4860 4302 4878
rect 4284 4878 4302 4896
rect 4284 4896 4302 4914
rect 4284 4914 4302 4932
rect 4284 4932 4302 4950
rect 4284 4950 4302 4968
rect 4284 4968 4302 4986
rect 4284 4986 4302 5004
rect 4284 5004 4302 5022
rect 4284 5022 4302 5040
rect 4284 5040 4302 5058
rect 4284 5058 4302 5076
rect 4284 5076 4302 5094
rect 4284 5094 4302 5112
rect 4284 5112 4302 5130
rect 4284 5130 4302 5148
rect 4284 5148 4302 5166
rect 4284 5166 4302 5184
rect 4284 5184 4302 5202
rect 4284 5202 4302 5220
rect 4284 5220 4302 5238
rect 4284 5238 4302 5256
rect 4284 5256 4302 5274
rect 4284 5274 4302 5292
rect 4284 5292 4302 5310
rect 4284 5310 4302 5328
rect 4284 5328 4302 5346
rect 4284 5346 4302 5364
rect 4284 5364 4302 5382
rect 4284 5382 4302 5400
rect 4284 5400 4302 5418
rect 4284 5418 4302 5436
rect 4284 5436 4302 5454
rect 4284 5454 4302 5472
rect 4284 5472 4302 5490
rect 4284 5490 4302 5508
rect 4284 5508 4302 5526
rect 4284 5526 4302 5544
rect 4284 5544 4302 5562
rect 4284 5562 4302 5580
rect 4284 5580 4302 5598
rect 4284 5598 4302 5616
rect 4284 5616 4302 5634
rect 4284 5634 4302 5652
rect 4284 5652 4302 5670
rect 4284 5670 4302 5688
rect 4284 5688 4302 5706
rect 4284 5706 4302 5724
rect 4284 5724 4302 5742
rect 4284 5742 4302 5760
rect 4284 5760 4302 5778
rect 4284 5778 4302 5796
rect 4284 5796 4302 5814
rect 4284 5814 4302 5832
rect 4284 5832 4302 5850
rect 4284 5850 4302 5868
rect 4284 5868 4302 5886
rect 4284 5886 4302 5904
rect 4284 5904 4302 5922
rect 4284 5922 4302 5940
rect 4284 5940 4302 5958
rect 4284 5958 4302 5976
rect 4284 5976 4302 5994
rect 4284 5994 4302 6012
rect 4284 6012 4302 6030
rect 4284 6030 4302 6048
rect 4284 6048 4302 6066
rect 4284 6066 4302 6084
rect 4284 6084 4302 6102
rect 4284 6102 4302 6120
rect 4284 6120 4302 6138
rect 4284 6138 4302 6156
rect 4284 6156 4302 6174
rect 4284 6174 4302 6192
rect 4284 6192 4302 6210
rect 4284 6210 4302 6228
rect 4284 6228 4302 6246
rect 4284 6246 4302 6264
rect 4284 6264 4302 6282
rect 4284 6282 4302 6300
rect 4284 6300 4302 6318
rect 4284 6318 4302 6336
rect 4284 6336 4302 6354
rect 4284 6354 4302 6372
rect 4284 6372 4302 6390
rect 4284 6390 4302 6408
rect 4284 6408 4302 6426
rect 4284 6426 4302 6444
rect 4284 6444 4302 6462
rect 4284 6462 4302 6480
rect 4284 6480 4302 6498
rect 4284 6498 4302 6516
rect 4284 6516 4302 6534
rect 4284 6534 4302 6552
rect 4284 6552 4302 6570
rect 4284 6570 4302 6588
rect 4284 6588 4302 6606
rect 4284 6606 4302 6624
rect 4284 6624 4302 6642
rect 4284 6642 4302 6660
rect 4284 6984 4302 7002
rect 4284 7002 4302 7020
rect 4284 7020 4302 7038
rect 4284 7038 4302 7056
rect 4284 7056 4302 7074
rect 4284 7074 4302 7092
rect 4284 7092 4302 7110
rect 4284 7110 4302 7128
rect 4284 7128 4302 7146
rect 4284 7146 4302 7164
rect 4284 7164 4302 7182
rect 4284 7182 4302 7200
rect 4284 7200 4302 7218
rect 4302 54 4320 72
rect 4302 72 4320 90
rect 4302 90 4320 108
rect 4302 108 4320 126
rect 4302 126 4320 144
rect 4302 144 4320 162
rect 4302 162 4320 180
rect 4302 180 4320 198
rect 4302 198 4320 216
rect 4302 216 4320 234
rect 4302 234 4320 252
rect 4302 252 4320 270
rect 4302 270 4320 288
rect 4302 288 4320 306
rect 4302 306 4320 324
rect 4302 324 4320 342
rect 4302 342 4320 360
rect 4302 360 4320 378
rect 4302 378 4320 396
rect 4302 396 4320 414
rect 4302 414 4320 432
rect 4302 432 4320 450
rect 4302 450 4320 468
rect 4302 468 4320 486
rect 4302 486 4320 504
rect 4302 504 4320 522
rect 4302 522 4320 540
rect 4302 540 4320 558
rect 4302 558 4320 576
rect 4302 576 4320 594
rect 4302 594 4320 612
rect 4302 612 4320 630
rect 4302 630 4320 648
rect 4302 648 4320 666
rect 4302 666 4320 684
rect 4302 864 4320 882
rect 4302 882 4320 900
rect 4302 900 4320 918
rect 4302 918 4320 936
rect 4302 936 4320 954
rect 4302 954 4320 972
rect 4302 972 4320 990
rect 4302 990 4320 1008
rect 4302 1008 4320 1026
rect 4302 1026 4320 1044
rect 4302 1044 4320 1062
rect 4302 1062 4320 1080
rect 4302 1080 4320 1098
rect 4302 1098 4320 1116
rect 4302 1116 4320 1134
rect 4302 1134 4320 1152
rect 4302 1152 4320 1170
rect 4302 1170 4320 1188
rect 4302 1188 4320 1206
rect 4302 1206 4320 1224
rect 4302 1224 4320 1242
rect 4302 1242 4320 1260
rect 4302 1260 4320 1278
rect 4302 1278 4320 1296
rect 4302 1296 4320 1314
rect 4302 1314 4320 1332
rect 4302 1332 4320 1350
rect 4302 1350 4320 1368
rect 4302 1368 4320 1386
rect 4302 1386 4320 1404
rect 4302 1404 4320 1422
rect 4302 1422 4320 1440
rect 4302 1440 4320 1458
rect 4302 1458 4320 1476
rect 4302 1476 4320 1494
rect 4302 1494 4320 1512
rect 4302 1512 4320 1530
rect 4302 1530 4320 1548
rect 4302 1548 4320 1566
rect 4302 1566 4320 1584
rect 4302 1584 4320 1602
rect 4302 1602 4320 1620
rect 4302 1620 4320 1638
rect 4302 1638 4320 1656
rect 4302 1656 4320 1674
rect 4302 1674 4320 1692
rect 4302 1692 4320 1710
rect 4302 1710 4320 1728
rect 4302 1728 4320 1746
rect 4302 1746 4320 1764
rect 4302 2016 4320 2034
rect 4302 2034 4320 2052
rect 4302 2052 4320 2070
rect 4302 2070 4320 2088
rect 4302 2088 4320 2106
rect 4302 2106 4320 2124
rect 4302 2124 4320 2142
rect 4302 2142 4320 2160
rect 4302 2160 4320 2178
rect 4302 2178 4320 2196
rect 4302 2196 4320 2214
rect 4302 2214 4320 2232
rect 4302 2232 4320 2250
rect 4302 2250 4320 2268
rect 4302 2268 4320 2286
rect 4302 2286 4320 2304
rect 4302 2304 4320 2322
rect 4302 2322 4320 2340
rect 4302 2340 4320 2358
rect 4302 2358 4320 2376
rect 4302 2376 4320 2394
rect 4302 2394 4320 2412
rect 4302 2412 4320 2430
rect 4302 2430 4320 2448
rect 4302 2448 4320 2466
rect 4302 2466 4320 2484
rect 4302 2484 4320 2502
rect 4302 2502 4320 2520
rect 4302 2520 4320 2538
rect 4302 2538 4320 2556
rect 4302 2556 4320 2574
rect 4302 2574 4320 2592
rect 4302 2592 4320 2610
rect 4302 2610 4320 2628
rect 4302 2628 4320 2646
rect 4302 2646 4320 2664
rect 4302 2664 4320 2682
rect 4302 2682 4320 2700
rect 4302 2700 4320 2718
rect 4302 2718 4320 2736
rect 4302 2736 4320 2754
rect 4302 2754 4320 2772
rect 4302 2772 4320 2790
rect 4302 2790 4320 2808
rect 4302 2808 4320 2826
rect 4302 2826 4320 2844
rect 4302 2844 4320 2862
rect 4302 2862 4320 2880
rect 4302 2880 4320 2898
rect 4302 2898 4320 2916
rect 4302 2916 4320 2934
rect 4302 2934 4320 2952
rect 4302 2952 4320 2970
rect 4302 2970 4320 2988
rect 4302 2988 4320 3006
rect 4302 3006 4320 3024
rect 4302 3024 4320 3042
rect 4302 3042 4320 3060
rect 4302 3060 4320 3078
rect 4302 3078 4320 3096
rect 4302 3096 4320 3114
rect 4302 3114 4320 3132
rect 4302 3132 4320 3150
rect 4302 3150 4320 3168
rect 4302 3168 4320 3186
rect 4302 3186 4320 3204
rect 4302 3204 4320 3222
rect 4302 3222 4320 3240
rect 4302 3240 4320 3258
rect 4302 3258 4320 3276
rect 4302 3276 4320 3294
rect 4302 3294 4320 3312
rect 4302 3312 4320 3330
rect 4302 3330 4320 3348
rect 4302 3348 4320 3366
rect 4302 3366 4320 3384
rect 4302 3384 4320 3402
rect 4302 3402 4320 3420
rect 4302 3420 4320 3438
rect 4302 3438 4320 3456
rect 4302 3456 4320 3474
rect 4302 3474 4320 3492
rect 4302 3492 4320 3510
rect 4302 3510 4320 3528
rect 4302 3744 4320 3762
rect 4302 3762 4320 3780
rect 4302 3780 4320 3798
rect 4302 3798 4320 3816
rect 4302 3816 4320 3834
rect 4302 3834 4320 3852
rect 4302 3852 4320 3870
rect 4302 3870 4320 3888
rect 4302 3888 4320 3906
rect 4302 3906 4320 3924
rect 4302 3924 4320 3942
rect 4302 3942 4320 3960
rect 4302 3960 4320 3978
rect 4302 3978 4320 3996
rect 4302 3996 4320 4014
rect 4302 4014 4320 4032
rect 4302 4032 4320 4050
rect 4302 4050 4320 4068
rect 4302 4068 4320 4086
rect 4302 4086 4320 4104
rect 4302 4104 4320 4122
rect 4302 4122 4320 4140
rect 4302 4140 4320 4158
rect 4302 4158 4320 4176
rect 4302 4176 4320 4194
rect 4302 4194 4320 4212
rect 4302 4212 4320 4230
rect 4302 4230 4320 4248
rect 4302 4248 4320 4266
rect 4302 4266 4320 4284
rect 4302 4284 4320 4302
rect 4302 4302 4320 4320
rect 4302 4320 4320 4338
rect 4302 4338 4320 4356
rect 4302 4356 4320 4374
rect 4302 4374 4320 4392
rect 4302 4392 4320 4410
rect 4302 4410 4320 4428
rect 4302 4428 4320 4446
rect 4302 4446 4320 4464
rect 4302 4464 4320 4482
rect 4302 4482 4320 4500
rect 4302 4500 4320 4518
rect 4302 4518 4320 4536
rect 4302 4536 4320 4554
rect 4302 4554 4320 4572
rect 4302 4572 4320 4590
rect 4302 4590 4320 4608
rect 4302 4608 4320 4626
rect 4302 4626 4320 4644
rect 4302 4644 4320 4662
rect 4302 4662 4320 4680
rect 4302 4680 4320 4698
rect 4302 4698 4320 4716
rect 4302 4716 4320 4734
rect 4302 4734 4320 4752
rect 4302 4752 4320 4770
rect 4302 4770 4320 4788
rect 4302 4788 4320 4806
rect 4302 4806 4320 4824
rect 4302 4824 4320 4842
rect 4302 4842 4320 4860
rect 4302 4860 4320 4878
rect 4302 4878 4320 4896
rect 4302 4896 4320 4914
rect 4302 4914 4320 4932
rect 4302 4932 4320 4950
rect 4302 4950 4320 4968
rect 4302 4968 4320 4986
rect 4302 4986 4320 5004
rect 4302 5004 4320 5022
rect 4302 5022 4320 5040
rect 4302 5040 4320 5058
rect 4302 5058 4320 5076
rect 4302 5076 4320 5094
rect 4302 5094 4320 5112
rect 4302 5112 4320 5130
rect 4302 5130 4320 5148
rect 4302 5148 4320 5166
rect 4302 5166 4320 5184
rect 4302 5184 4320 5202
rect 4302 5202 4320 5220
rect 4302 5220 4320 5238
rect 4302 5238 4320 5256
rect 4302 5256 4320 5274
rect 4302 5274 4320 5292
rect 4302 5292 4320 5310
rect 4302 5310 4320 5328
rect 4302 5328 4320 5346
rect 4302 5346 4320 5364
rect 4302 5364 4320 5382
rect 4302 5382 4320 5400
rect 4302 5400 4320 5418
rect 4302 5418 4320 5436
rect 4302 5436 4320 5454
rect 4302 5454 4320 5472
rect 4302 5472 4320 5490
rect 4302 5490 4320 5508
rect 4302 5508 4320 5526
rect 4302 5526 4320 5544
rect 4302 5544 4320 5562
rect 4302 5562 4320 5580
rect 4302 5580 4320 5598
rect 4302 5598 4320 5616
rect 4302 5616 4320 5634
rect 4302 5634 4320 5652
rect 4302 5652 4320 5670
rect 4302 5670 4320 5688
rect 4302 5688 4320 5706
rect 4302 5706 4320 5724
rect 4302 5724 4320 5742
rect 4302 5742 4320 5760
rect 4302 5760 4320 5778
rect 4302 5778 4320 5796
rect 4302 5796 4320 5814
rect 4302 5814 4320 5832
rect 4302 5832 4320 5850
rect 4302 5850 4320 5868
rect 4302 5868 4320 5886
rect 4302 5886 4320 5904
rect 4302 5904 4320 5922
rect 4302 5922 4320 5940
rect 4302 5940 4320 5958
rect 4302 5958 4320 5976
rect 4302 5976 4320 5994
rect 4302 5994 4320 6012
rect 4302 6012 4320 6030
rect 4302 6030 4320 6048
rect 4302 6048 4320 6066
rect 4302 6066 4320 6084
rect 4302 6084 4320 6102
rect 4302 6102 4320 6120
rect 4302 6120 4320 6138
rect 4302 6138 4320 6156
rect 4302 6156 4320 6174
rect 4302 6174 4320 6192
rect 4302 6192 4320 6210
rect 4302 6210 4320 6228
rect 4302 6228 4320 6246
rect 4302 6246 4320 6264
rect 4302 6264 4320 6282
rect 4302 6282 4320 6300
rect 4302 6300 4320 6318
rect 4302 6318 4320 6336
rect 4302 6336 4320 6354
rect 4302 6354 4320 6372
rect 4302 6372 4320 6390
rect 4302 6390 4320 6408
rect 4302 6408 4320 6426
rect 4302 6426 4320 6444
rect 4302 6444 4320 6462
rect 4302 6462 4320 6480
rect 4302 6480 4320 6498
rect 4302 6498 4320 6516
rect 4302 6516 4320 6534
rect 4302 6534 4320 6552
rect 4302 6552 4320 6570
rect 4302 6570 4320 6588
rect 4302 6588 4320 6606
rect 4302 6606 4320 6624
rect 4302 6624 4320 6642
rect 4302 6642 4320 6660
rect 4302 6660 4320 6678
rect 4302 6678 4320 6696
rect 4302 7020 4320 7038
rect 4302 7038 4320 7056
rect 4302 7056 4320 7074
rect 4302 7074 4320 7092
rect 4302 7092 4320 7110
rect 4302 7110 4320 7128
rect 4302 7128 4320 7146
rect 4302 7146 4320 7164
rect 4302 7164 4320 7182
rect 4302 7182 4320 7200
rect 4302 7200 4320 7218
rect 4320 54 4338 72
rect 4320 72 4338 90
rect 4320 90 4338 108
rect 4320 108 4338 126
rect 4320 126 4338 144
rect 4320 144 4338 162
rect 4320 162 4338 180
rect 4320 180 4338 198
rect 4320 198 4338 216
rect 4320 216 4338 234
rect 4320 234 4338 252
rect 4320 252 4338 270
rect 4320 270 4338 288
rect 4320 288 4338 306
rect 4320 306 4338 324
rect 4320 324 4338 342
rect 4320 342 4338 360
rect 4320 360 4338 378
rect 4320 378 4338 396
rect 4320 396 4338 414
rect 4320 414 4338 432
rect 4320 432 4338 450
rect 4320 450 4338 468
rect 4320 468 4338 486
rect 4320 486 4338 504
rect 4320 504 4338 522
rect 4320 522 4338 540
rect 4320 540 4338 558
rect 4320 558 4338 576
rect 4320 576 4338 594
rect 4320 594 4338 612
rect 4320 612 4338 630
rect 4320 630 4338 648
rect 4320 648 4338 666
rect 4320 666 4338 684
rect 4320 684 4338 702
rect 4320 864 4338 882
rect 4320 882 4338 900
rect 4320 900 4338 918
rect 4320 918 4338 936
rect 4320 936 4338 954
rect 4320 954 4338 972
rect 4320 972 4338 990
rect 4320 990 4338 1008
rect 4320 1008 4338 1026
rect 4320 1026 4338 1044
rect 4320 1044 4338 1062
rect 4320 1062 4338 1080
rect 4320 1080 4338 1098
rect 4320 1098 4338 1116
rect 4320 1116 4338 1134
rect 4320 1134 4338 1152
rect 4320 1152 4338 1170
rect 4320 1170 4338 1188
rect 4320 1188 4338 1206
rect 4320 1206 4338 1224
rect 4320 1224 4338 1242
rect 4320 1242 4338 1260
rect 4320 1260 4338 1278
rect 4320 1278 4338 1296
rect 4320 1296 4338 1314
rect 4320 1314 4338 1332
rect 4320 1332 4338 1350
rect 4320 1350 4338 1368
rect 4320 1368 4338 1386
rect 4320 1386 4338 1404
rect 4320 1404 4338 1422
rect 4320 1422 4338 1440
rect 4320 1440 4338 1458
rect 4320 1458 4338 1476
rect 4320 1476 4338 1494
rect 4320 1494 4338 1512
rect 4320 1512 4338 1530
rect 4320 1530 4338 1548
rect 4320 1548 4338 1566
rect 4320 1566 4338 1584
rect 4320 1584 4338 1602
rect 4320 1602 4338 1620
rect 4320 1620 4338 1638
rect 4320 1638 4338 1656
rect 4320 1656 4338 1674
rect 4320 1674 4338 1692
rect 4320 1692 4338 1710
rect 4320 1710 4338 1728
rect 4320 1728 4338 1746
rect 4320 1746 4338 1764
rect 4320 1764 4338 1782
rect 4320 2016 4338 2034
rect 4320 2034 4338 2052
rect 4320 2052 4338 2070
rect 4320 2070 4338 2088
rect 4320 2088 4338 2106
rect 4320 2106 4338 2124
rect 4320 2124 4338 2142
rect 4320 2142 4338 2160
rect 4320 2160 4338 2178
rect 4320 2178 4338 2196
rect 4320 2196 4338 2214
rect 4320 2214 4338 2232
rect 4320 2232 4338 2250
rect 4320 2250 4338 2268
rect 4320 2268 4338 2286
rect 4320 2286 4338 2304
rect 4320 2304 4338 2322
rect 4320 2322 4338 2340
rect 4320 2340 4338 2358
rect 4320 2358 4338 2376
rect 4320 2376 4338 2394
rect 4320 2394 4338 2412
rect 4320 2412 4338 2430
rect 4320 2430 4338 2448
rect 4320 2448 4338 2466
rect 4320 2466 4338 2484
rect 4320 2484 4338 2502
rect 4320 2502 4338 2520
rect 4320 2520 4338 2538
rect 4320 2538 4338 2556
rect 4320 2556 4338 2574
rect 4320 2574 4338 2592
rect 4320 2592 4338 2610
rect 4320 2610 4338 2628
rect 4320 2628 4338 2646
rect 4320 2646 4338 2664
rect 4320 2664 4338 2682
rect 4320 2682 4338 2700
rect 4320 2700 4338 2718
rect 4320 2718 4338 2736
rect 4320 2736 4338 2754
rect 4320 2754 4338 2772
rect 4320 2772 4338 2790
rect 4320 2790 4338 2808
rect 4320 2808 4338 2826
rect 4320 2826 4338 2844
rect 4320 2844 4338 2862
rect 4320 2862 4338 2880
rect 4320 2880 4338 2898
rect 4320 2898 4338 2916
rect 4320 2916 4338 2934
rect 4320 2934 4338 2952
rect 4320 2952 4338 2970
rect 4320 2970 4338 2988
rect 4320 2988 4338 3006
rect 4320 3006 4338 3024
rect 4320 3024 4338 3042
rect 4320 3042 4338 3060
rect 4320 3060 4338 3078
rect 4320 3078 4338 3096
rect 4320 3096 4338 3114
rect 4320 3114 4338 3132
rect 4320 3132 4338 3150
rect 4320 3150 4338 3168
rect 4320 3168 4338 3186
rect 4320 3186 4338 3204
rect 4320 3204 4338 3222
rect 4320 3222 4338 3240
rect 4320 3240 4338 3258
rect 4320 3258 4338 3276
rect 4320 3276 4338 3294
rect 4320 3294 4338 3312
rect 4320 3312 4338 3330
rect 4320 3330 4338 3348
rect 4320 3348 4338 3366
rect 4320 3366 4338 3384
rect 4320 3384 4338 3402
rect 4320 3402 4338 3420
rect 4320 3420 4338 3438
rect 4320 3438 4338 3456
rect 4320 3456 4338 3474
rect 4320 3474 4338 3492
rect 4320 3492 4338 3510
rect 4320 3510 4338 3528
rect 4320 3528 4338 3546
rect 4320 3762 4338 3780
rect 4320 3780 4338 3798
rect 4320 3798 4338 3816
rect 4320 3816 4338 3834
rect 4320 3834 4338 3852
rect 4320 3852 4338 3870
rect 4320 3870 4338 3888
rect 4320 3888 4338 3906
rect 4320 3906 4338 3924
rect 4320 3924 4338 3942
rect 4320 3942 4338 3960
rect 4320 3960 4338 3978
rect 4320 3978 4338 3996
rect 4320 3996 4338 4014
rect 4320 4014 4338 4032
rect 4320 4032 4338 4050
rect 4320 4050 4338 4068
rect 4320 4068 4338 4086
rect 4320 4086 4338 4104
rect 4320 4104 4338 4122
rect 4320 4122 4338 4140
rect 4320 4140 4338 4158
rect 4320 4158 4338 4176
rect 4320 4176 4338 4194
rect 4320 4194 4338 4212
rect 4320 4212 4338 4230
rect 4320 4230 4338 4248
rect 4320 4248 4338 4266
rect 4320 4266 4338 4284
rect 4320 4284 4338 4302
rect 4320 4302 4338 4320
rect 4320 4320 4338 4338
rect 4320 4338 4338 4356
rect 4320 4356 4338 4374
rect 4320 4374 4338 4392
rect 4320 4392 4338 4410
rect 4320 4410 4338 4428
rect 4320 4428 4338 4446
rect 4320 4446 4338 4464
rect 4320 4464 4338 4482
rect 4320 4482 4338 4500
rect 4320 4500 4338 4518
rect 4320 4518 4338 4536
rect 4320 4536 4338 4554
rect 4320 4554 4338 4572
rect 4320 4572 4338 4590
rect 4320 4590 4338 4608
rect 4320 4608 4338 4626
rect 4320 4626 4338 4644
rect 4320 4644 4338 4662
rect 4320 4662 4338 4680
rect 4320 4680 4338 4698
rect 4320 4698 4338 4716
rect 4320 4716 4338 4734
rect 4320 4734 4338 4752
rect 4320 4752 4338 4770
rect 4320 4770 4338 4788
rect 4320 4788 4338 4806
rect 4320 4806 4338 4824
rect 4320 4824 4338 4842
rect 4320 4842 4338 4860
rect 4320 4860 4338 4878
rect 4320 4878 4338 4896
rect 4320 4896 4338 4914
rect 4320 4914 4338 4932
rect 4320 4932 4338 4950
rect 4320 4950 4338 4968
rect 4320 4968 4338 4986
rect 4320 4986 4338 5004
rect 4320 5004 4338 5022
rect 4320 5022 4338 5040
rect 4320 5040 4338 5058
rect 4320 5058 4338 5076
rect 4320 5076 4338 5094
rect 4320 5094 4338 5112
rect 4320 5112 4338 5130
rect 4320 5130 4338 5148
rect 4320 5148 4338 5166
rect 4320 5166 4338 5184
rect 4320 5184 4338 5202
rect 4320 5202 4338 5220
rect 4320 5220 4338 5238
rect 4320 5238 4338 5256
rect 4320 5256 4338 5274
rect 4320 5274 4338 5292
rect 4320 5292 4338 5310
rect 4320 5310 4338 5328
rect 4320 5328 4338 5346
rect 4320 5346 4338 5364
rect 4320 5364 4338 5382
rect 4320 5382 4338 5400
rect 4320 5400 4338 5418
rect 4320 5418 4338 5436
rect 4320 5436 4338 5454
rect 4320 5454 4338 5472
rect 4320 5472 4338 5490
rect 4320 5490 4338 5508
rect 4320 5508 4338 5526
rect 4320 5526 4338 5544
rect 4320 5544 4338 5562
rect 4320 5562 4338 5580
rect 4320 5580 4338 5598
rect 4320 5598 4338 5616
rect 4320 5616 4338 5634
rect 4320 5634 4338 5652
rect 4320 5652 4338 5670
rect 4320 5670 4338 5688
rect 4320 5688 4338 5706
rect 4320 5706 4338 5724
rect 4320 5724 4338 5742
rect 4320 5742 4338 5760
rect 4320 5760 4338 5778
rect 4320 5778 4338 5796
rect 4320 5796 4338 5814
rect 4320 5814 4338 5832
rect 4320 5832 4338 5850
rect 4320 5850 4338 5868
rect 4320 5868 4338 5886
rect 4320 5886 4338 5904
rect 4320 5904 4338 5922
rect 4320 5922 4338 5940
rect 4320 5940 4338 5958
rect 4320 5958 4338 5976
rect 4320 5976 4338 5994
rect 4320 5994 4338 6012
rect 4320 6012 4338 6030
rect 4320 6030 4338 6048
rect 4320 6048 4338 6066
rect 4320 6066 4338 6084
rect 4320 6084 4338 6102
rect 4320 6102 4338 6120
rect 4320 6120 4338 6138
rect 4320 6138 4338 6156
rect 4320 6156 4338 6174
rect 4320 6174 4338 6192
rect 4320 6192 4338 6210
rect 4320 6210 4338 6228
rect 4320 6228 4338 6246
rect 4320 6246 4338 6264
rect 4320 6264 4338 6282
rect 4320 6282 4338 6300
rect 4320 6300 4338 6318
rect 4320 6318 4338 6336
rect 4320 6336 4338 6354
rect 4320 6354 4338 6372
rect 4320 6372 4338 6390
rect 4320 6390 4338 6408
rect 4320 6408 4338 6426
rect 4320 6426 4338 6444
rect 4320 6444 4338 6462
rect 4320 6462 4338 6480
rect 4320 6480 4338 6498
rect 4320 6498 4338 6516
rect 4320 6516 4338 6534
rect 4320 6534 4338 6552
rect 4320 6552 4338 6570
rect 4320 6570 4338 6588
rect 4320 6588 4338 6606
rect 4320 6606 4338 6624
rect 4320 6624 4338 6642
rect 4320 6642 4338 6660
rect 4320 6660 4338 6678
rect 4320 6678 4338 6696
rect 4320 6696 4338 6714
rect 4320 7056 4338 7074
rect 4320 7074 4338 7092
rect 4320 7092 4338 7110
rect 4320 7110 4338 7128
rect 4320 7128 4338 7146
rect 4320 7146 4338 7164
rect 4320 7164 4338 7182
rect 4320 7182 4338 7200
rect 4320 7200 4338 7218
rect 4338 72 4356 90
rect 4338 90 4356 108
rect 4338 108 4356 126
rect 4338 126 4356 144
rect 4338 144 4356 162
rect 4338 162 4356 180
rect 4338 180 4356 198
rect 4338 198 4356 216
rect 4338 216 4356 234
rect 4338 234 4356 252
rect 4338 252 4356 270
rect 4338 270 4356 288
rect 4338 288 4356 306
rect 4338 306 4356 324
rect 4338 324 4356 342
rect 4338 342 4356 360
rect 4338 360 4356 378
rect 4338 378 4356 396
rect 4338 396 4356 414
rect 4338 414 4356 432
rect 4338 432 4356 450
rect 4338 450 4356 468
rect 4338 468 4356 486
rect 4338 486 4356 504
rect 4338 504 4356 522
rect 4338 522 4356 540
rect 4338 540 4356 558
rect 4338 558 4356 576
rect 4338 576 4356 594
rect 4338 594 4356 612
rect 4338 612 4356 630
rect 4338 630 4356 648
rect 4338 648 4356 666
rect 4338 666 4356 684
rect 4338 684 4356 702
rect 4338 864 4356 882
rect 4338 882 4356 900
rect 4338 900 4356 918
rect 4338 918 4356 936
rect 4338 936 4356 954
rect 4338 954 4356 972
rect 4338 972 4356 990
rect 4338 990 4356 1008
rect 4338 1008 4356 1026
rect 4338 1026 4356 1044
rect 4338 1044 4356 1062
rect 4338 1062 4356 1080
rect 4338 1080 4356 1098
rect 4338 1098 4356 1116
rect 4338 1116 4356 1134
rect 4338 1134 4356 1152
rect 4338 1152 4356 1170
rect 4338 1170 4356 1188
rect 4338 1188 4356 1206
rect 4338 1206 4356 1224
rect 4338 1224 4356 1242
rect 4338 1242 4356 1260
rect 4338 1260 4356 1278
rect 4338 1278 4356 1296
rect 4338 1296 4356 1314
rect 4338 1314 4356 1332
rect 4338 1332 4356 1350
rect 4338 1350 4356 1368
rect 4338 1368 4356 1386
rect 4338 1386 4356 1404
rect 4338 1404 4356 1422
rect 4338 1422 4356 1440
rect 4338 1440 4356 1458
rect 4338 1458 4356 1476
rect 4338 1476 4356 1494
rect 4338 1494 4356 1512
rect 4338 1512 4356 1530
rect 4338 1530 4356 1548
rect 4338 1548 4356 1566
rect 4338 1566 4356 1584
rect 4338 1584 4356 1602
rect 4338 1602 4356 1620
rect 4338 1620 4356 1638
rect 4338 1638 4356 1656
rect 4338 1656 4356 1674
rect 4338 1674 4356 1692
rect 4338 1692 4356 1710
rect 4338 1710 4356 1728
rect 4338 1728 4356 1746
rect 4338 1746 4356 1764
rect 4338 1764 4356 1782
rect 4338 1782 4356 1800
rect 4338 2034 4356 2052
rect 4338 2052 4356 2070
rect 4338 2070 4356 2088
rect 4338 2088 4356 2106
rect 4338 2106 4356 2124
rect 4338 2124 4356 2142
rect 4338 2142 4356 2160
rect 4338 2160 4356 2178
rect 4338 2178 4356 2196
rect 4338 2196 4356 2214
rect 4338 2214 4356 2232
rect 4338 2232 4356 2250
rect 4338 2250 4356 2268
rect 4338 2268 4356 2286
rect 4338 2286 4356 2304
rect 4338 2304 4356 2322
rect 4338 2322 4356 2340
rect 4338 2340 4356 2358
rect 4338 2358 4356 2376
rect 4338 2376 4356 2394
rect 4338 2394 4356 2412
rect 4338 2412 4356 2430
rect 4338 2430 4356 2448
rect 4338 2448 4356 2466
rect 4338 2466 4356 2484
rect 4338 2484 4356 2502
rect 4338 2502 4356 2520
rect 4338 2520 4356 2538
rect 4338 2538 4356 2556
rect 4338 2556 4356 2574
rect 4338 2574 4356 2592
rect 4338 2592 4356 2610
rect 4338 2610 4356 2628
rect 4338 2628 4356 2646
rect 4338 2646 4356 2664
rect 4338 2664 4356 2682
rect 4338 2682 4356 2700
rect 4338 2700 4356 2718
rect 4338 2718 4356 2736
rect 4338 2736 4356 2754
rect 4338 2754 4356 2772
rect 4338 2772 4356 2790
rect 4338 2790 4356 2808
rect 4338 2808 4356 2826
rect 4338 2826 4356 2844
rect 4338 2844 4356 2862
rect 4338 2862 4356 2880
rect 4338 2880 4356 2898
rect 4338 2898 4356 2916
rect 4338 2916 4356 2934
rect 4338 2934 4356 2952
rect 4338 2952 4356 2970
rect 4338 2970 4356 2988
rect 4338 2988 4356 3006
rect 4338 3006 4356 3024
rect 4338 3024 4356 3042
rect 4338 3042 4356 3060
rect 4338 3060 4356 3078
rect 4338 3078 4356 3096
rect 4338 3096 4356 3114
rect 4338 3114 4356 3132
rect 4338 3132 4356 3150
rect 4338 3150 4356 3168
rect 4338 3168 4356 3186
rect 4338 3186 4356 3204
rect 4338 3204 4356 3222
rect 4338 3222 4356 3240
rect 4338 3240 4356 3258
rect 4338 3258 4356 3276
rect 4338 3276 4356 3294
rect 4338 3294 4356 3312
rect 4338 3312 4356 3330
rect 4338 3330 4356 3348
rect 4338 3348 4356 3366
rect 4338 3366 4356 3384
rect 4338 3384 4356 3402
rect 4338 3402 4356 3420
rect 4338 3420 4356 3438
rect 4338 3438 4356 3456
rect 4338 3456 4356 3474
rect 4338 3474 4356 3492
rect 4338 3492 4356 3510
rect 4338 3510 4356 3528
rect 4338 3528 4356 3546
rect 4338 3546 4356 3564
rect 4338 3564 4356 3582
rect 4338 3780 4356 3798
rect 4338 3798 4356 3816
rect 4338 3816 4356 3834
rect 4338 3834 4356 3852
rect 4338 3852 4356 3870
rect 4338 3870 4356 3888
rect 4338 3888 4356 3906
rect 4338 3906 4356 3924
rect 4338 3924 4356 3942
rect 4338 3942 4356 3960
rect 4338 3960 4356 3978
rect 4338 3978 4356 3996
rect 4338 3996 4356 4014
rect 4338 4014 4356 4032
rect 4338 4032 4356 4050
rect 4338 4050 4356 4068
rect 4338 4068 4356 4086
rect 4338 4086 4356 4104
rect 4338 4104 4356 4122
rect 4338 4122 4356 4140
rect 4338 4140 4356 4158
rect 4338 4158 4356 4176
rect 4338 4176 4356 4194
rect 4338 4194 4356 4212
rect 4338 4212 4356 4230
rect 4338 4230 4356 4248
rect 4338 4248 4356 4266
rect 4338 4266 4356 4284
rect 4338 4284 4356 4302
rect 4338 4302 4356 4320
rect 4338 4320 4356 4338
rect 4338 4338 4356 4356
rect 4338 4356 4356 4374
rect 4338 4374 4356 4392
rect 4338 4392 4356 4410
rect 4338 4410 4356 4428
rect 4338 4428 4356 4446
rect 4338 4446 4356 4464
rect 4338 4464 4356 4482
rect 4338 4482 4356 4500
rect 4338 4500 4356 4518
rect 4338 4518 4356 4536
rect 4338 4536 4356 4554
rect 4338 4554 4356 4572
rect 4338 4572 4356 4590
rect 4338 4590 4356 4608
rect 4338 4608 4356 4626
rect 4338 4626 4356 4644
rect 4338 4644 4356 4662
rect 4338 4662 4356 4680
rect 4338 4680 4356 4698
rect 4338 4698 4356 4716
rect 4338 4716 4356 4734
rect 4338 4734 4356 4752
rect 4338 4752 4356 4770
rect 4338 4770 4356 4788
rect 4338 4788 4356 4806
rect 4338 4806 4356 4824
rect 4338 4824 4356 4842
rect 4338 4842 4356 4860
rect 4338 4860 4356 4878
rect 4338 4878 4356 4896
rect 4338 4896 4356 4914
rect 4338 4914 4356 4932
rect 4338 4932 4356 4950
rect 4338 4950 4356 4968
rect 4338 4968 4356 4986
rect 4338 4986 4356 5004
rect 4338 5004 4356 5022
rect 4338 5022 4356 5040
rect 4338 5040 4356 5058
rect 4338 5058 4356 5076
rect 4338 5076 4356 5094
rect 4338 5094 4356 5112
rect 4338 5112 4356 5130
rect 4338 5130 4356 5148
rect 4338 5148 4356 5166
rect 4338 5166 4356 5184
rect 4338 5184 4356 5202
rect 4338 5202 4356 5220
rect 4338 5220 4356 5238
rect 4338 5238 4356 5256
rect 4338 5256 4356 5274
rect 4338 5274 4356 5292
rect 4338 5292 4356 5310
rect 4338 5310 4356 5328
rect 4338 5328 4356 5346
rect 4338 5346 4356 5364
rect 4338 5364 4356 5382
rect 4338 5382 4356 5400
rect 4338 5400 4356 5418
rect 4338 5418 4356 5436
rect 4338 5436 4356 5454
rect 4338 5454 4356 5472
rect 4338 5472 4356 5490
rect 4338 5490 4356 5508
rect 4338 5508 4356 5526
rect 4338 5526 4356 5544
rect 4338 5544 4356 5562
rect 4338 5562 4356 5580
rect 4338 5580 4356 5598
rect 4338 5598 4356 5616
rect 4338 5616 4356 5634
rect 4338 5634 4356 5652
rect 4338 5652 4356 5670
rect 4338 5670 4356 5688
rect 4338 5688 4356 5706
rect 4338 5706 4356 5724
rect 4338 5724 4356 5742
rect 4338 5742 4356 5760
rect 4338 5760 4356 5778
rect 4338 5778 4356 5796
rect 4338 5796 4356 5814
rect 4338 5814 4356 5832
rect 4338 5832 4356 5850
rect 4338 5850 4356 5868
rect 4338 5868 4356 5886
rect 4338 5886 4356 5904
rect 4338 5904 4356 5922
rect 4338 5922 4356 5940
rect 4338 5940 4356 5958
rect 4338 5958 4356 5976
rect 4338 5976 4356 5994
rect 4338 5994 4356 6012
rect 4338 6012 4356 6030
rect 4338 6030 4356 6048
rect 4338 6048 4356 6066
rect 4338 6066 4356 6084
rect 4338 6084 4356 6102
rect 4338 6102 4356 6120
rect 4338 6120 4356 6138
rect 4338 6138 4356 6156
rect 4338 6156 4356 6174
rect 4338 6174 4356 6192
rect 4338 6192 4356 6210
rect 4338 6210 4356 6228
rect 4338 6228 4356 6246
rect 4338 6246 4356 6264
rect 4338 6264 4356 6282
rect 4338 6282 4356 6300
rect 4338 6300 4356 6318
rect 4338 6318 4356 6336
rect 4338 6336 4356 6354
rect 4338 6354 4356 6372
rect 4338 6372 4356 6390
rect 4338 6390 4356 6408
rect 4338 6408 4356 6426
rect 4338 6426 4356 6444
rect 4338 6444 4356 6462
rect 4338 6462 4356 6480
rect 4338 6480 4356 6498
rect 4338 6498 4356 6516
rect 4338 6516 4356 6534
rect 4338 6534 4356 6552
rect 4338 6552 4356 6570
rect 4338 6570 4356 6588
rect 4338 6588 4356 6606
rect 4338 6606 4356 6624
rect 4338 6624 4356 6642
rect 4338 6642 4356 6660
rect 4338 6660 4356 6678
rect 4338 6678 4356 6696
rect 4338 6696 4356 6714
rect 4338 6714 4356 6732
rect 4338 6732 4356 6750
rect 4338 7074 4356 7092
rect 4338 7092 4356 7110
rect 4338 7110 4356 7128
rect 4338 7128 4356 7146
rect 4338 7146 4356 7164
rect 4338 7164 4356 7182
rect 4338 7182 4356 7200
rect 4338 7200 4356 7218
rect 4356 72 4374 90
rect 4356 90 4374 108
rect 4356 108 4374 126
rect 4356 126 4374 144
rect 4356 144 4374 162
rect 4356 162 4374 180
rect 4356 180 4374 198
rect 4356 198 4374 216
rect 4356 216 4374 234
rect 4356 234 4374 252
rect 4356 252 4374 270
rect 4356 270 4374 288
rect 4356 288 4374 306
rect 4356 306 4374 324
rect 4356 324 4374 342
rect 4356 342 4374 360
rect 4356 360 4374 378
rect 4356 378 4374 396
rect 4356 396 4374 414
rect 4356 414 4374 432
rect 4356 432 4374 450
rect 4356 450 4374 468
rect 4356 468 4374 486
rect 4356 486 4374 504
rect 4356 504 4374 522
rect 4356 522 4374 540
rect 4356 540 4374 558
rect 4356 558 4374 576
rect 4356 576 4374 594
rect 4356 594 4374 612
rect 4356 612 4374 630
rect 4356 630 4374 648
rect 4356 648 4374 666
rect 4356 666 4374 684
rect 4356 684 4374 702
rect 4356 864 4374 882
rect 4356 882 4374 900
rect 4356 900 4374 918
rect 4356 918 4374 936
rect 4356 936 4374 954
rect 4356 954 4374 972
rect 4356 972 4374 990
rect 4356 990 4374 1008
rect 4356 1008 4374 1026
rect 4356 1026 4374 1044
rect 4356 1044 4374 1062
rect 4356 1062 4374 1080
rect 4356 1080 4374 1098
rect 4356 1098 4374 1116
rect 4356 1116 4374 1134
rect 4356 1134 4374 1152
rect 4356 1152 4374 1170
rect 4356 1170 4374 1188
rect 4356 1188 4374 1206
rect 4356 1206 4374 1224
rect 4356 1224 4374 1242
rect 4356 1242 4374 1260
rect 4356 1260 4374 1278
rect 4356 1278 4374 1296
rect 4356 1296 4374 1314
rect 4356 1314 4374 1332
rect 4356 1332 4374 1350
rect 4356 1350 4374 1368
rect 4356 1368 4374 1386
rect 4356 1386 4374 1404
rect 4356 1404 4374 1422
rect 4356 1422 4374 1440
rect 4356 1440 4374 1458
rect 4356 1458 4374 1476
rect 4356 1476 4374 1494
rect 4356 1494 4374 1512
rect 4356 1512 4374 1530
rect 4356 1530 4374 1548
rect 4356 1548 4374 1566
rect 4356 1566 4374 1584
rect 4356 1584 4374 1602
rect 4356 1602 4374 1620
rect 4356 1620 4374 1638
rect 4356 1638 4374 1656
rect 4356 1656 4374 1674
rect 4356 1674 4374 1692
rect 4356 1692 4374 1710
rect 4356 1710 4374 1728
rect 4356 1728 4374 1746
rect 4356 1746 4374 1764
rect 4356 1764 4374 1782
rect 4356 1782 4374 1800
rect 4356 2052 4374 2070
rect 4356 2070 4374 2088
rect 4356 2088 4374 2106
rect 4356 2106 4374 2124
rect 4356 2124 4374 2142
rect 4356 2142 4374 2160
rect 4356 2160 4374 2178
rect 4356 2178 4374 2196
rect 4356 2196 4374 2214
rect 4356 2214 4374 2232
rect 4356 2232 4374 2250
rect 4356 2250 4374 2268
rect 4356 2268 4374 2286
rect 4356 2286 4374 2304
rect 4356 2304 4374 2322
rect 4356 2322 4374 2340
rect 4356 2340 4374 2358
rect 4356 2358 4374 2376
rect 4356 2376 4374 2394
rect 4356 2394 4374 2412
rect 4356 2412 4374 2430
rect 4356 2430 4374 2448
rect 4356 2448 4374 2466
rect 4356 2466 4374 2484
rect 4356 2484 4374 2502
rect 4356 2502 4374 2520
rect 4356 2520 4374 2538
rect 4356 2538 4374 2556
rect 4356 2556 4374 2574
rect 4356 2574 4374 2592
rect 4356 2592 4374 2610
rect 4356 2610 4374 2628
rect 4356 2628 4374 2646
rect 4356 2646 4374 2664
rect 4356 2664 4374 2682
rect 4356 2682 4374 2700
rect 4356 2700 4374 2718
rect 4356 2718 4374 2736
rect 4356 2736 4374 2754
rect 4356 2754 4374 2772
rect 4356 2772 4374 2790
rect 4356 2790 4374 2808
rect 4356 2808 4374 2826
rect 4356 2826 4374 2844
rect 4356 2844 4374 2862
rect 4356 2862 4374 2880
rect 4356 2880 4374 2898
rect 4356 2898 4374 2916
rect 4356 2916 4374 2934
rect 4356 2934 4374 2952
rect 4356 2952 4374 2970
rect 4356 2970 4374 2988
rect 4356 2988 4374 3006
rect 4356 3006 4374 3024
rect 4356 3024 4374 3042
rect 4356 3042 4374 3060
rect 4356 3060 4374 3078
rect 4356 3078 4374 3096
rect 4356 3096 4374 3114
rect 4356 3114 4374 3132
rect 4356 3132 4374 3150
rect 4356 3150 4374 3168
rect 4356 3168 4374 3186
rect 4356 3186 4374 3204
rect 4356 3204 4374 3222
rect 4356 3222 4374 3240
rect 4356 3240 4374 3258
rect 4356 3258 4374 3276
rect 4356 3276 4374 3294
rect 4356 3294 4374 3312
rect 4356 3312 4374 3330
rect 4356 3330 4374 3348
rect 4356 3348 4374 3366
rect 4356 3366 4374 3384
rect 4356 3384 4374 3402
rect 4356 3402 4374 3420
rect 4356 3420 4374 3438
rect 4356 3438 4374 3456
rect 4356 3456 4374 3474
rect 4356 3474 4374 3492
rect 4356 3492 4374 3510
rect 4356 3510 4374 3528
rect 4356 3528 4374 3546
rect 4356 3546 4374 3564
rect 4356 3564 4374 3582
rect 4356 3582 4374 3600
rect 4356 3816 4374 3834
rect 4356 3834 4374 3852
rect 4356 3852 4374 3870
rect 4356 3870 4374 3888
rect 4356 3888 4374 3906
rect 4356 3906 4374 3924
rect 4356 3924 4374 3942
rect 4356 3942 4374 3960
rect 4356 3960 4374 3978
rect 4356 3978 4374 3996
rect 4356 3996 4374 4014
rect 4356 4014 4374 4032
rect 4356 4032 4374 4050
rect 4356 4050 4374 4068
rect 4356 4068 4374 4086
rect 4356 4086 4374 4104
rect 4356 4104 4374 4122
rect 4356 4122 4374 4140
rect 4356 4140 4374 4158
rect 4356 4158 4374 4176
rect 4356 4176 4374 4194
rect 4356 4194 4374 4212
rect 4356 4212 4374 4230
rect 4356 4230 4374 4248
rect 4356 4248 4374 4266
rect 4356 4266 4374 4284
rect 4356 4284 4374 4302
rect 4356 4302 4374 4320
rect 4356 4320 4374 4338
rect 4356 4338 4374 4356
rect 4356 4356 4374 4374
rect 4356 4374 4374 4392
rect 4356 4392 4374 4410
rect 4356 4410 4374 4428
rect 4356 4428 4374 4446
rect 4356 4446 4374 4464
rect 4356 4464 4374 4482
rect 4356 4482 4374 4500
rect 4356 4500 4374 4518
rect 4356 4518 4374 4536
rect 4356 4536 4374 4554
rect 4356 4554 4374 4572
rect 4356 4572 4374 4590
rect 4356 4590 4374 4608
rect 4356 4608 4374 4626
rect 4356 4626 4374 4644
rect 4356 4644 4374 4662
rect 4356 4662 4374 4680
rect 4356 4680 4374 4698
rect 4356 4698 4374 4716
rect 4356 4716 4374 4734
rect 4356 4734 4374 4752
rect 4356 4752 4374 4770
rect 4356 4770 4374 4788
rect 4356 4788 4374 4806
rect 4356 4806 4374 4824
rect 4356 4824 4374 4842
rect 4356 4842 4374 4860
rect 4356 4860 4374 4878
rect 4356 4878 4374 4896
rect 4356 4896 4374 4914
rect 4356 4914 4374 4932
rect 4356 4932 4374 4950
rect 4356 4950 4374 4968
rect 4356 4968 4374 4986
rect 4356 4986 4374 5004
rect 4356 5004 4374 5022
rect 4356 5022 4374 5040
rect 4356 5040 4374 5058
rect 4356 5058 4374 5076
rect 4356 5076 4374 5094
rect 4356 5094 4374 5112
rect 4356 5112 4374 5130
rect 4356 5130 4374 5148
rect 4356 5148 4374 5166
rect 4356 5166 4374 5184
rect 4356 5184 4374 5202
rect 4356 5202 4374 5220
rect 4356 5220 4374 5238
rect 4356 5238 4374 5256
rect 4356 5256 4374 5274
rect 4356 5274 4374 5292
rect 4356 5292 4374 5310
rect 4356 5310 4374 5328
rect 4356 5328 4374 5346
rect 4356 5346 4374 5364
rect 4356 5364 4374 5382
rect 4356 5382 4374 5400
rect 4356 5400 4374 5418
rect 4356 5418 4374 5436
rect 4356 5436 4374 5454
rect 4356 5454 4374 5472
rect 4356 5472 4374 5490
rect 4356 5490 4374 5508
rect 4356 5508 4374 5526
rect 4356 5526 4374 5544
rect 4356 5544 4374 5562
rect 4356 5562 4374 5580
rect 4356 5580 4374 5598
rect 4356 5598 4374 5616
rect 4356 5616 4374 5634
rect 4356 5634 4374 5652
rect 4356 5652 4374 5670
rect 4356 5670 4374 5688
rect 4356 5688 4374 5706
rect 4356 5706 4374 5724
rect 4356 5724 4374 5742
rect 4356 5742 4374 5760
rect 4356 5760 4374 5778
rect 4356 5778 4374 5796
rect 4356 5796 4374 5814
rect 4356 5814 4374 5832
rect 4356 5832 4374 5850
rect 4356 5850 4374 5868
rect 4356 5868 4374 5886
rect 4356 5886 4374 5904
rect 4356 5904 4374 5922
rect 4356 5922 4374 5940
rect 4356 5940 4374 5958
rect 4356 5958 4374 5976
rect 4356 5976 4374 5994
rect 4356 5994 4374 6012
rect 4356 6012 4374 6030
rect 4356 6030 4374 6048
rect 4356 6048 4374 6066
rect 4356 6066 4374 6084
rect 4356 6084 4374 6102
rect 4356 6102 4374 6120
rect 4356 6120 4374 6138
rect 4356 6138 4374 6156
rect 4356 6156 4374 6174
rect 4356 6174 4374 6192
rect 4356 6192 4374 6210
rect 4356 6210 4374 6228
rect 4356 6228 4374 6246
rect 4356 6246 4374 6264
rect 4356 6264 4374 6282
rect 4356 6282 4374 6300
rect 4356 6300 4374 6318
rect 4356 6318 4374 6336
rect 4356 6336 4374 6354
rect 4356 6354 4374 6372
rect 4356 6372 4374 6390
rect 4356 6390 4374 6408
rect 4356 6408 4374 6426
rect 4356 6426 4374 6444
rect 4356 6444 4374 6462
rect 4356 6462 4374 6480
rect 4356 6480 4374 6498
rect 4356 6498 4374 6516
rect 4356 6516 4374 6534
rect 4356 6534 4374 6552
rect 4356 6552 4374 6570
rect 4356 6570 4374 6588
rect 4356 6588 4374 6606
rect 4356 6606 4374 6624
rect 4356 6624 4374 6642
rect 4356 6642 4374 6660
rect 4356 6660 4374 6678
rect 4356 6678 4374 6696
rect 4356 6696 4374 6714
rect 4356 6714 4374 6732
rect 4356 6732 4374 6750
rect 4356 6750 4374 6768
rect 4356 6768 4374 6786
rect 4356 7110 4374 7128
rect 4356 7128 4374 7146
rect 4356 7146 4374 7164
rect 4356 7164 4374 7182
rect 4356 7182 4374 7200
rect 4356 7200 4374 7218
rect 4374 72 4392 90
rect 4374 90 4392 108
rect 4374 108 4392 126
rect 4374 126 4392 144
rect 4374 144 4392 162
rect 4374 162 4392 180
rect 4374 180 4392 198
rect 4374 198 4392 216
rect 4374 216 4392 234
rect 4374 234 4392 252
rect 4374 252 4392 270
rect 4374 270 4392 288
rect 4374 288 4392 306
rect 4374 306 4392 324
rect 4374 324 4392 342
rect 4374 342 4392 360
rect 4374 360 4392 378
rect 4374 378 4392 396
rect 4374 396 4392 414
rect 4374 414 4392 432
rect 4374 432 4392 450
rect 4374 450 4392 468
rect 4374 468 4392 486
rect 4374 486 4392 504
rect 4374 504 4392 522
rect 4374 522 4392 540
rect 4374 540 4392 558
rect 4374 558 4392 576
rect 4374 576 4392 594
rect 4374 594 4392 612
rect 4374 612 4392 630
rect 4374 630 4392 648
rect 4374 648 4392 666
rect 4374 666 4392 684
rect 4374 684 4392 702
rect 4374 864 4392 882
rect 4374 882 4392 900
rect 4374 900 4392 918
rect 4374 918 4392 936
rect 4374 936 4392 954
rect 4374 954 4392 972
rect 4374 972 4392 990
rect 4374 990 4392 1008
rect 4374 1008 4392 1026
rect 4374 1026 4392 1044
rect 4374 1044 4392 1062
rect 4374 1062 4392 1080
rect 4374 1080 4392 1098
rect 4374 1098 4392 1116
rect 4374 1116 4392 1134
rect 4374 1134 4392 1152
rect 4374 1152 4392 1170
rect 4374 1170 4392 1188
rect 4374 1188 4392 1206
rect 4374 1206 4392 1224
rect 4374 1224 4392 1242
rect 4374 1242 4392 1260
rect 4374 1260 4392 1278
rect 4374 1278 4392 1296
rect 4374 1296 4392 1314
rect 4374 1314 4392 1332
rect 4374 1332 4392 1350
rect 4374 1350 4392 1368
rect 4374 1368 4392 1386
rect 4374 1386 4392 1404
rect 4374 1404 4392 1422
rect 4374 1422 4392 1440
rect 4374 1440 4392 1458
rect 4374 1458 4392 1476
rect 4374 1476 4392 1494
rect 4374 1494 4392 1512
rect 4374 1512 4392 1530
rect 4374 1530 4392 1548
rect 4374 1548 4392 1566
rect 4374 1566 4392 1584
rect 4374 1584 4392 1602
rect 4374 1602 4392 1620
rect 4374 1620 4392 1638
rect 4374 1638 4392 1656
rect 4374 1656 4392 1674
rect 4374 1674 4392 1692
rect 4374 1692 4392 1710
rect 4374 1710 4392 1728
rect 4374 1728 4392 1746
rect 4374 1746 4392 1764
rect 4374 1764 4392 1782
rect 4374 1782 4392 1800
rect 4374 1800 4392 1818
rect 4374 2052 4392 2070
rect 4374 2070 4392 2088
rect 4374 2088 4392 2106
rect 4374 2106 4392 2124
rect 4374 2124 4392 2142
rect 4374 2142 4392 2160
rect 4374 2160 4392 2178
rect 4374 2178 4392 2196
rect 4374 2196 4392 2214
rect 4374 2214 4392 2232
rect 4374 2232 4392 2250
rect 4374 2250 4392 2268
rect 4374 2268 4392 2286
rect 4374 2286 4392 2304
rect 4374 2304 4392 2322
rect 4374 2322 4392 2340
rect 4374 2340 4392 2358
rect 4374 2358 4392 2376
rect 4374 2376 4392 2394
rect 4374 2394 4392 2412
rect 4374 2412 4392 2430
rect 4374 2430 4392 2448
rect 4374 2448 4392 2466
rect 4374 2466 4392 2484
rect 4374 2484 4392 2502
rect 4374 2502 4392 2520
rect 4374 2520 4392 2538
rect 4374 2538 4392 2556
rect 4374 2556 4392 2574
rect 4374 2574 4392 2592
rect 4374 2592 4392 2610
rect 4374 2610 4392 2628
rect 4374 2628 4392 2646
rect 4374 2646 4392 2664
rect 4374 2664 4392 2682
rect 4374 2682 4392 2700
rect 4374 2700 4392 2718
rect 4374 2718 4392 2736
rect 4374 2736 4392 2754
rect 4374 2754 4392 2772
rect 4374 2772 4392 2790
rect 4374 2790 4392 2808
rect 4374 2808 4392 2826
rect 4374 2826 4392 2844
rect 4374 2844 4392 2862
rect 4374 2862 4392 2880
rect 4374 2880 4392 2898
rect 4374 2898 4392 2916
rect 4374 2916 4392 2934
rect 4374 2934 4392 2952
rect 4374 2952 4392 2970
rect 4374 2970 4392 2988
rect 4374 2988 4392 3006
rect 4374 3006 4392 3024
rect 4374 3024 4392 3042
rect 4374 3042 4392 3060
rect 4374 3060 4392 3078
rect 4374 3078 4392 3096
rect 4374 3096 4392 3114
rect 4374 3114 4392 3132
rect 4374 3132 4392 3150
rect 4374 3150 4392 3168
rect 4374 3168 4392 3186
rect 4374 3186 4392 3204
rect 4374 3204 4392 3222
rect 4374 3222 4392 3240
rect 4374 3240 4392 3258
rect 4374 3258 4392 3276
rect 4374 3276 4392 3294
rect 4374 3294 4392 3312
rect 4374 3312 4392 3330
rect 4374 3330 4392 3348
rect 4374 3348 4392 3366
rect 4374 3366 4392 3384
rect 4374 3384 4392 3402
rect 4374 3402 4392 3420
rect 4374 3420 4392 3438
rect 4374 3438 4392 3456
rect 4374 3456 4392 3474
rect 4374 3474 4392 3492
rect 4374 3492 4392 3510
rect 4374 3510 4392 3528
rect 4374 3528 4392 3546
rect 4374 3546 4392 3564
rect 4374 3564 4392 3582
rect 4374 3582 4392 3600
rect 4374 3600 4392 3618
rect 4374 3618 4392 3636
rect 4374 3834 4392 3852
rect 4374 3852 4392 3870
rect 4374 3870 4392 3888
rect 4374 3888 4392 3906
rect 4374 3906 4392 3924
rect 4374 3924 4392 3942
rect 4374 3942 4392 3960
rect 4374 3960 4392 3978
rect 4374 3978 4392 3996
rect 4374 3996 4392 4014
rect 4374 4014 4392 4032
rect 4374 4032 4392 4050
rect 4374 4050 4392 4068
rect 4374 4068 4392 4086
rect 4374 4086 4392 4104
rect 4374 4104 4392 4122
rect 4374 4122 4392 4140
rect 4374 4140 4392 4158
rect 4374 4158 4392 4176
rect 4374 4176 4392 4194
rect 4374 4194 4392 4212
rect 4374 4212 4392 4230
rect 4374 4230 4392 4248
rect 4374 4248 4392 4266
rect 4374 4266 4392 4284
rect 4374 4284 4392 4302
rect 4374 4302 4392 4320
rect 4374 4320 4392 4338
rect 4374 4338 4392 4356
rect 4374 4356 4392 4374
rect 4374 4374 4392 4392
rect 4374 4392 4392 4410
rect 4374 4410 4392 4428
rect 4374 4428 4392 4446
rect 4374 4446 4392 4464
rect 4374 4464 4392 4482
rect 4374 4482 4392 4500
rect 4374 4500 4392 4518
rect 4374 4518 4392 4536
rect 4374 4536 4392 4554
rect 4374 4554 4392 4572
rect 4374 4572 4392 4590
rect 4374 4590 4392 4608
rect 4374 4608 4392 4626
rect 4374 4626 4392 4644
rect 4374 4644 4392 4662
rect 4374 4662 4392 4680
rect 4374 4680 4392 4698
rect 4374 4698 4392 4716
rect 4374 4716 4392 4734
rect 4374 4734 4392 4752
rect 4374 4752 4392 4770
rect 4374 4770 4392 4788
rect 4374 4788 4392 4806
rect 4374 4806 4392 4824
rect 4374 4824 4392 4842
rect 4374 4842 4392 4860
rect 4374 4860 4392 4878
rect 4374 4878 4392 4896
rect 4374 4896 4392 4914
rect 4374 4914 4392 4932
rect 4374 4932 4392 4950
rect 4374 4950 4392 4968
rect 4374 4968 4392 4986
rect 4374 4986 4392 5004
rect 4374 5004 4392 5022
rect 4374 5022 4392 5040
rect 4374 5040 4392 5058
rect 4374 5058 4392 5076
rect 4374 5076 4392 5094
rect 4374 5094 4392 5112
rect 4374 5112 4392 5130
rect 4374 5130 4392 5148
rect 4374 5148 4392 5166
rect 4374 5166 4392 5184
rect 4374 5184 4392 5202
rect 4374 5202 4392 5220
rect 4374 5220 4392 5238
rect 4374 5238 4392 5256
rect 4374 5256 4392 5274
rect 4374 5274 4392 5292
rect 4374 5292 4392 5310
rect 4374 5310 4392 5328
rect 4374 5328 4392 5346
rect 4374 5346 4392 5364
rect 4374 5364 4392 5382
rect 4374 5382 4392 5400
rect 4374 5400 4392 5418
rect 4374 5418 4392 5436
rect 4374 5436 4392 5454
rect 4374 5454 4392 5472
rect 4374 5472 4392 5490
rect 4374 5490 4392 5508
rect 4374 5508 4392 5526
rect 4374 5526 4392 5544
rect 4374 5544 4392 5562
rect 4374 5562 4392 5580
rect 4374 5580 4392 5598
rect 4374 5598 4392 5616
rect 4374 5616 4392 5634
rect 4374 5634 4392 5652
rect 4374 5652 4392 5670
rect 4374 5670 4392 5688
rect 4374 5688 4392 5706
rect 4374 5706 4392 5724
rect 4374 5724 4392 5742
rect 4374 5742 4392 5760
rect 4374 5760 4392 5778
rect 4374 5778 4392 5796
rect 4374 5796 4392 5814
rect 4374 5814 4392 5832
rect 4374 5832 4392 5850
rect 4374 5850 4392 5868
rect 4374 5868 4392 5886
rect 4374 5886 4392 5904
rect 4374 5904 4392 5922
rect 4374 5922 4392 5940
rect 4374 5940 4392 5958
rect 4374 5958 4392 5976
rect 4374 5976 4392 5994
rect 4374 5994 4392 6012
rect 4374 6012 4392 6030
rect 4374 6030 4392 6048
rect 4374 6048 4392 6066
rect 4374 6066 4392 6084
rect 4374 6084 4392 6102
rect 4374 6102 4392 6120
rect 4374 6120 4392 6138
rect 4374 6138 4392 6156
rect 4374 6156 4392 6174
rect 4374 6174 4392 6192
rect 4374 6192 4392 6210
rect 4374 6210 4392 6228
rect 4374 6228 4392 6246
rect 4374 6246 4392 6264
rect 4374 6264 4392 6282
rect 4374 6282 4392 6300
rect 4374 6300 4392 6318
rect 4374 6318 4392 6336
rect 4374 6336 4392 6354
rect 4374 6354 4392 6372
rect 4374 6372 4392 6390
rect 4374 6390 4392 6408
rect 4374 6408 4392 6426
rect 4374 6426 4392 6444
rect 4374 6444 4392 6462
rect 4374 6462 4392 6480
rect 4374 6480 4392 6498
rect 4374 6498 4392 6516
rect 4374 6516 4392 6534
rect 4374 6534 4392 6552
rect 4374 6552 4392 6570
rect 4374 6570 4392 6588
rect 4374 6588 4392 6606
rect 4374 6606 4392 6624
rect 4374 6624 4392 6642
rect 4374 6642 4392 6660
rect 4374 6660 4392 6678
rect 4374 6678 4392 6696
rect 4374 6696 4392 6714
rect 4374 6714 4392 6732
rect 4374 6732 4392 6750
rect 4374 6750 4392 6768
rect 4374 6768 4392 6786
rect 4374 6786 4392 6804
rect 4374 6804 4392 6822
rect 4374 7146 4392 7164
rect 4374 7164 4392 7182
rect 4374 7182 4392 7200
rect 4374 7200 4392 7218
rect 4392 72 4410 90
rect 4392 90 4410 108
rect 4392 108 4410 126
rect 4392 126 4410 144
rect 4392 144 4410 162
rect 4392 162 4410 180
rect 4392 180 4410 198
rect 4392 198 4410 216
rect 4392 216 4410 234
rect 4392 234 4410 252
rect 4392 252 4410 270
rect 4392 270 4410 288
rect 4392 288 4410 306
rect 4392 306 4410 324
rect 4392 324 4410 342
rect 4392 342 4410 360
rect 4392 360 4410 378
rect 4392 378 4410 396
rect 4392 396 4410 414
rect 4392 414 4410 432
rect 4392 432 4410 450
rect 4392 450 4410 468
rect 4392 468 4410 486
rect 4392 486 4410 504
rect 4392 504 4410 522
rect 4392 522 4410 540
rect 4392 540 4410 558
rect 4392 558 4410 576
rect 4392 576 4410 594
rect 4392 594 4410 612
rect 4392 612 4410 630
rect 4392 630 4410 648
rect 4392 648 4410 666
rect 4392 666 4410 684
rect 4392 684 4410 702
rect 4392 702 4410 720
rect 4392 864 4410 882
rect 4392 882 4410 900
rect 4392 900 4410 918
rect 4392 918 4410 936
rect 4392 936 4410 954
rect 4392 954 4410 972
rect 4392 972 4410 990
rect 4392 990 4410 1008
rect 4392 1008 4410 1026
rect 4392 1026 4410 1044
rect 4392 1044 4410 1062
rect 4392 1062 4410 1080
rect 4392 1080 4410 1098
rect 4392 1098 4410 1116
rect 4392 1116 4410 1134
rect 4392 1134 4410 1152
rect 4392 1152 4410 1170
rect 4392 1170 4410 1188
rect 4392 1188 4410 1206
rect 4392 1206 4410 1224
rect 4392 1224 4410 1242
rect 4392 1242 4410 1260
rect 4392 1260 4410 1278
rect 4392 1278 4410 1296
rect 4392 1296 4410 1314
rect 4392 1314 4410 1332
rect 4392 1332 4410 1350
rect 4392 1350 4410 1368
rect 4392 1368 4410 1386
rect 4392 1386 4410 1404
rect 4392 1404 4410 1422
rect 4392 1422 4410 1440
rect 4392 1440 4410 1458
rect 4392 1458 4410 1476
rect 4392 1476 4410 1494
rect 4392 1494 4410 1512
rect 4392 1512 4410 1530
rect 4392 1530 4410 1548
rect 4392 1548 4410 1566
rect 4392 1566 4410 1584
rect 4392 1584 4410 1602
rect 4392 1602 4410 1620
rect 4392 1620 4410 1638
rect 4392 1638 4410 1656
rect 4392 1656 4410 1674
rect 4392 1674 4410 1692
rect 4392 1692 4410 1710
rect 4392 1710 4410 1728
rect 4392 1728 4410 1746
rect 4392 1746 4410 1764
rect 4392 1764 4410 1782
rect 4392 1782 4410 1800
rect 4392 1800 4410 1818
rect 4392 1818 4410 1836
rect 4392 2070 4410 2088
rect 4392 2088 4410 2106
rect 4392 2106 4410 2124
rect 4392 2124 4410 2142
rect 4392 2142 4410 2160
rect 4392 2160 4410 2178
rect 4392 2178 4410 2196
rect 4392 2196 4410 2214
rect 4392 2214 4410 2232
rect 4392 2232 4410 2250
rect 4392 2250 4410 2268
rect 4392 2268 4410 2286
rect 4392 2286 4410 2304
rect 4392 2304 4410 2322
rect 4392 2322 4410 2340
rect 4392 2340 4410 2358
rect 4392 2358 4410 2376
rect 4392 2376 4410 2394
rect 4392 2394 4410 2412
rect 4392 2412 4410 2430
rect 4392 2430 4410 2448
rect 4392 2448 4410 2466
rect 4392 2466 4410 2484
rect 4392 2484 4410 2502
rect 4392 2502 4410 2520
rect 4392 2520 4410 2538
rect 4392 2538 4410 2556
rect 4392 2556 4410 2574
rect 4392 2574 4410 2592
rect 4392 2592 4410 2610
rect 4392 2610 4410 2628
rect 4392 2628 4410 2646
rect 4392 2646 4410 2664
rect 4392 2664 4410 2682
rect 4392 2682 4410 2700
rect 4392 2700 4410 2718
rect 4392 2718 4410 2736
rect 4392 2736 4410 2754
rect 4392 2754 4410 2772
rect 4392 2772 4410 2790
rect 4392 2790 4410 2808
rect 4392 2808 4410 2826
rect 4392 2826 4410 2844
rect 4392 2844 4410 2862
rect 4392 2862 4410 2880
rect 4392 2880 4410 2898
rect 4392 2898 4410 2916
rect 4392 2916 4410 2934
rect 4392 2934 4410 2952
rect 4392 2952 4410 2970
rect 4392 2970 4410 2988
rect 4392 2988 4410 3006
rect 4392 3006 4410 3024
rect 4392 3024 4410 3042
rect 4392 3042 4410 3060
rect 4392 3060 4410 3078
rect 4392 3078 4410 3096
rect 4392 3096 4410 3114
rect 4392 3114 4410 3132
rect 4392 3132 4410 3150
rect 4392 3150 4410 3168
rect 4392 3168 4410 3186
rect 4392 3186 4410 3204
rect 4392 3204 4410 3222
rect 4392 3222 4410 3240
rect 4392 3240 4410 3258
rect 4392 3258 4410 3276
rect 4392 3276 4410 3294
rect 4392 3294 4410 3312
rect 4392 3312 4410 3330
rect 4392 3330 4410 3348
rect 4392 3348 4410 3366
rect 4392 3366 4410 3384
rect 4392 3384 4410 3402
rect 4392 3402 4410 3420
rect 4392 3420 4410 3438
rect 4392 3438 4410 3456
rect 4392 3456 4410 3474
rect 4392 3474 4410 3492
rect 4392 3492 4410 3510
rect 4392 3510 4410 3528
rect 4392 3528 4410 3546
rect 4392 3546 4410 3564
rect 4392 3564 4410 3582
rect 4392 3582 4410 3600
rect 4392 3600 4410 3618
rect 4392 3618 4410 3636
rect 4392 3636 4410 3654
rect 4392 3852 4410 3870
rect 4392 3870 4410 3888
rect 4392 3888 4410 3906
rect 4392 3906 4410 3924
rect 4392 3924 4410 3942
rect 4392 3942 4410 3960
rect 4392 3960 4410 3978
rect 4392 3978 4410 3996
rect 4392 3996 4410 4014
rect 4392 4014 4410 4032
rect 4392 4032 4410 4050
rect 4392 4050 4410 4068
rect 4392 4068 4410 4086
rect 4392 4086 4410 4104
rect 4392 4104 4410 4122
rect 4392 4122 4410 4140
rect 4392 4140 4410 4158
rect 4392 4158 4410 4176
rect 4392 4176 4410 4194
rect 4392 4194 4410 4212
rect 4392 4212 4410 4230
rect 4392 4230 4410 4248
rect 4392 4248 4410 4266
rect 4392 4266 4410 4284
rect 4392 4284 4410 4302
rect 4392 4302 4410 4320
rect 4392 4320 4410 4338
rect 4392 4338 4410 4356
rect 4392 4356 4410 4374
rect 4392 4374 4410 4392
rect 4392 4392 4410 4410
rect 4392 4410 4410 4428
rect 4392 4428 4410 4446
rect 4392 4446 4410 4464
rect 4392 4464 4410 4482
rect 4392 4482 4410 4500
rect 4392 4500 4410 4518
rect 4392 4518 4410 4536
rect 4392 4536 4410 4554
rect 4392 4554 4410 4572
rect 4392 4572 4410 4590
rect 4392 4590 4410 4608
rect 4392 4608 4410 4626
rect 4392 4626 4410 4644
rect 4392 4644 4410 4662
rect 4392 4662 4410 4680
rect 4392 4680 4410 4698
rect 4392 4698 4410 4716
rect 4392 4716 4410 4734
rect 4392 4734 4410 4752
rect 4392 4752 4410 4770
rect 4392 4770 4410 4788
rect 4392 4788 4410 4806
rect 4392 4806 4410 4824
rect 4392 4824 4410 4842
rect 4392 4842 4410 4860
rect 4392 4860 4410 4878
rect 4392 4878 4410 4896
rect 4392 4896 4410 4914
rect 4392 4914 4410 4932
rect 4392 4932 4410 4950
rect 4392 4950 4410 4968
rect 4392 4968 4410 4986
rect 4392 4986 4410 5004
rect 4392 5004 4410 5022
rect 4392 5022 4410 5040
rect 4392 5040 4410 5058
rect 4392 5058 4410 5076
rect 4392 5076 4410 5094
rect 4392 5094 4410 5112
rect 4392 5112 4410 5130
rect 4392 5130 4410 5148
rect 4392 5148 4410 5166
rect 4392 5166 4410 5184
rect 4392 5184 4410 5202
rect 4392 5202 4410 5220
rect 4392 5220 4410 5238
rect 4392 5238 4410 5256
rect 4392 5256 4410 5274
rect 4392 5274 4410 5292
rect 4392 5292 4410 5310
rect 4392 5310 4410 5328
rect 4392 5328 4410 5346
rect 4392 5346 4410 5364
rect 4392 5364 4410 5382
rect 4392 5382 4410 5400
rect 4392 5400 4410 5418
rect 4392 5418 4410 5436
rect 4392 5436 4410 5454
rect 4392 5454 4410 5472
rect 4392 5472 4410 5490
rect 4392 5490 4410 5508
rect 4392 5508 4410 5526
rect 4392 5526 4410 5544
rect 4392 5544 4410 5562
rect 4392 5562 4410 5580
rect 4392 5580 4410 5598
rect 4392 5598 4410 5616
rect 4392 5616 4410 5634
rect 4392 5634 4410 5652
rect 4392 5652 4410 5670
rect 4392 5670 4410 5688
rect 4392 5688 4410 5706
rect 4392 5706 4410 5724
rect 4392 5724 4410 5742
rect 4392 5742 4410 5760
rect 4392 5760 4410 5778
rect 4392 5778 4410 5796
rect 4392 5796 4410 5814
rect 4392 5814 4410 5832
rect 4392 5832 4410 5850
rect 4392 5850 4410 5868
rect 4392 5868 4410 5886
rect 4392 5886 4410 5904
rect 4392 5904 4410 5922
rect 4392 5922 4410 5940
rect 4392 5940 4410 5958
rect 4392 5958 4410 5976
rect 4392 5976 4410 5994
rect 4392 5994 4410 6012
rect 4392 6012 4410 6030
rect 4392 6030 4410 6048
rect 4392 6048 4410 6066
rect 4392 6066 4410 6084
rect 4392 6084 4410 6102
rect 4392 6102 4410 6120
rect 4392 6120 4410 6138
rect 4392 6138 4410 6156
rect 4392 6156 4410 6174
rect 4392 6174 4410 6192
rect 4392 6192 4410 6210
rect 4392 6210 4410 6228
rect 4392 6228 4410 6246
rect 4392 6246 4410 6264
rect 4392 6264 4410 6282
rect 4392 6282 4410 6300
rect 4392 6300 4410 6318
rect 4392 6318 4410 6336
rect 4392 6336 4410 6354
rect 4392 6354 4410 6372
rect 4392 6372 4410 6390
rect 4392 6390 4410 6408
rect 4392 6408 4410 6426
rect 4392 6426 4410 6444
rect 4392 6444 4410 6462
rect 4392 6462 4410 6480
rect 4392 6480 4410 6498
rect 4392 6498 4410 6516
rect 4392 6516 4410 6534
rect 4392 6534 4410 6552
rect 4392 6552 4410 6570
rect 4392 6570 4410 6588
rect 4392 6588 4410 6606
rect 4392 6606 4410 6624
rect 4392 6624 4410 6642
rect 4392 6642 4410 6660
rect 4392 6660 4410 6678
rect 4392 6678 4410 6696
rect 4392 6696 4410 6714
rect 4392 6714 4410 6732
rect 4392 6732 4410 6750
rect 4392 6750 4410 6768
rect 4392 6768 4410 6786
rect 4392 6786 4410 6804
rect 4392 6804 4410 6822
rect 4392 6822 4410 6840
rect 4392 6840 4410 6858
rect 4392 7182 4410 7200
rect 4392 7200 4410 7218
rect 4410 90 4428 108
rect 4410 108 4428 126
rect 4410 126 4428 144
rect 4410 144 4428 162
rect 4410 162 4428 180
rect 4410 180 4428 198
rect 4410 198 4428 216
rect 4410 216 4428 234
rect 4410 234 4428 252
rect 4410 252 4428 270
rect 4410 270 4428 288
rect 4410 288 4428 306
rect 4410 306 4428 324
rect 4410 324 4428 342
rect 4410 342 4428 360
rect 4410 360 4428 378
rect 4410 378 4428 396
rect 4410 396 4428 414
rect 4410 414 4428 432
rect 4410 432 4428 450
rect 4410 450 4428 468
rect 4410 468 4428 486
rect 4410 486 4428 504
rect 4410 504 4428 522
rect 4410 522 4428 540
rect 4410 540 4428 558
rect 4410 558 4428 576
rect 4410 576 4428 594
rect 4410 594 4428 612
rect 4410 612 4428 630
rect 4410 630 4428 648
rect 4410 648 4428 666
rect 4410 666 4428 684
rect 4410 684 4428 702
rect 4410 702 4428 720
rect 4410 864 4428 882
rect 4410 882 4428 900
rect 4410 900 4428 918
rect 4410 918 4428 936
rect 4410 936 4428 954
rect 4410 954 4428 972
rect 4410 972 4428 990
rect 4410 990 4428 1008
rect 4410 1008 4428 1026
rect 4410 1026 4428 1044
rect 4410 1044 4428 1062
rect 4410 1062 4428 1080
rect 4410 1080 4428 1098
rect 4410 1098 4428 1116
rect 4410 1116 4428 1134
rect 4410 1134 4428 1152
rect 4410 1152 4428 1170
rect 4410 1170 4428 1188
rect 4410 1188 4428 1206
rect 4410 1206 4428 1224
rect 4410 1224 4428 1242
rect 4410 1242 4428 1260
rect 4410 1260 4428 1278
rect 4410 1278 4428 1296
rect 4410 1296 4428 1314
rect 4410 1314 4428 1332
rect 4410 1332 4428 1350
rect 4410 1350 4428 1368
rect 4410 1368 4428 1386
rect 4410 1386 4428 1404
rect 4410 1404 4428 1422
rect 4410 1422 4428 1440
rect 4410 1440 4428 1458
rect 4410 1458 4428 1476
rect 4410 1476 4428 1494
rect 4410 1494 4428 1512
rect 4410 1512 4428 1530
rect 4410 1530 4428 1548
rect 4410 1548 4428 1566
rect 4410 1566 4428 1584
rect 4410 1584 4428 1602
rect 4410 1602 4428 1620
rect 4410 1620 4428 1638
rect 4410 1638 4428 1656
rect 4410 1656 4428 1674
rect 4410 1674 4428 1692
rect 4410 1692 4428 1710
rect 4410 1710 4428 1728
rect 4410 1728 4428 1746
rect 4410 1746 4428 1764
rect 4410 1764 4428 1782
rect 4410 1782 4428 1800
rect 4410 1800 4428 1818
rect 4410 1818 4428 1836
rect 4410 2088 4428 2106
rect 4410 2106 4428 2124
rect 4410 2124 4428 2142
rect 4410 2142 4428 2160
rect 4410 2160 4428 2178
rect 4410 2178 4428 2196
rect 4410 2196 4428 2214
rect 4410 2214 4428 2232
rect 4410 2232 4428 2250
rect 4410 2250 4428 2268
rect 4410 2268 4428 2286
rect 4410 2286 4428 2304
rect 4410 2304 4428 2322
rect 4410 2322 4428 2340
rect 4410 2340 4428 2358
rect 4410 2358 4428 2376
rect 4410 2376 4428 2394
rect 4410 2394 4428 2412
rect 4410 2412 4428 2430
rect 4410 2430 4428 2448
rect 4410 2448 4428 2466
rect 4410 2466 4428 2484
rect 4410 2484 4428 2502
rect 4410 2502 4428 2520
rect 4410 2520 4428 2538
rect 4410 2538 4428 2556
rect 4410 2556 4428 2574
rect 4410 2574 4428 2592
rect 4410 2592 4428 2610
rect 4410 2610 4428 2628
rect 4410 2628 4428 2646
rect 4410 2646 4428 2664
rect 4410 2664 4428 2682
rect 4410 2682 4428 2700
rect 4410 2700 4428 2718
rect 4410 2718 4428 2736
rect 4410 2736 4428 2754
rect 4410 2754 4428 2772
rect 4410 2772 4428 2790
rect 4410 2790 4428 2808
rect 4410 2808 4428 2826
rect 4410 2826 4428 2844
rect 4410 2844 4428 2862
rect 4410 2862 4428 2880
rect 4410 2880 4428 2898
rect 4410 2898 4428 2916
rect 4410 2916 4428 2934
rect 4410 2934 4428 2952
rect 4410 2952 4428 2970
rect 4410 2970 4428 2988
rect 4410 2988 4428 3006
rect 4410 3006 4428 3024
rect 4410 3024 4428 3042
rect 4410 3042 4428 3060
rect 4410 3060 4428 3078
rect 4410 3078 4428 3096
rect 4410 3096 4428 3114
rect 4410 3114 4428 3132
rect 4410 3132 4428 3150
rect 4410 3150 4428 3168
rect 4410 3168 4428 3186
rect 4410 3186 4428 3204
rect 4410 3204 4428 3222
rect 4410 3222 4428 3240
rect 4410 3240 4428 3258
rect 4410 3258 4428 3276
rect 4410 3276 4428 3294
rect 4410 3294 4428 3312
rect 4410 3312 4428 3330
rect 4410 3330 4428 3348
rect 4410 3348 4428 3366
rect 4410 3366 4428 3384
rect 4410 3384 4428 3402
rect 4410 3402 4428 3420
rect 4410 3420 4428 3438
rect 4410 3438 4428 3456
rect 4410 3456 4428 3474
rect 4410 3474 4428 3492
rect 4410 3492 4428 3510
rect 4410 3510 4428 3528
rect 4410 3528 4428 3546
rect 4410 3546 4428 3564
rect 4410 3564 4428 3582
rect 4410 3582 4428 3600
rect 4410 3600 4428 3618
rect 4410 3618 4428 3636
rect 4410 3636 4428 3654
rect 4410 3654 4428 3672
rect 4410 3888 4428 3906
rect 4410 3906 4428 3924
rect 4410 3924 4428 3942
rect 4410 3942 4428 3960
rect 4410 3960 4428 3978
rect 4410 3978 4428 3996
rect 4410 3996 4428 4014
rect 4410 4014 4428 4032
rect 4410 4032 4428 4050
rect 4410 4050 4428 4068
rect 4410 4068 4428 4086
rect 4410 4086 4428 4104
rect 4410 4104 4428 4122
rect 4410 4122 4428 4140
rect 4410 4140 4428 4158
rect 4410 4158 4428 4176
rect 4410 4176 4428 4194
rect 4410 4194 4428 4212
rect 4410 4212 4428 4230
rect 4410 4230 4428 4248
rect 4410 4248 4428 4266
rect 4410 4266 4428 4284
rect 4410 4284 4428 4302
rect 4410 4302 4428 4320
rect 4410 4320 4428 4338
rect 4410 4338 4428 4356
rect 4410 4356 4428 4374
rect 4410 4374 4428 4392
rect 4410 4392 4428 4410
rect 4410 4410 4428 4428
rect 4410 4428 4428 4446
rect 4410 4446 4428 4464
rect 4410 4464 4428 4482
rect 4410 4482 4428 4500
rect 4410 4500 4428 4518
rect 4410 4518 4428 4536
rect 4410 4536 4428 4554
rect 4410 4554 4428 4572
rect 4410 4572 4428 4590
rect 4410 4590 4428 4608
rect 4410 4608 4428 4626
rect 4410 4626 4428 4644
rect 4410 4644 4428 4662
rect 4410 4662 4428 4680
rect 4410 4680 4428 4698
rect 4410 4698 4428 4716
rect 4410 4716 4428 4734
rect 4410 4734 4428 4752
rect 4410 4752 4428 4770
rect 4410 4770 4428 4788
rect 4410 4788 4428 4806
rect 4410 4806 4428 4824
rect 4410 4824 4428 4842
rect 4410 4842 4428 4860
rect 4410 4860 4428 4878
rect 4410 4878 4428 4896
rect 4410 4896 4428 4914
rect 4410 4914 4428 4932
rect 4410 4932 4428 4950
rect 4410 4950 4428 4968
rect 4410 4968 4428 4986
rect 4410 4986 4428 5004
rect 4410 5004 4428 5022
rect 4410 5022 4428 5040
rect 4410 5040 4428 5058
rect 4410 5058 4428 5076
rect 4410 5076 4428 5094
rect 4410 5094 4428 5112
rect 4410 5112 4428 5130
rect 4410 5130 4428 5148
rect 4410 5148 4428 5166
rect 4410 5166 4428 5184
rect 4410 5184 4428 5202
rect 4410 5202 4428 5220
rect 4410 5220 4428 5238
rect 4410 5238 4428 5256
rect 4410 5256 4428 5274
rect 4410 5274 4428 5292
rect 4410 5292 4428 5310
rect 4410 5310 4428 5328
rect 4410 5328 4428 5346
rect 4410 5346 4428 5364
rect 4410 5364 4428 5382
rect 4410 5382 4428 5400
rect 4410 5400 4428 5418
rect 4410 5418 4428 5436
rect 4410 5436 4428 5454
rect 4410 5454 4428 5472
rect 4410 5472 4428 5490
rect 4410 5490 4428 5508
rect 4410 5508 4428 5526
rect 4410 5526 4428 5544
rect 4410 5544 4428 5562
rect 4410 5562 4428 5580
rect 4410 5580 4428 5598
rect 4410 5598 4428 5616
rect 4410 5616 4428 5634
rect 4410 5634 4428 5652
rect 4410 5652 4428 5670
rect 4410 5670 4428 5688
rect 4410 5688 4428 5706
rect 4410 5706 4428 5724
rect 4410 5724 4428 5742
rect 4410 5742 4428 5760
rect 4410 5760 4428 5778
rect 4410 5778 4428 5796
rect 4410 5796 4428 5814
rect 4410 5814 4428 5832
rect 4410 5832 4428 5850
rect 4410 5850 4428 5868
rect 4410 5868 4428 5886
rect 4410 5886 4428 5904
rect 4410 5904 4428 5922
rect 4410 5922 4428 5940
rect 4410 5940 4428 5958
rect 4410 5958 4428 5976
rect 4410 5976 4428 5994
rect 4410 5994 4428 6012
rect 4410 6012 4428 6030
rect 4410 6030 4428 6048
rect 4410 6048 4428 6066
rect 4410 6066 4428 6084
rect 4410 6084 4428 6102
rect 4410 6102 4428 6120
rect 4410 6120 4428 6138
rect 4410 6138 4428 6156
rect 4410 6156 4428 6174
rect 4410 6174 4428 6192
rect 4410 6192 4428 6210
rect 4410 6210 4428 6228
rect 4410 6228 4428 6246
rect 4410 6246 4428 6264
rect 4410 6264 4428 6282
rect 4410 6282 4428 6300
rect 4410 6300 4428 6318
rect 4410 6318 4428 6336
rect 4410 6336 4428 6354
rect 4410 6354 4428 6372
rect 4410 6372 4428 6390
rect 4410 6390 4428 6408
rect 4410 6408 4428 6426
rect 4410 6426 4428 6444
rect 4410 6444 4428 6462
rect 4410 6462 4428 6480
rect 4410 6480 4428 6498
rect 4410 6498 4428 6516
rect 4410 6516 4428 6534
rect 4410 6534 4428 6552
rect 4410 6552 4428 6570
rect 4410 6570 4428 6588
rect 4410 6588 4428 6606
rect 4410 6606 4428 6624
rect 4410 6624 4428 6642
rect 4410 6642 4428 6660
rect 4410 6660 4428 6678
rect 4410 6678 4428 6696
rect 4410 6696 4428 6714
rect 4410 6714 4428 6732
rect 4410 6732 4428 6750
rect 4410 6750 4428 6768
rect 4410 6768 4428 6786
rect 4410 6786 4428 6804
rect 4410 6804 4428 6822
rect 4410 6822 4428 6840
rect 4410 6840 4428 6858
rect 4410 6858 4428 6876
rect 4428 90 4446 108
rect 4428 108 4446 126
rect 4428 126 4446 144
rect 4428 144 4446 162
rect 4428 162 4446 180
rect 4428 180 4446 198
rect 4428 198 4446 216
rect 4428 216 4446 234
rect 4428 234 4446 252
rect 4428 252 4446 270
rect 4428 270 4446 288
rect 4428 288 4446 306
rect 4428 306 4446 324
rect 4428 324 4446 342
rect 4428 342 4446 360
rect 4428 360 4446 378
rect 4428 378 4446 396
rect 4428 396 4446 414
rect 4428 414 4446 432
rect 4428 432 4446 450
rect 4428 450 4446 468
rect 4428 468 4446 486
rect 4428 486 4446 504
rect 4428 504 4446 522
rect 4428 522 4446 540
rect 4428 540 4446 558
rect 4428 558 4446 576
rect 4428 576 4446 594
rect 4428 594 4446 612
rect 4428 612 4446 630
rect 4428 630 4446 648
rect 4428 648 4446 666
rect 4428 666 4446 684
rect 4428 684 4446 702
rect 4428 702 4446 720
rect 4428 864 4446 882
rect 4428 882 4446 900
rect 4428 900 4446 918
rect 4428 918 4446 936
rect 4428 936 4446 954
rect 4428 954 4446 972
rect 4428 972 4446 990
rect 4428 990 4446 1008
rect 4428 1008 4446 1026
rect 4428 1026 4446 1044
rect 4428 1044 4446 1062
rect 4428 1062 4446 1080
rect 4428 1080 4446 1098
rect 4428 1098 4446 1116
rect 4428 1116 4446 1134
rect 4428 1134 4446 1152
rect 4428 1152 4446 1170
rect 4428 1170 4446 1188
rect 4428 1188 4446 1206
rect 4428 1206 4446 1224
rect 4428 1224 4446 1242
rect 4428 1242 4446 1260
rect 4428 1260 4446 1278
rect 4428 1278 4446 1296
rect 4428 1296 4446 1314
rect 4428 1314 4446 1332
rect 4428 1332 4446 1350
rect 4428 1350 4446 1368
rect 4428 1368 4446 1386
rect 4428 1386 4446 1404
rect 4428 1404 4446 1422
rect 4428 1422 4446 1440
rect 4428 1440 4446 1458
rect 4428 1458 4446 1476
rect 4428 1476 4446 1494
rect 4428 1494 4446 1512
rect 4428 1512 4446 1530
rect 4428 1530 4446 1548
rect 4428 1548 4446 1566
rect 4428 1566 4446 1584
rect 4428 1584 4446 1602
rect 4428 1602 4446 1620
rect 4428 1620 4446 1638
rect 4428 1638 4446 1656
rect 4428 1656 4446 1674
rect 4428 1674 4446 1692
rect 4428 1692 4446 1710
rect 4428 1710 4446 1728
rect 4428 1728 4446 1746
rect 4428 1746 4446 1764
rect 4428 1764 4446 1782
rect 4428 1782 4446 1800
rect 4428 1800 4446 1818
rect 4428 1818 4446 1836
rect 4428 1836 4446 1854
rect 4428 2088 4446 2106
rect 4428 2106 4446 2124
rect 4428 2124 4446 2142
rect 4428 2142 4446 2160
rect 4428 2160 4446 2178
rect 4428 2178 4446 2196
rect 4428 2196 4446 2214
rect 4428 2214 4446 2232
rect 4428 2232 4446 2250
rect 4428 2250 4446 2268
rect 4428 2268 4446 2286
rect 4428 2286 4446 2304
rect 4428 2304 4446 2322
rect 4428 2322 4446 2340
rect 4428 2340 4446 2358
rect 4428 2358 4446 2376
rect 4428 2376 4446 2394
rect 4428 2394 4446 2412
rect 4428 2412 4446 2430
rect 4428 2430 4446 2448
rect 4428 2448 4446 2466
rect 4428 2466 4446 2484
rect 4428 2484 4446 2502
rect 4428 2502 4446 2520
rect 4428 2520 4446 2538
rect 4428 2538 4446 2556
rect 4428 2556 4446 2574
rect 4428 2574 4446 2592
rect 4428 2592 4446 2610
rect 4428 2610 4446 2628
rect 4428 2628 4446 2646
rect 4428 2646 4446 2664
rect 4428 2664 4446 2682
rect 4428 2682 4446 2700
rect 4428 2700 4446 2718
rect 4428 2718 4446 2736
rect 4428 2736 4446 2754
rect 4428 2754 4446 2772
rect 4428 2772 4446 2790
rect 4428 2790 4446 2808
rect 4428 2808 4446 2826
rect 4428 2826 4446 2844
rect 4428 2844 4446 2862
rect 4428 2862 4446 2880
rect 4428 2880 4446 2898
rect 4428 2898 4446 2916
rect 4428 2916 4446 2934
rect 4428 2934 4446 2952
rect 4428 2952 4446 2970
rect 4428 2970 4446 2988
rect 4428 2988 4446 3006
rect 4428 3006 4446 3024
rect 4428 3024 4446 3042
rect 4428 3042 4446 3060
rect 4428 3060 4446 3078
rect 4428 3078 4446 3096
rect 4428 3096 4446 3114
rect 4428 3114 4446 3132
rect 4428 3132 4446 3150
rect 4428 3150 4446 3168
rect 4428 3168 4446 3186
rect 4428 3186 4446 3204
rect 4428 3204 4446 3222
rect 4428 3222 4446 3240
rect 4428 3240 4446 3258
rect 4428 3258 4446 3276
rect 4428 3276 4446 3294
rect 4428 3294 4446 3312
rect 4428 3312 4446 3330
rect 4428 3330 4446 3348
rect 4428 3348 4446 3366
rect 4428 3366 4446 3384
rect 4428 3384 4446 3402
rect 4428 3402 4446 3420
rect 4428 3420 4446 3438
rect 4428 3438 4446 3456
rect 4428 3456 4446 3474
rect 4428 3474 4446 3492
rect 4428 3492 4446 3510
rect 4428 3510 4446 3528
rect 4428 3528 4446 3546
rect 4428 3546 4446 3564
rect 4428 3564 4446 3582
rect 4428 3582 4446 3600
rect 4428 3600 4446 3618
rect 4428 3618 4446 3636
rect 4428 3636 4446 3654
rect 4428 3654 4446 3672
rect 4428 3672 4446 3690
rect 4428 3690 4446 3708
rect 4428 3906 4446 3924
rect 4428 3924 4446 3942
rect 4428 3942 4446 3960
rect 4428 3960 4446 3978
rect 4428 3978 4446 3996
rect 4428 3996 4446 4014
rect 4428 4014 4446 4032
rect 4428 4032 4446 4050
rect 4428 4050 4446 4068
rect 4428 4068 4446 4086
rect 4428 4086 4446 4104
rect 4428 4104 4446 4122
rect 4428 4122 4446 4140
rect 4428 4140 4446 4158
rect 4428 4158 4446 4176
rect 4428 4176 4446 4194
rect 4428 4194 4446 4212
rect 4428 4212 4446 4230
rect 4428 4230 4446 4248
rect 4428 4248 4446 4266
rect 4428 4266 4446 4284
rect 4428 4284 4446 4302
rect 4428 4302 4446 4320
rect 4428 4320 4446 4338
rect 4428 4338 4446 4356
rect 4428 4356 4446 4374
rect 4428 4374 4446 4392
rect 4428 4392 4446 4410
rect 4428 4410 4446 4428
rect 4428 4428 4446 4446
rect 4428 4446 4446 4464
rect 4428 4464 4446 4482
rect 4428 4482 4446 4500
rect 4428 4500 4446 4518
rect 4428 4518 4446 4536
rect 4428 4536 4446 4554
rect 4428 4554 4446 4572
rect 4428 4572 4446 4590
rect 4428 4590 4446 4608
rect 4428 4608 4446 4626
rect 4428 4626 4446 4644
rect 4428 4644 4446 4662
rect 4428 4662 4446 4680
rect 4428 4680 4446 4698
rect 4428 4698 4446 4716
rect 4428 4716 4446 4734
rect 4428 4734 4446 4752
rect 4428 4752 4446 4770
rect 4428 4770 4446 4788
rect 4428 4788 4446 4806
rect 4428 4806 4446 4824
rect 4428 4824 4446 4842
rect 4428 4842 4446 4860
rect 4428 4860 4446 4878
rect 4428 4878 4446 4896
rect 4428 4896 4446 4914
rect 4428 4914 4446 4932
rect 4428 4932 4446 4950
rect 4428 4950 4446 4968
rect 4428 4968 4446 4986
rect 4428 4986 4446 5004
rect 4428 5004 4446 5022
rect 4428 5022 4446 5040
rect 4428 5040 4446 5058
rect 4428 5058 4446 5076
rect 4428 5076 4446 5094
rect 4428 5094 4446 5112
rect 4428 5112 4446 5130
rect 4428 5130 4446 5148
rect 4428 5148 4446 5166
rect 4428 5166 4446 5184
rect 4428 5184 4446 5202
rect 4428 5202 4446 5220
rect 4428 5220 4446 5238
rect 4428 5238 4446 5256
rect 4428 5256 4446 5274
rect 4428 5274 4446 5292
rect 4428 5292 4446 5310
rect 4428 5310 4446 5328
rect 4428 5328 4446 5346
rect 4428 5346 4446 5364
rect 4428 5364 4446 5382
rect 4428 5382 4446 5400
rect 4428 5400 4446 5418
rect 4428 5418 4446 5436
rect 4428 5436 4446 5454
rect 4428 5454 4446 5472
rect 4428 5472 4446 5490
rect 4428 5490 4446 5508
rect 4428 5508 4446 5526
rect 4428 5526 4446 5544
rect 4428 5544 4446 5562
rect 4428 5562 4446 5580
rect 4428 5580 4446 5598
rect 4428 5598 4446 5616
rect 4428 5616 4446 5634
rect 4428 5634 4446 5652
rect 4428 5652 4446 5670
rect 4428 5670 4446 5688
rect 4428 5688 4446 5706
rect 4428 5706 4446 5724
rect 4428 5724 4446 5742
rect 4428 5742 4446 5760
rect 4428 5760 4446 5778
rect 4428 5778 4446 5796
rect 4428 5796 4446 5814
rect 4428 5814 4446 5832
rect 4428 5832 4446 5850
rect 4428 5850 4446 5868
rect 4428 5868 4446 5886
rect 4428 5886 4446 5904
rect 4428 5904 4446 5922
rect 4428 5922 4446 5940
rect 4428 5940 4446 5958
rect 4428 5958 4446 5976
rect 4428 5976 4446 5994
rect 4428 5994 4446 6012
rect 4428 6012 4446 6030
rect 4428 6030 4446 6048
rect 4428 6048 4446 6066
rect 4428 6066 4446 6084
rect 4428 6084 4446 6102
rect 4428 6102 4446 6120
rect 4428 6120 4446 6138
rect 4428 6138 4446 6156
rect 4428 6156 4446 6174
rect 4428 6174 4446 6192
rect 4428 6192 4446 6210
rect 4428 6210 4446 6228
rect 4428 6228 4446 6246
rect 4428 6246 4446 6264
rect 4428 6264 4446 6282
rect 4428 6282 4446 6300
rect 4428 6300 4446 6318
rect 4428 6318 4446 6336
rect 4428 6336 4446 6354
rect 4428 6354 4446 6372
rect 4428 6372 4446 6390
rect 4428 6390 4446 6408
rect 4428 6408 4446 6426
rect 4428 6426 4446 6444
rect 4428 6444 4446 6462
rect 4428 6462 4446 6480
rect 4428 6480 4446 6498
rect 4428 6498 4446 6516
rect 4428 6516 4446 6534
rect 4428 6534 4446 6552
rect 4428 6552 4446 6570
rect 4428 6570 4446 6588
rect 4428 6588 4446 6606
rect 4428 6606 4446 6624
rect 4428 6624 4446 6642
rect 4428 6642 4446 6660
rect 4428 6660 4446 6678
rect 4428 6678 4446 6696
rect 4428 6696 4446 6714
rect 4428 6714 4446 6732
rect 4428 6732 4446 6750
rect 4428 6750 4446 6768
rect 4428 6768 4446 6786
rect 4428 6786 4446 6804
rect 4428 6804 4446 6822
rect 4428 6822 4446 6840
rect 4428 6840 4446 6858
rect 4428 6858 4446 6876
rect 4428 6876 4446 6894
rect 4428 6894 4446 6912
rect 4446 90 4464 108
rect 4446 108 4464 126
rect 4446 126 4464 144
rect 4446 144 4464 162
rect 4446 162 4464 180
rect 4446 180 4464 198
rect 4446 198 4464 216
rect 4446 216 4464 234
rect 4446 234 4464 252
rect 4446 252 4464 270
rect 4446 270 4464 288
rect 4446 288 4464 306
rect 4446 306 4464 324
rect 4446 324 4464 342
rect 4446 342 4464 360
rect 4446 360 4464 378
rect 4446 378 4464 396
rect 4446 396 4464 414
rect 4446 414 4464 432
rect 4446 432 4464 450
rect 4446 450 4464 468
rect 4446 468 4464 486
rect 4446 486 4464 504
rect 4446 504 4464 522
rect 4446 522 4464 540
rect 4446 540 4464 558
rect 4446 558 4464 576
rect 4446 576 4464 594
rect 4446 594 4464 612
rect 4446 612 4464 630
rect 4446 630 4464 648
rect 4446 648 4464 666
rect 4446 666 4464 684
rect 4446 684 4464 702
rect 4446 702 4464 720
rect 4446 720 4464 738
rect 4446 864 4464 882
rect 4446 882 4464 900
rect 4446 900 4464 918
rect 4446 918 4464 936
rect 4446 936 4464 954
rect 4446 954 4464 972
rect 4446 972 4464 990
rect 4446 990 4464 1008
rect 4446 1008 4464 1026
rect 4446 1026 4464 1044
rect 4446 1044 4464 1062
rect 4446 1062 4464 1080
rect 4446 1080 4464 1098
rect 4446 1098 4464 1116
rect 4446 1116 4464 1134
rect 4446 1134 4464 1152
rect 4446 1152 4464 1170
rect 4446 1170 4464 1188
rect 4446 1188 4464 1206
rect 4446 1206 4464 1224
rect 4446 1224 4464 1242
rect 4446 1242 4464 1260
rect 4446 1260 4464 1278
rect 4446 1278 4464 1296
rect 4446 1296 4464 1314
rect 4446 1314 4464 1332
rect 4446 1332 4464 1350
rect 4446 1350 4464 1368
rect 4446 1368 4464 1386
rect 4446 1386 4464 1404
rect 4446 1404 4464 1422
rect 4446 1422 4464 1440
rect 4446 1440 4464 1458
rect 4446 1458 4464 1476
rect 4446 1476 4464 1494
rect 4446 1494 4464 1512
rect 4446 1512 4464 1530
rect 4446 1530 4464 1548
rect 4446 1548 4464 1566
rect 4446 1566 4464 1584
rect 4446 1584 4464 1602
rect 4446 1602 4464 1620
rect 4446 1620 4464 1638
rect 4446 1638 4464 1656
rect 4446 1656 4464 1674
rect 4446 1674 4464 1692
rect 4446 1692 4464 1710
rect 4446 1710 4464 1728
rect 4446 1728 4464 1746
rect 4446 1746 4464 1764
rect 4446 1764 4464 1782
rect 4446 1782 4464 1800
rect 4446 1800 4464 1818
rect 4446 1818 4464 1836
rect 4446 1836 4464 1854
rect 4446 1854 4464 1872
rect 4446 2106 4464 2124
rect 4446 2124 4464 2142
rect 4446 2142 4464 2160
rect 4446 2160 4464 2178
rect 4446 2178 4464 2196
rect 4446 2196 4464 2214
rect 4446 2214 4464 2232
rect 4446 2232 4464 2250
rect 4446 2250 4464 2268
rect 4446 2268 4464 2286
rect 4446 2286 4464 2304
rect 4446 2304 4464 2322
rect 4446 2322 4464 2340
rect 4446 2340 4464 2358
rect 4446 2358 4464 2376
rect 4446 2376 4464 2394
rect 4446 2394 4464 2412
rect 4446 2412 4464 2430
rect 4446 2430 4464 2448
rect 4446 2448 4464 2466
rect 4446 2466 4464 2484
rect 4446 2484 4464 2502
rect 4446 2502 4464 2520
rect 4446 2520 4464 2538
rect 4446 2538 4464 2556
rect 4446 2556 4464 2574
rect 4446 2574 4464 2592
rect 4446 2592 4464 2610
rect 4446 2610 4464 2628
rect 4446 2628 4464 2646
rect 4446 2646 4464 2664
rect 4446 2664 4464 2682
rect 4446 2682 4464 2700
rect 4446 2700 4464 2718
rect 4446 2718 4464 2736
rect 4446 2736 4464 2754
rect 4446 2754 4464 2772
rect 4446 2772 4464 2790
rect 4446 2790 4464 2808
rect 4446 2808 4464 2826
rect 4446 2826 4464 2844
rect 4446 2844 4464 2862
rect 4446 2862 4464 2880
rect 4446 2880 4464 2898
rect 4446 2898 4464 2916
rect 4446 2916 4464 2934
rect 4446 2934 4464 2952
rect 4446 2952 4464 2970
rect 4446 2970 4464 2988
rect 4446 2988 4464 3006
rect 4446 3006 4464 3024
rect 4446 3024 4464 3042
rect 4446 3042 4464 3060
rect 4446 3060 4464 3078
rect 4446 3078 4464 3096
rect 4446 3096 4464 3114
rect 4446 3114 4464 3132
rect 4446 3132 4464 3150
rect 4446 3150 4464 3168
rect 4446 3168 4464 3186
rect 4446 3186 4464 3204
rect 4446 3204 4464 3222
rect 4446 3222 4464 3240
rect 4446 3240 4464 3258
rect 4446 3258 4464 3276
rect 4446 3276 4464 3294
rect 4446 3294 4464 3312
rect 4446 3312 4464 3330
rect 4446 3330 4464 3348
rect 4446 3348 4464 3366
rect 4446 3366 4464 3384
rect 4446 3384 4464 3402
rect 4446 3402 4464 3420
rect 4446 3420 4464 3438
rect 4446 3438 4464 3456
rect 4446 3456 4464 3474
rect 4446 3474 4464 3492
rect 4446 3492 4464 3510
rect 4446 3510 4464 3528
rect 4446 3528 4464 3546
rect 4446 3546 4464 3564
rect 4446 3564 4464 3582
rect 4446 3582 4464 3600
rect 4446 3600 4464 3618
rect 4446 3618 4464 3636
rect 4446 3636 4464 3654
rect 4446 3654 4464 3672
rect 4446 3672 4464 3690
rect 4446 3690 4464 3708
rect 4446 3708 4464 3726
rect 4446 3924 4464 3942
rect 4446 3942 4464 3960
rect 4446 3960 4464 3978
rect 4446 3978 4464 3996
rect 4446 3996 4464 4014
rect 4446 4014 4464 4032
rect 4446 4032 4464 4050
rect 4446 4050 4464 4068
rect 4446 4068 4464 4086
rect 4446 4086 4464 4104
rect 4446 4104 4464 4122
rect 4446 4122 4464 4140
rect 4446 4140 4464 4158
rect 4446 4158 4464 4176
rect 4446 4176 4464 4194
rect 4446 4194 4464 4212
rect 4446 4212 4464 4230
rect 4446 4230 4464 4248
rect 4446 4248 4464 4266
rect 4446 4266 4464 4284
rect 4446 4284 4464 4302
rect 4446 4302 4464 4320
rect 4446 4320 4464 4338
rect 4446 4338 4464 4356
rect 4446 4356 4464 4374
rect 4446 4374 4464 4392
rect 4446 4392 4464 4410
rect 4446 4410 4464 4428
rect 4446 4428 4464 4446
rect 4446 4446 4464 4464
rect 4446 4464 4464 4482
rect 4446 4482 4464 4500
rect 4446 4500 4464 4518
rect 4446 4518 4464 4536
rect 4446 4536 4464 4554
rect 4446 4554 4464 4572
rect 4446 4572 4464 4590
rect 4446 4590 4464 4608
rect 4446 4608 4464 4626
rect 4446 4626 4464 4644
rect 4446 4644 4464 4662
rect 4446 4662 4464 4680
rect 4446 4680 4464 4698
rect 4446 4698 4464 4716
rect 4446 4716 4464 4734
rect 4446 4734 4464 4752
rect 4446 4752 4464 4770
rect 4446 4770 4464 4788
rect 4446 4788 4464 4806
rect 4446 4806 4464 4824
rect 4446 4824 4464 4842
rect 4446 4842 4464 4860
rect 4446 4860 4464 4878
rect 4446 4878 4464 4896
rect 4446 4896 4464 4914
rect 4446 4914 4464 4932
rect 4446 4932 4464 4950
rect 4446 4950 4464 4968
rect 4446 4968 4464 4986
rect 4446 4986 4464 5004
rect 4446 5004 4464 5022
rect 4446 5022 4464 5040
rect 4446 5040 4464 5058
rect 4446 5058 4464 5076
rect 4446 5076 4464 5094
rect 4446 5094 4464 5112
rect 4446 5112 4464 5130
rect 4446 5130 4464 5148
rect 4446 5148 4464 5166
rect 4446 5166 4464 5184
rect 4446 5184 4464 5202
rect 4446 5202 4464 5220
rect 4446 5220 4464 5238
rect 4446 5238 4464 5256
rect 4446 5256 4464 5274
rect 4446 5274 4464 5292
rect 4446 5292 4464 5310
rect 4446 5310 4464 5328
rect 4446 5328 4464 5346
rect 4446 5346 4464 5364
rect 4446 5364 4464 5382
rect 4446 5382 4464 5400
rect 4446 5400 4464 5418
rect 4446 5418 4464 5436
rect 4446 5436 4464 5454
rect 4446 5454 4464 5472
rect 4446 5472 4464 5490
rect 4446 5490 4464 5508
rect 4446 5508 4464 5526
rect 4446 5526 4464 5544
rect 4446 5544 4464 5562
rect 4446 5562 4464 5580
rect 4446 5580 4464 5598
rect 4446 5598 4464 5616
rect 4446 5616 4464 5634
rect 4446 5634 4464 5652
rect 4446 5652 4464 5670
rect 4446 5670 4464 5688
rect 4446 5688 4464 5706
rect 4446 5706 4464 5724
rect 4446 5724 4464 5742
rect 4446 5742 4464 5760
rect 4446 5760 4464 5778
rect 4446 5778 4464 5796
rect 4446 5796 4464 5814
rect 4446 5814 4464 5832
rect 4446 5832 4464 5850
rect 4446 5850 4464 5868
rect 4446 5868 4464 5886
rect 4446 5886 4464 5904
rect 4446 5904 4464 5922
rect 4446 5922 4464 5940
rect 4446 5940 4464 5958
rect 4446 5958 4464 5976
rect 4446 5976 4464 5994
rect 4446 5994 4464 6012
rect 4446 6012 4464 6030
rect 4446 6030 4464 6048
rect 4446 6048 4464 6066
rect 4446 6066 4464 6084
rect 4446 6084 4464 6102
rect 4446 6102 4464 6120
rect 4446 6120 4464 6138
rect 4446 6138 4464 6156
rect 4446 6156 4464 6174
rect 4446 6174 4464 6192
rect 4446 6192 4464 6210
rect 4446 6210 4464 6228
rect 4446 6228 4464 6246
rect 4446 6246 4464 6264
rect 4446 6264 4464 6282
rect 4446 6282 4464 6300
rect 4446 6300 4464 6318
rect 4446 6318 4464 6336
rect 4446 6336 4464 6354
rect 4446 6354 4464 6372
rect 4446 6372 4464 6390
rect 4446 6390 4464 6408
rect 4446 6408 4464 6426
rect 4446 6426 4464 6444
rect 4446 6444 4464 6462
rect 4446 6462 4464 6480
rect 4446 6480 4464 6498
rect 4446 6498 4464 6516
rect 4446 6516 4464 6534
rect 4446 6534 4464 6552
rect 4446 6552 4464 6570
rect 4446 6570 4464 6588
rect 4446 6588 4464 6606
rect 4446 6606 4464 6624
rect 4446 6624 4464 6642
rect 4446 6642 4464 6660
rect 4446 6660 4464 6678
rect 4446 6678 4464 6696
rect 4446 6696 4464 6714
rect 4446 6714 4464 6732
rect 4446 6732 4464 6750
rect 4446 6750 4464 6768
rect 4446 6768 4464 6786
rect 4446 6786 4464 6804
rect 4446 6804 4464 6822
rect 4446 6822 4464 6840
rect 4446 6840 4464 6858
rect 4446 6858 4464 6876
rect 4446 6876 4464 6894
rect 4446 6894 4464 6912
rect 4446 6912 4464 6930
rect 4446 6930 4464 6948
rect 4464 90 4482 108
rect 4464 108 4482 126
rect 4464 126 4482 144
rect 4464 144 4482 162
rect 4464 162 4482 180
rect 4464 180 4482 198
rect 4464 198 4482 216
rect 4464 216 4482 234
rect 4464 234 4482 252
rect 4464 252 4482 270
rect 4464 270 4482 288
rect 4464 288 4482 306
rect 4464 306 4482 324
rect 4464 324 4482 342
rect 4464 342 4482 360
rect 4464 360 4482 378
rect 4464 378 4482 396
rect 4464 396 4482 414
rect 4464 414 4482 432
rect 4464 432 4482 450
rect 4464 450 4482 468
rect 4464 468 4482 486
rect 4464 486 4482 504
rect 4464 504 4482 522
rect 4464 522 4482 540
rect 4464 540 4482 558
rect 4464 558 4482 576
rect 4464 576 4482 594
rect 4464 594 4482 612
rect 4464 612 4482 630
rect 4464 630 4482 648
rect 4464 648 4482 666
rect 4464 666 4482 684
rect 4464 684 4482 702
rect 4464 702 4482 720
rect 4464 720 4482 738
rect 4464 864 4482 882
rect 4464 882 4482 900
rect 4464 900 4482 918
rect 4464 918 4482 936
rect 4464 936 4482 954
rect 4464 954 4482 972
rect 4464 972 4482 990
rect 4464 990 4482 1008
rect 4464 1008 4482 1026
rect 4464 1026 4482 1044
rect 4464 1044 4482 1062
rect 4464 1062 4482 1080
rect 4464 1080 4482 1098
rect 4464 1098 4482 1116
rect 4464 1116 4482 1134
rect 4464 1134 4482 1152
rect 4464 1152 4482 1170
rect 4464 1170 4482 1188
rect 4464 1188 4482 1206
rect 4464 1206 4482 1224
rect 4464 1224 4482 1242
rect 4464 1242 4482 1260
rect 4464 1260 4482 1278
rect 4464 1278 4482 1296
rect 4464 1296 4482 1314
rect 4464 1314 4482 1332
rect 4464 1332 4482 1350
rect 4464 1350 4482 1368
rect 4464 1368 4482 1386
rect 4464 1386 4482 1404
rect 4464 1404 4482 1422
rect 4464 1422 4482 1440
rect 4464 1440 4482 1458
rect 4464 1458 4482 1476
rect 4464 1476 4482 1494
rect 4464 1494 4482 1512
rect 4464 1512 4482 1530
rect 4464 1530 4482 1548
rect 4464 1548 4482 1566
rect 4464 1566 4482 1584
rect 4464 1584 4482 1602
rect 4464 1602 4482 1620
rect 4464 1620 4482 1638
rect 4464 1638 4482 1656
rect 4464 1656 4482 1674
rect 4464 1674 4482 1692
rect 4464 1692 4482 1710
rect 4464 1710 4482 1728
rect 4464 1728 4482 1746
rect 4464 1746 4482 1764
rect 4464 1764 4482 1782
rect 4464 1782 4482 1800
rect 4464 1800 4482 1818
rect 4464 1818 4482 1836
rect 4464 1836 4482 1854
rect 4464 1854 4482 1872
rect 4464 2124 4482 2142
rect 4464 2142 4482 2160
rect 4464 2160 4482 2178
rect 4464 2178 4482 2196
rect 4464 2196 4482 2214
rect 4464 2214 4482 2232
rect 4464 2232 4482 2250
rect 4464 2250 4482 2268
rect 4464 2268 4482 2286
rect 4464 2286 4482 2304
rect 4464 2304 4482 2322
rect 4464 2322 4482 2340
rect 4464 2340 4482 2358
rect 4464 2358 4482 2376
rect 4464 2376 4482 2394
rect 4464 2394 4482 2412
rect 4464 2412 4482 2430
rect 4464 2430 4482 2448
rect 4464 2448 4482 2466
rect 4464 2466 4482 2484
rect 4464 2484 4482 2502
rect 4464 2502 4482 2520
rect 4464 2520 4482 2538
rect 4464 2538 4482 2556
rect 4464 2556 4482 2574
rect 4464 2574 4482 2592
rect 4464 2592 4482 2610
rect 4464 2610 4482 2628
rect 4464 2628 4482 2646
rect 4464 2646 4482 2664
rect 4464 2664 4482 2682
rect 4464 2682 4482 2700
rect 4464 2700 4482 2718
rect 4464 2718 4482 2736
rect 4464 2736 4482 2754
rect 4464 2754 4482 2772
rect 4464 2772 4482 2790
rect 4464 2790 4482 2808
rect 4464 2808 4482 2826
rect 4464 2826 4482 2844
rect 4464 2844 4482 2862
rect 4464 2862 4482 2880
rect 4464 2880 4482 2898
rect 4464 2898 4482 2916
rect 4464 2916 4482 2934
rect 4464 2934 4482 2952
rect 4464 2952 4482 2970
rect 4464 2970 4482 2988
rect 4464 2988 4482 3006
rect 4464 3006 4482 3024
rect 4464 3024 4482 3042
rect 4464 3042 4482 3060
rect 4464 3060 4482 3078
rect 4464 3078 4482 3096
rect 4464 3096 4482 3114
rect 4464 3114 4482 3132
rect 4464 3132 4482 3150
rect 4464 3150 4482 3168
rect 4464 3168 4482 3186
rect 4464 3186 4482 3204
rect 4464 3204 4482 3222
rect 4464 3222 4482 3240
rect 4464 3240 4482 3258
rect 4464 3258 4482 3276
rect 4464 3276 4482 3294
rect 4464 3294 4482 3312
rect 4464 3312 4482 3330
rect 4464 3330 4482 3348
rect 4464 3348 4482 3366
rect 4464 3366 4482 3384
rect 4464 3384 4482 3402
rect 4464 3402 4482 3420
rect 4464 3420 4482 3438
rect 4464 3438 4482 3456
rect 4464 3456 4482 3474
rect 4464 3474 4482 3492
rect 4464 3492 4482 3510
rect 4464 3510 4482 3528
rect 4464 3528 4482 3546
rect 4464 3546 4482 3564
rect 4464 3564 4482 3582
rect 4464 3582 4482 3600
rect 4464 3600 4482 3618
rect 4464 3618 4482 3636
rect 4464 3636 4482 3654
rect 4464 3654 4482 3672
rect 4464 3672 4482 3690
rect 4464 3690 4482 3708
rect 4464 3708 4482 3726
rect 4464 3726 4482 3744
rect 4464 3942 4482 3960
rect 4464 3960 4482 3978
rect 4464 3978 4482 3996
rect 4464 3996 4482 4014
rect 4464 4014 4482 4032
rect 4464 4032 4482 4050
rect 4464 4050 4482 4068
rect 4464 4068 4482 4086
rect 4464 4086 4482 4104
rect 4464 4104 4482 4122
rect 4464 4122 4482 4140
rect 4464 4140 4482 4158
rect 4464 4158 4482 4176
rect 4464 4176 4482 4194
rect 4464 4194 4482 4212
rect 4464 4212 4482 4230
rect 4464 4230 4482 4248
rect 4464 4248 4482 4266
rect 4464 4266 4482 4284
rect 4464 4284 4482 4302
rect 4464 4302 4482 4320
rect 4464 4320 4482 4338
rect 4464 4338 4482 4356
rect 4464 4356 4482 4374
rect 4464 4374 4482 4392
rect 4464 4392 4482 4410
rect 4464 4410 4482 4428
rect 4464 4428 4482 4446
rect 4464 4446 4482 4464
rect 4464 4464 4482 4482
rect 4464 4482 4482 4500
rect 4464 4500 4482 4518
rect 4464 4518 4482 4536
rect 4464 4536 4482 4554
rect 4464 4554 4482 4572
rect 4464 4572 4482 4590
rect 4464 4590 4482 4608
rect 4464 4608 4482 4626
rect 4464 4626 4482 4644
rect 4464 4644 4482 4662
rect 4464 4662 4482 4680
rect 4464 4680 4482 4698
rect 4464 4698 4482 4716
rect 4464 4716 4482 4734
rect 4464 4734 4482 4752
rect 4464 4752 4482 4770
rect 4464 4770 4482 4788
rect 4464 4788 4482 4806
rect 4464 4806 4482 4824
rect 4464 4824 4482 4842
rect 4464 4842 4482 4860
rect 4464 4860 4482 4878
rect 4464 4878 4482 4896
rect 4464 4896 4482 4914
rect 4464 4914 4482 4932
rect 4464 4932 4482 4950
rect 4464 4950 4482 4968
rect 4464 4968 4482 4986
rect 4464 4986 4482 5004
rect 4464 5004 4482 5022
rect 4464 5022 4482 5040
rect 4464 5040 4482 5058
rect 4464 5058 4482 5076
rect 4464 5076 4482 5094
rect 4464 5094 4482 5112
rect 4464 5112 4482 5130
rect 4464 5130 4482 5148
rect 4464 5148 4482 5166
rect 4464 5166 4482 5184
rect 4464 5184 4482 5202
rect 4464 5202 4482 5220
rect 4464 5220 4482 5238
rect 4464 5238 4482 5256
rect 4464 5256 4482 5274
rect 4464 5274 4482 5292
rect 4464 5292 4482 5310
rect 4464 5310 4482 5328
rect 4464 5328 4482 5346
rect 4464 5346 4482 5364
rect 4464 5364 4482 5382
rect 4464 5382 4482 5400
rect 4464 5400 4482 5418
rect 4464 5418 4482 5436
rect 4464 5436 4482 5454
rect 4464 5454 4482 5472
rect 4464 5472 4482 5490
rect 4464 5490 4482 5508
rect 4464 5508 4482 5526
rect 4464 5526 4482 5544
rect 4464 5544 4482 5562
rect 4464 5562 4482 5580
rect 4464 5580 4482 5598
rect 4464 5598 4482 5616
rect 4464 5616 4482 5634
rect 4464 5634 4482 5652
rect 4464 5652 4482 5670
rect 4464 5670 4482 5688
rect 4464 5688 4482 5706
rect 4464 5706 4482 5724
rect 4464 5724 4482 5742
rect 4464 5742 4482 5760
rect 4464 5760 4482 5778
rect 4464 5778 4482 5796
rect 4464 5796 4482 5814
rect 4464 5814 4482 5832
rect 4464 5832 4482 5850
rect 4464 5850 4482 5868
rect 4464 5868 4482 5886
rect 4464 5886 4482 5904
rect 4464 5904 4482 5922
rect 4464 5922 4482 5940
rect 4464 5940 4482 5958
rect 4464 5958 4482 5976
rect 4464 5976 4482 5994
rect 4464 5994 4482 6012
rect 4464 6012 4482 6030
rect 4464 6030 4482 6048
rect 4464 6048 4482 6066
rect 4464 6066 4482 6084
rect 4464 6084 4482 6102
rect 4464 6102 4482 6120
rect 4464 6120 4482 6138
rect 4464 6138 4482 6156
rect 4464 6156 4482 6174
rect 4464 6174 4482 6192
rect 4464 6192 4482 6210
rect 4464 6210 4482 6228
rect 4464 6228 4482 6246
rect 4464 6246 4482 6264
rect 4464 6264 4482 6282
rect 4464 6282 4482 6300
rect 4464 6300 4482 6318
rect 4464 6318 4482 6336
rect 4464 6336 4482 6354
rect 4464 6354 4482 6372
rect 4464 6372 4482 6390
rect 4464 6390 4482 6408
rect 4464 6408 4482 6426
rect 4464 6426 4482 6444
rect 4464 6444 4482 6462
rect 4464 6462 4482 6480
rect 4464 6480 4482 6498
rect 4464 6498 4482 6516
rect 4464 6516 4482 6534
rect 4464 6534 4482 6552
rect 4464 6552 4482 6570
rect 4464 6570 4482 6588
rect 4464 6588 4482 6606
rect 4464 6606 4482 6624
rect 4464 6624 4482 6642
rect 4464 6642 4482 6660
rect 4464 6660 4482 6678
rect 4464 6678 4482 6696
rect 4464 6696 4482 6714
rect 4464 6714 4482 6732
rect 4464 6732 4482 6750
rect 4464 6750 4482 6768
rect 4464 6768 4482 6786
rect 4464 6786 4482 6804
rect 4464 6804 4482 6822
rect 4464 6822 4482 6840
rect 4464 6840 4482 6858
rect 4464 6858 4482 6876
rect 4464 6876 4482 6894
rect 4464 6894 4482 6912
rect 4464 6912 4482 6930
rect 4464 6930 4482 6948
rect 4464 6948 4482 6966
rect 4464 6966 4482 6984
rect 4482 90 4500 108
rect 4482 108 4500 126
rect 4482 126 4500 144
rect 4482 144 4500 162
rect 4482 162 4500 180
rect 4482 180 4500 198
rect 4482 198 4500 216
rect 4482 216 4500 234
rect 4482 234 4500 252
rect 4482 252 4500 270
rect 4482 270 4500 288
rect 4482 288 4500 306
rect 4482 306 4500 324
rect 4482 324 4500 342
rect 4482 342 4500 360
rect 4482 360 4500 378
rect 4482 378 4500 396
rect 4482 396 4500 414
rect 4482 414 4500 432
rect 4482 432 4500 450
rect 4482 450 4500 468
rect 4482 468 4500 486
rect 4482 486 4500 504
rect 4482 504 4500 522
rect 4482 522 4500 540
rect 4482 540 4500 558
rect 4482 558 4500 576
rect 4482 576 4500 594
rect 4482 594 4500 612
rect 4482 612 4500 630
rect 4482 630 4500 648
rect 4482 648 4500 666
rect 4482 666 4500 684
rect 4482 684 4500 702
rect 4482 702 4500 720
rect 4482 720 4500 738
rect 4482 864 4500 882
rect 4482 882 4500 900
rect 4482 900 4500 918
rect 4482 918 4500 936
rect 4482 936 4500 954
rect 4482 954 4500 972
rect 4482 972 4500 990
rect 4482 990 4500 1008
rect 4482 1008 4500 1026
rect 4482 1026 4500 1044
rect 4482 1044 4500 1062
rect 4482 1062 4500 1080
rect 4482 1080 4500 1098
rect 4482 1098 4500 1116
rect 4482 1116 4500 1134
rect 4482 1134 4500 1152
rect 4482 1152 4500 1170
rect 4482 1170 4500 1188
rect 4482 1188 4500 1206
rect 4482 1206 4500 1224
rect 4482 1224 4500 1242
rect 4482 1242 4500 1260
rect 4482 1260 4500 1278
rect 4482 1278 4500 1296
rect 4482 1296 4500 1314
rect 4482 1314 4500 1332
rect 4482 1332 4500 1350
rect 4482 1350 4500 1368
rect 4482 1368 4500 1386
rect 4482 1386 4500 1404
rect 4482 1404 4500 1422
rect 4482 1422 4500 1440
rect 4482 1440 4500 1458
rect 4482 1458 4500 1476
rect 4482 1476 4500 1494
rect 4482 1494 4500 1512
rect 4482 1512 4500 1530
rect 4482 1530 4500 1548
rect 4482 1548 4500 1566
rect 4482 1566 4500 1584
rect 4482 1584 4500 1602
rect 4482 1602 4500 1620
rect 4482 1620 4500 1638
rect 4482 1638 4500 1656
rect 4482 1656 4500 1674
rect 4482 1674 4500 1692
rect 4482 1692 4500 1710
rect 4482 1710 4500 1728
rect 4482 1728 4500 1746
rect 4482 1746 4500 1764
rect 4482 1764 4500 1782
rect 4482 1782 4500 1800
rect 4482 1800 4500 1818
rect 4482 1818 4500 1836
rect 4482 1836 4500 1854
rect 4482 1854 4500 1872
rect 4482 1872 4500 1890
rect 4482 2124 4500 2142
rect 4482 2142 4500 2160
rect 4482 2160 4500 2178
rect 4482 2178 4500 2196
rect 4482 2196 4500 2214
rect 4482 2214 4500 2232
rect 4482 2232 4500 2250
rect 4482 2250 4500 2268
rect 4482 2268 4500 2286
rect 4482 2286 4500 2304
rect 4482 2304 4500 2322
rect 4482 2322 4500 2340
rect 4482 2340 4500 2358
rect 4482 2358 4500 2376
rect 4482 2376 4500 2394
rect 4482 2394 4500 2412
rect 4482 2412 4500 2430
rect 4482 2430 4500 2448
rect 4482 2448 4500 2466
rect 4482 2466 4500 2484
rect 4482 2484 4500 2502
rect 4482 2502 4500 2520
rect 4482 2520 4500 2538
rect 4482 2538 4500 2556
rect 4482 2556 4500 2574
rect 4482 2574 4500 2592
rect 4482 2592 4500 2610
rect 4482 2610 4500 2628
rect 4482 2628 4500 2646
rect 4482 2646 4500 2664
rect 4482 2664 4500 2682
rect 4482 2682 4500 2700
rect 4482 2700 4500 2718
rect 4482 2718 4500 2736
rect 4482 2736 4500 2754
rect 4482 2754 4500 2772
rect 4482 2772 4500 2790
rect 4482 2790 4500 2808
rect 4482 2808 4500 2826
rect 4482 2826 4500 2844
rect 4482 2844 4500 2862
rect 4482 2862 4500 2880
rect 4482 2880 4500 2898
rect 4482 2898 4500 2916
rect 4482 2916 4500 2934
rect 4482 2934 4500 2952
rect 4482 2952 4500 2970
rect 4482 2970 4500 2988
rect 4482 2988 4500 3006
rect 4482 3006 4500 3024
rect 4482 3024 4500 3042
rect 4482 3042 4500 3060
rect 4482 3060 4500 3078
rect 4482 3078 4500 3096
rect 4482 3096 4500 3114
rect 4482 3114 4500 3132
rect 4482 3132 4500 3150
rect 4482 3150 4500 3168
rect 4482 3168 4500 3186
rect 4482 3186 4500 3204
rect 4482 3204 4500 3222
rect 4482 3222 4500 3240
rect 4482 3240 4500 3258
rect 4482 3258 4500 3276
rect 4482 3276 4500 3294
rect 4482 3294 4500 3312
rect 4482 3312 4500 3330
rect 4482 3330 4500 3348
rect 4482 3348 4500 3366
rect 4482 3366 4500 3384
rect 4482 3384 4500 3402
rect 4482 3402 4500 3420
rect 4482 3420 4500 3438
rect 4482 3438 4500 3456
rect 4482 3456 4500 3474
rect 4482 3474 4500 3492
rect 4482 3492 4500 3510
rect 4482 3510 4500 3528
rect 4482 3528 4500 3546
rect 4482 3546 4500 3564
rect 4482 3564 4500 3582
rect 4482 3582 4500 3600
rect 4482 3600 4500 3618
rect 4482 3618 4500 3636
rect 4482 3636 4500 3654
rect 4482 3654 4500 3672
rect 4482 3672 4500 3690
rect 4482 3690 4500 3708
rect 4482 3708 4500 3726
rect 4482 3726 4500 3744
rect 4482 3744 4500 3762
rect 4482 3978 4500 3996
rect 4482 3996 4500 4014
rect 4482 4014 4500 4032
rect 4482 4032 4500 4050
rect 4482 4050 4500 4068
rect 4482 4068 4500 4086
rect 4482 4086 4500 4104
rect 4482 4104 4500 4122
rect 4482 4122 4500 4140
rect 4482 4140 4500 4158
rect 4482 4158 4500 4176
rect 4482 4176 4500 4194
rect 4482 4194 4500 4212
rect 4482 4212 4500 4230
rect 4482 4230 4500 4248
rect 4482 4248 4500 4266
rect 4482 4266 4500 4284
rect 4482 4284 4500 4302
rect 4482 4302 4500 4320
rect 4482 4320 4500 4338
rect 4482 4338 4500 4356
rect 4482 4356 4500 4374
rect 4482 4374 4500 4392
rect 4482 4392 4500 4410
rect 4482 4410 4500 4428
rect 4482 4428 4500 4446
rect 4482 4446 4500 4464
rect 4482 4464 4500 4482
rect 4482 4482 4500 4500
rect 4482 4500 4500 4518
rect 4482 4518 4500 4536
rect 4482 4536 4500 4554
rect 4482 4554 4500 4572
rect 4482 4572 4500 4590
rect 4482 4590 4500 4608
rect 4482 4608 4500 4626
rect 4482 4626 4500 4644
rect 4482 4644 4500 4662
rect 4482 4662 4500 4680
rect 4482 4680 4500 4698
rect 4482 4698 4500 4716
rect 4482 4716 4500 4734
rect 4482 4734 4500 4752
rect 4482 4752 4500 4770
rect 4482 4770 4500 4788
rect 4482 4788 4500 4806
rect 4482 4806 4500 4824
rect 4482 4824 4500 4842
rect 4482 4842 4500 4860
rect 4482 4860 4500 4878
rect 4482 4878 4500 4896
rect 4482 4896 4500 4914
rect 4482 4914 4500 4932
rect 4482 4932 4500 4950
rect 4482 4950 4500 4968
rect 4482 4968 4500 4986
rect 4482 4986 4500 5004
rect 4482 5004 4500 5022
rect 4482 5022 4500 5040
rect 4482 5040 4500 5058
rect 4482 5058 4500 5076
rect 4482 5076 4500 5094
rect 4482 5094 4500 5112
rect 4482 5112 4500 5130
rect 4482 5130 4500 5148
rect 4482 5148 4500 5166
rect 4482 5166 4500 5184
rect 4482 5184 4500 5202
rect 4482 5202 4500 5220
rect 4482 5220 4500 5238
rect 4482 5238 4500 5256
rect 4482 5256 4500 5274
rect 4482 5274 4500 5292
rect 4482 5292 4500 5310
rect 4482 5310 4500 5328
rect 4482 5328 4500 5346
rect 4482 5346 4500 5364
rect 4482 5364 4500 5382
rect 4482 5382 4500 5400
rect 4482 5400 4500 5418
rect 4482 5418 4500 5436
rect 4482 5436 4500 5454
rect 4482 5454 4500 5472
rect 4482 5472 4500 5490
rect 4482 5490 4500 5508
rect 4482 5508 4500 5526
rect 4482 5526 4500 5544
rect 4482 5544 4500 5562
rect 4482 5562 4500 5580
rect 4482 5580 4500 5598
rect 4482 5598 4500 5616
rect 4482 5616 4500 5634
rect 4482 5634 4500 5652
rect 4482 5652 4500 5670
rect 4482 5670 4500 5688
rect 4482 5688 4500 5706
rect 4482 5706 4500 5724
rect 4482 5724 4500 5742
rect 4482 5742 4500 5760
rect 4482 5760 4500 5778
rect 4482 5778 4500 5796
rect 4482 5796 4500 5814
rect 4482 5814 4500 5832
rect 4482 5832 4500 5850
rect 4482 5850 4500 5868
rect 4482 5868 4500 5886
rect 4482 5886 4500 5904
rect 4482 5904 4500 5922
rect 4482 5922 4500 5940
rect 4482 5940 4500 5958
rect 4482 5958 4500 5976
rect 4482 5976 4500 5994
rect 4482 5994 4500 6012
rect 4482 6012 4500 6030
rect 4482 6030 4500 6048
rect 4482 6048 4500 6066
rect 4482 6066 4500 6084
rect 4482 6084 4500 6102
rect 4482 6102 4500 6120
rect 4482 6120 4500 6138
rect 4482 6138 4500 6156
rect 4482 6156 4500 6174
rect 4482 6174 4500 6192
rect 4482 6192 4500 6210
rect 4482 6210 4500 6228
rect 4482 6228 4500 6246
rect 4482 6246 4500 6264
rect 4482 6264 4500 6282
rect 4482 6282 4500 6300
rect 4482 6300 4500 6318
rect 4482 6318 4500 6336
rect 4482 6336 4500 6354
rect 4482 6354 4500 6372
rect 4482 6372 4500 6390
rect 4482 6390 4500 6408
rect 4482 6408 4500 6426
rect 4482 6426 4500 6444
rect 4482 6444 4500 6462
rect 4482 6462 4500 6480
rect 4482 6480 4500 6498
rect 4482 6498 4500 6516
rect 4482 6516 4500 6534
rect 4482 6534 4500 6552
rect 4482 6552 4500 6570
rect 4482 6570 4500 6588
rect 4482 6588 4500 6606
rect 4482 6606 4500 6624
rect 4482 6624 4500 6642
rect 4482 6642 4500 6660
rect 4482 6660 4500 6678
rect 4482 6678 4500 6696
rect 4482 6696 4500 6714
rect 4482 6714 4500 6732
rect 4482 6732 4500 6750
rect 4482 6750 4500 6768
rect 4482 6768 4500 6786
rect 4482 6786 4500 6804
rect 4482 6804 4500 6822
rect 4482 6822 4500 6840
rect 4482 6840 4500 6858
rect 4482 6858 4500 6876
rect 4482 6876 4500 6894
rect 4482 6894 4500 6912
rect 4482 6912 4500 6930
rect 4482 6930 4500 6948
rect 4482 6948 4500 6966
rect 4482 6966 4500 6984
rect 4482 6984 4500 7002
rect 4482 7002 4500 7020
rect 4500 108 4518 126
rect 4500 126 4518 144
rect 4500 144 4518 162
rect 4500 162 4518 180
rect 4500 180 4518 198
rect 4500 198 4518 216
rect 4500 216 4518 234
rect 4500 234 4518 252
rect 4500 252 4518 270
rect 4500 270 4518 288
rect 4500 288 4518 306
rect 4500 306 4518 324
rect 4500 324 4518 342
rect 4500 342 4518 360
rect 4500 360 4518 378
rect 4500 378 4518 396
rect 4500 396 4518 414
rect 4500 414 4518 432
rect 4500 432 4518 450
rect 4500 450 4518 468
rect 4500 468 4518 486
rect 4500 486 4518 504
rect 4500 504 4518 522
rect 4500 522 4518 540
rect 4500 540 4518 558
rect 4500 558 4518 576
rect 4500 576 4518 594
rect 4500 594 4518 612
rect 4500 612 4518 630
rect 4500 630 4518 648
rect 4500 648 4518 666
rect 4500 666 4518 684
rect 4500 684 4518 702
rect 4500 702 4518 720
rect 4500 720 4518 738
rect 4500 864 4518 882
rect 4500 882 4518 900
rect 4500 900 4518 918
rect 4500 918 4518 936
rect 4500 936 4518 954
rect 4500 954 4518 972
rect 4500 972 4518 990
rect 4500 990 4518 1008
rect 4500 1008 4518 1026
rect 4500 1026 4518 1044
rect 4500 1044 4518 1062
rect 4500 1062 4518 1080
rect 4500 1080 4518 1098
rect 4500 1098 4518 1116
rect 4500 1116 4518 1134
rect 4500 1134 4518 1152
rect 4500 1152 4518 1170
rect 4500 1170 4518 1188
rect 4500 1188 4518 1206
rect 4500 1206 4518 1224
rect 4500 1224 4518 1242
rect 4500 1242 4518 1260
rect 4500 1260 4518 1278
rect 4500 1278 4518 1296
rect 4500 1296 4518 1314
rect 4500 1314 4518 1332
rect 4500 1332 4518 1350
rect 4500 1350 4518 1368
rect 4500 1368 4518 1386
rect 4500 1386 4518 1404
rect 4500 1404 4518 1422
rect 4500 1422 4518 1440
rect 4500 1440 4518 1458
rect 4500 1458 4518 1476
rect 4500 1476 4518 1494
rect 4500 1494 4518 1512
rect 4500 1512 4518 1530
rect 4500 1530 4518 1548
rect 4500 1548 4518 1566
rect 4500 1566 4518 1584
rect 4500 1584 4518 1602
rect 4500 1602 4518 1620
rect 4500 1620 4518 1638
rect 4500 1638 4518 1656
rect 4500 1656 4518 1674
rect 4500 1674 4518 1692
rect 4500 1692 4518 1710
rect 4500 1710 4518 1728
rect 4500 1728 4518 1746
rect 4500 1746 4518 1764
rect 4500 1764 4518 1782
rect 4500 1782 4518 1800
rect 4500 1800 4518 1818
rect 4500 1818 4518 1836
rect 4500 1836 4518 1854
rect 4500 1854 4518 1872
rect 4500 1872 4518 1890
rect 4500 1890 4518 1908
rect 4500 2142 4518 2160
rect 4500 2160 4518 2178
rect 4500 2178 4518 2196
rect 4500 2196 4518 2214
rect 4500 2214 4518 2232
rect 4500 2232 4518 2250
rect 4500 2250 4518 2268
rect 4500 2268 4518 2286
rect 4500 2286 4518 2304
rect 4500 2304 4518 2322
rect 4500 2322 4518 2340
rect 4500 2340 4518 2358
rect 4500 2358 4518 2376
rect 4500 2376 4518 2394
rect 4500 2394 4518 2412
rect 4500 2412 4518 2430
rect 4500 2430 4518 2448
rect 4500 2448 4518 2466
rect 4500 2466 4518 2484
rect 4500 2484 4518 2502
rect 4500 2502 4518 2520
rect 4500 2520 4518 2538
rect 4500 2538 4518 2556
rect 4500 2556 4518 2574
rect 4500 2574 4518 2592
rect 4500 2592 4518 2610
rect 4500 2610 4518 2628
rect 4500 2628 4518 2646
rect 4500 2646 4518 2664
rect 4500 2664 4518 2682
rect 4500 2682 4518 2700
rect 4500 2700 4518 2718
rect 4500 2718 4518 2736
rect 4500 2736 4518 2754
rect 4500 2754 4518 2772
rect 4500 2772 4518 2790
rect 4500 2790 4518 2808
rect 4500 2808 4518 2826
rect 4500 2826 4518 2844
rect 4500 2844 4518 2862
rect 4500 2862 4518 2880
rect 4500 2880 4518 2898
rect 4500 2898 4518 2916
rect 4500 2916 4518 2934
rect 4500 2934 4518 2952
rect 4500 2952 4518 2970
rect 4500 2970 4518 2988
rect 4500 2988 4518 3006
rect 4500 3006 4518 3024
rect 4500 3024 4518 3042
rect 4500 3042 4518 3060
rect 4500 3060 4518 3078
rect 4500 3078 4518 3096
rect 4500 3096 4518 3114
rect 4500 3114 4518 3132
rect 4500 3132 4518 3150
rect 4500 3150 4518 3168
rect 4500 3168 4518 3186
rect 4500 3186 4518 3204
rect 4500 3204 4518 3222
rect 4500 3222 4518 3240
rect 4500 3240 4518 3258
rect 4500 3258 4518 3276
rect 4500 3276 4518 3294
rect 4500 3294 4518 3312
rect 4500 3312 4518 3330
rect 4500 3330 4518 3348
rect 4500 3348 4518 3366
rect 4500 3366 4518 3384
rect 4500 3384 4518 3402
rect 4500 3402 4518 3420
rect 4500 3420 4518 3438
rect 4500 3438 4518 3456
rect 4500 3456 4518 3474
rect 4500 3474 4518 3492
rect 4500 3492 4518 3510
rect 4500 3510 4518 3528
rect 4500 3528 4518 3546
rect 4500 3546 4518 3564
rect 4500 3564 4518 3582
rect 4500 3582 4518 3600
rect 4500 3600 4518 3618
rect 4500 3618 4518 3636
rect 4500 3636 4518 3654
rect 4500 3654 4518 3672
rect 4500 3672 4518 3690
rect 4500 3690 4518 3708
rect 4500 3708 4518 3726
rect 4500 3726 4518 3744
rect 4500 3744 4518 3762
rect 4500 3762 4518 3780
rect 4500 3780 4518 3798
rect 4500 3996 4518 4014
rect 4500 4014 4518 4032
rect 4500 4032 4518 4050
rect 4500 4050 4518 4068
rect 4500 4068 4518 4086
rect 4500 4086 4518 4104
rect 4500 4104 4518 4122
rect 4500 4122 4518 4140
rect 4500 4140 4518 4158
rect 4500 4158 4518 4176
rect 4500 4176 4518 4194
rect 4500 4194 4518 4212
rect 4500 4212 4518 4230
rect 4500 4230 4518 4248
rect 4500 4248 4518 4266
rect 4500 4266 4518 4284
rect 4500 4284 4518 4302
rect 4500 4302 4518 4320
rect 4500 4320 4518 4338
rect 4500 4338 4518 4356
rect 4500 4356 4518 4374
rect 4500 4374 4518 4392
rect 4500 4392 4518 4410
rect 4500 4410 4518 4428
rect 4500 4428 4518 4446
rect 4500 4446 4518 4464
rect 4500 4464 4518 4482
rect 4500 4482 4518 4500
rect 4500 4500 4518 4518
rect 4500 4518 4518 4536
rect 4500 4536 4518 4554
rect 4500 4554 4518 4572
rect 4500 4572 4518 4590
rect 4500 4590 4518 4608
rect 4500 4608 4518 4626
rect 4500 4626 4518 4644
rect 4500 4644 4518 4662
rect 4500 4662 4518 4680
rect 4500 4680 4518 4698
rect 4500 4698 4518 4716
rect 4500 4716 4518 4734
rect 4500 4734 4518 4752
rect 4500 4752 4518 4770
rect 4500 4770 4518 4788
rect 4500 4788 4518 4806
rect 4500 4806 4518 4824
rect 4500 4824 4518 4842
rect 4500 4842 4518 4860
rect 4500 4860 4518 4878
rect 4500 4878 4518 4896
rect 4500 4896 4518 4914
rect 4500 4914 4518 4932
rect 4500 4932 4518 4950
rect 4500 4950 4518 4968
rect 4500 4968 4518 4986
rect 4500 4986 4518 5004
rect 4500 5004 4518 5022
rect 4500 5022 4518 5040
rect 4500 5040 4518 5058
rect 4500 5058 4518 5076
rect 4500 5076 4518 5094
rect 4500 5094 4518 5112
rect 4500 5112 4518 5130
rect 4500 5130 4518 5148
rect 4500 5148 4518 5166
rect 4500 5166 4518 5184
rect 4500 5184 4518 5202
rect 4500 5202 4518 5220
rect 4500 5220 4518 5238
rect 4500 5238 4518 5256
rect 4500 5256 4518 5274
rect 4500 5274 4518 5292
rect 4500 5292 4518 5310
rect 4500 5310 4518 5328
rect 4500 5328 4518 5346
rect 4500 5346 4518 5364
rect 4500 5364 4518 5382
rect 4500 5382 4518 5400
rect 4500 5400 4518 5418
rect 4500 5418 4518 5436
rect 4500 5436 4518 5454
rect 4500 5454 4518 5472
rect 4500 5472 4518 5490
rect 4500 5490 4518 5508
rect 4500 5508 4518 5526
rect 4500 5526 4518 5544
rect 4500 5544 4518 5562
rect 4500 5562 4518 5580
rect 4500 5580 4518 5598
rect 4500 5598 4518 5616
rect 4500 5616 4518 5634
rect 4500 5634 4518 5652
rect 4500 5652 4518 5670
rect 4500 5670 4518 5688
rect 4500 5688 4518 5706
rect 4500 5706 4518 5724
rect 4500 5724 4518 5742
rect 4500 5742 4518 5760
rect 4500 5760 4518 5778
rect 4500 5778 4518 5796
rect 4500 5796 4518 5814
rect 4500 5814 4518 5832
rect 4500 5832 4518 5850
rect 4500 5850 4518 5868
rect 4500 5868 4518 5886
rect 4500 5886 4518 5904
rect 4500 5904 4518 5922
rect 4500 5922 4518 5940
rect 4500 5940 4518 5958
rect 4500 5958 4518 5976
rect 4500 5976 4518 5994
rect 4500 5994 4518 6012
rect 4500 6012 4518 6030
rect 4500 6030 4518 6048
rect 4500 6048 4518 6066
rect 4500 6066 4518 6084
rect 4500 6084 4518 6102
rect 4500 6102 4518 6120
rect 4500 6120 4518 6138
rect 4500 6138 4518 6156
rect 4500 6156 4518 6174
rect 4500 6174 4518 6192
rect 4500 6192 4518 6210
rect 4500 6210 4518 6228
rect 4500 6228 4518 6246
rect 4500 6246 4518 6264
rect 4500 6264 4518 6282
rect 4500 6282 4518 6300
rect 4500 6300 4518 6318
rect 4500 6318 4518 6336
rect 4500 6336 4518 6354
rect 4500 6354 4518 6372
rect 4500 6372 4518 6390
rect 4500 6390 4518 6408
rect 4500 6408 4518 6426
rect 4500 6426 4518 6444
rect 4500 6444 4518 6462
rect 4500 6462 4518 6480
rect 4500 6480 4518 6498
rect 4500 6498 4518 6516
rect 4500 6516 4518 6534
rect 4500 6534 4518 6552
rect 4500 6552 4518 6570
rect 4500 6570 4518 6588
rect 4500 6588 4518 6606
rect 4500 6606 4518 6624
rect 4500 6624 4518 6642
rect 4500 6642 4518 6660
rect 4500 6660 4518 6678
rect 4500 6678 4518 6696
rect 4500 6696 4518 6714
rect 4500 6714 4518 6732
rect 4500 6732 4518 6750
rect 4500 6750 4518 6768
rect 4500 6768 4518 6786
rect 4500 6786 4518 6804
rect 4500 6804 4518 6822
rect 4500 6822 4518 6840
rect 4500 6840 4518 6858
rect 4500 6858 4518 6876
rect 4500 6876 4518 6894
rect 4500 6894 4518 6912
rect 4500 6912 4518 6930
rect 4500 6930 4518 6948
rect 4500 6948 4518 6966
rect 4500 6966 4518 6984
rect 4500 6984 4518 7002
rect 4500 7002 4518 7020
rect 4500 7020 4518 7038
rect 4518 108 4536 126
rect 4518 126 4536 144
rect 4518 144 4536 162
rect 4518 162 4536 180
rect 4518 180 4536 198
rect 4518 198 4536 216
rect 4518 216 4536 234
rect 4518 234 4536 252
rect 4518 252 4536 270
rect 4518 270 4536 288
rect 4518 288 4536 306
rect 4518 306 4536 324
rect 4518 324 4536 342
rect 4518 342 4536 360
rect 4518 360 4536 378
rect 4518 378 4536 396
rect 4518 396 4536 414
rect 4518 414 4536 432
rect 4518 432 4536 450
rect 4518 450 4536 468
rect 4518 468 4536 486
rect 4518 486 4536 504
rect 4518 504 4536 522
rect 4518 522 4536 540
rect 4518 540 4536 558
rect 4518 558 4536 576
rect 4518 576 4536 594
rect 4518 594 4536 612
rect 4518 612 4536 630
rect 4518 630 4536 648
rect 4518 648 4536 666
rect 4518 666 4536 684
rect 4518 684 4536 702
rect 4518 702 4536 720
rect 4518 720 4536 738
rect 4518 738 4536 756
rect 4518 864 4536 882
rect 4518 882 4536 900
rect 4518 900 4536 918
rect 4518 918 4536 936
rect 4518 936 4536 954
rect 4518 954 4536 972
rect 4518 972 4536 990
rect 4518 990 4536 1008
rect 4518 1008 4536 1026
rect 4518 1026 4536 1044
rect 4518 1044 4536 1062
rect 4518 1062 4536 1080
rect 4518 1080 4536 1098
rect 4518 1098 4536 1116
rect 4518 1116 4536 1134
rect 4518 1134 4536 1152
rect 4518 1152 4536 1170
rect 4518 1170 4536 1188
rect 4518 1188 4536 1206
rect 4518 1206 4536 1224
rect 4518 1224 4536 1242
rect 4518 1242 4536 1260
rect 4518 1260 4536 1278
rect 4518 1278 4536 1296
rect 4518 1296 4536 1314
rect 4518 1314 4536 1332
rect 4518 1332 4536 1350
rect 4518 1350 4536 1368
rect 4518 1368 4536 1386
rect 4518 1386 4536 1404
rect 4518 1404 4536 1422
rect 4518 1422 4536 1440
rect 4518 1440 4536 1458
rect 4518 1458 4536 1476
rect 4518 1476 4536 1494
rect 4518 1494 4536 1512
rect 4518 1512 4536 1530
rect 4518 1530 4536 1548
rect 4518 1548 4536 1566
rect 4518 1566 4536 1584
rect 4518 1584 4536 1602
rect 4518 1602 4536 1620
rect 4518 1620 4536 1638
rect 4518 1638 4536 1656
rect 4518 1656 4536 1674
rect 4518 1674 4536 1692
rect 4518 1692 4536 1710
rect 4518 1710 4536 1728
rect 4518 1728 4536 1746
rect 4518 1746 4536 1764
rect 4518 1764 4536 1782
rect 4518 1782 4536 1800
rect 4518 1800 4536 1818
rect 4518 1818 4536 1836
rect 4518 1836 4536 1854
rect 4518 1854 4536 1872
rect 4518 1872 4536 1890
rect 4518 1890 4536 1908
rect 4518 2142 4536 2160
rect 4518 2160 4536 2178
rect 4518 2178 4536 2196
rect 4518 2196 4536 2214
rect 4518 2214 4536 2232
rect 4518 2232 4536 2250
rect 4518 2250 4536 2268
rect 4518 2268 4536 2286
rect 4518 2286 4536 2304
rect 4518 2304 4536 2322
rect 4518 2322 4536 2340
rect 4518 2340 4536 2358
rect 4518 2358 4536 2376
rect 4518 2376 4536 2394
rect 4518 2394 4536 2412
rect 4518 2412 4536 2430
rect 4518 2430 4536 2448
rect 4518 2448 4536 2466
rect 4518 2466 4536 2484
rect 4518 2484 4536 2502
rect 4518 2502 4536 2520
rect 4518 2520 4536 2538
rect 4518 2538 4536 2556
rect 4518 2556 4536 2574
rect 4518 2574 4536 2592
rect 4518 2592 4536 2610
rect 4518 2610 4536 2628
rect 4518 2628 4536 2646
rect 4518 2646 4536 2664
rect 4518 2664 4536 2682
rect 4518 2682 4536 2700
rect 4518 2700 4536 2718
rect 4518 2718 4536 2736
rect 4518 2736 4536 2754
rect 4518 2754 4536 2772
rect 4518 2772 4536 2790
rect 4518 2790 4536 2808
rect 4518 2808 4536 2826
rect 4518 2826 4536 2844
rect 4518 2844 4536 2862
rect 4518 2862 4536 2880
rect 4518 2880 4536 2898
rect 4518 2898 4536 2916
rect 4518 2916 4536 2934
rect 4518 2934 4536 2952
rect 4518 2952 4536 2970
rect 4518 2970 4536 2988
rect 4518 2988 4536 3006
rect 4518 3006 4536 3024
rect 4518 3024 4536 3042
rect 4518 3042 4536 3060
rect 4518 3060 4536 3078
rect 4518 3078 4536 3096
rect 4518 3096 4536 3114
rect 4518 3114 4536 3132
rect 4518 3132 4536 3150
rect 4518 3150 4536 3168
rect 4518 3168 4536 3186
rect 4518 3186 4536 3204
rect 4518 3204 4536 3222
rect 4518 3222 4536 3240
rect 4518 3240 4536 3258
rect 4518 3258 4536 3276
rect 4518 3276 4536 3294
rect 4518 3294 4536 3312
rect 4518 3312 4536 3330
rect 4518 3330 4536 3348
rect 4518 3348 4536 3366
rect 4518 3366 4536 3384
rect 4518 3384 4536 3402
rect 4518 3402 4536 3420
rect 4518 3420 4536 3438
rect 4518 3438 4536 3456
rect 4518 3456 4536 3474
rect 4518 3474 4536 3492
rect 4518 3492 4536 3510
rect 4518 3510 4536 3528
rect 4518 3528 4536 3546
rect 4518 3546 4536 3564
rect 4518 3564 4536 3582
rect 4518 3582 4536 3600
rect 4518 3600 4536 3618
rect 4518 3618 4536 3636
rect 4518 3636 4536 3654
rect 4518 3654 4536 3672
rect 4518 3672 4536 3690
rect 4518 3690 4536 3708
rect 4518 3708 4536 3726
rect 4518 3726 4536 3744
rect 4518 3744 4536 3762
rect 4518 3762 4536 3780
rect 4518 3780 4536 3798
rect 4518 3798 4536 3816
rect 4518 4014 4536 4032
rect 4518 4032 4536 4050
rect 4518 4050 4536 4068
rect 4518 4068 4536 4086
rect 4518 4086 4536 4104
rect 4518 4104 4536 4122
rect 4518 4122 4536 4140
rect 4518 4140 4536 4158
rect 4518 4158 4536 4176
rect 4518 4176 4536 4194
rect 4518 4194 4536 4212
rect 4518 4212 4536 4230
rect 4518 4230 4536 4248
rect 4518 4248 4536 4266
rect 4518 4266 4536 4284
rect 4518 4284 4536 4302
rect 4518 4302 4536 4320
rect 4518 4320 4536 4338
rect 4518 4338 4536 4356
rect 4518 4356 4536 4374
rect 4518 4374 4536 4392
rect 4518 4392 4536 4410
rect 4518 4410 4536 4428
rect 4518 4428 4536 4446
rect 4518 4446 4536 4464
rect 4518 4464 4536 4482
rect 4518 4482 4536 4500
rect 4518 4500 4536 4518
rect 4518 4518 4536 4536
rect 4518 4536 4536 4554
rect 4518 4554 4536 4572
rect 4518 4572 4536 4590
rect 4518 4590 4536 4608
rect 4518 4608 4536 4626
rect 4518 4626 4536 4644
rect 4518 4644 4536 4662
rect 4518 4662 4536 4680
rect 4518 4680 4536 4698
rect 4518 4698 4536 4716
rect 4518 4716 4536 4734
rect 4518 4734 4536 4752
rect 4518 4752 4536 4770
rect 4518 4770 4536 4788
rect 4518 4788 4536 4806
rect 4518 4806 4536 4824
rect 4518 4824 4536 4842
rect 4518 4842 4536 4860
rect 4518 4860 4536 4878
rect 4518 4878 4536 4896
rect 4518 4896 4536 4914
rect 4518 4914 4536 4932
rect 4518 4932 4536 4950
rect 4518 4950 4536 4968
rect 4518 4968 4536 4986
rect 4518 4986 4536 5004
rect 4518 5004 4536 5022
rect 4518 5022 4536 5040
rect 4518 5040 4536 5058
rect 4518 5058 4536 5076
rect 4518 5076 4536 5094
rect 4518 5094 4536 5112
rect 4518 5112 4536 5130
rect 4518 5130 4536 5148
rect 4518 5148 4536 5166
rect 4518 5166 4536 5184
rect 4518 5184 4536 5202
rect 4518 5202 4536 5220
rect 4518 5220 4536 5238
rect 4518 5238 4536 5256
rect 4518 5256 4536 5274
rect 4518 5274 4536 5292
rect 4518 5292 4536 5310
rect 4518 5310 4536 5328
rect 4518 5328 4536 5346
rect 4518 5346 4536 5364
rect 4518 5364 4536 5382
rect 4518 5382 4536 5400
rect 4518 5400 4536 5418
rect 4518 5418 4536 5436
rect 4518 5436 4536 5454
rect 4518 5454 4536 5472
rect 4518 5472 4536 5490
rect 4518 5490 4536 5508
rect 4518 5508 4536 5526
rect 4518 5526 4536 5544
rect 4518 5544 4536 5562
rect 4518 5562 4536 5580
rect 4518 5580 4536 5598
rect 4518 5598 4536 5616
rect 4518 5616 4536 5634
rect 4518 5634 4536 5652
rect 4518 5652 4536 5670
rect 4518 5670 4536 5688
rect 4518 5688 4536 5706
rect 4518 5706 4536 5724
rect 4518 5724 4536 5742
rect 4518 5742 4536 5760
rect 4518 5760 4536 5778
rect 4518 5778 4536 5796
rect 4518 5796 4536 5814
rect 4518 5814 4536 5832
rect 4518 5832 4536 5850
rect 4518 5850 4536 5868
rect 4518 5868 4536 5886
rect 4518 5886 4536 5904
rect 4518 5904 4536 5922
rect 4518 5922 4536 5940
rect 4518 5940 4536 5958
rect 4518 5958 4536 5976
rect 4518 5976 4536 5994
rect 4518 5994 4536 6012
rect 4518 6012 4536 6030
rect 4518 6030 4536 6048
rect 4518 6048 4536 6066
rect 4518 6066 4536 6084
rect 4518 6084 4536 6102
rect 4518 6102 4536 6120
rect 4518 6120 4536 6138
rect 4518 6138 4536 6156
rect 4518 6156 4536 6174
rect 4518 6174 4536 6192
rect 4518 6192 4536 6210
rect 4518 6210 4536 6228
rect 4518 6228 4536 6246
rect 4518 6246 4536 6264
rect 4518 6264 4536 6282
rect 4518 6282 4536 6300
rect 4518 6300 4536 6318
rect 4518 6318 4536 6336
rect 4518 6336 4536 6354
rect 4518 6354 4536 6372
rect 4518 6372 4536 6390
rect 4518 6390 4536 6408
rect 4518 6408 4536 6426
rect 4518 6426 4536 6444
rect 4518 6444 4536 6462
rect 4518 6462 4536 6480
rect 4518 6480 4536 6498
rect 4518 6498 4536 6516
rect 4518 6516 4536 6534
rect 4518 6534 4536 6552
rect 4518 6552 4536 6570
rect 4518 6570 4536 6588
rect 4518 6588 4536 6606
rect 4518 6606 4536 6624
rect 4518 6624 4536 6642
rect 4518 6642 4536 6660
rect 4518 6660 4536 6678
rect 4518 6678 4536 6696
rect 4518 6696 4536 6714
rect 4518 6714 4536 6732
rect 4518 6732 4536 6750
rect 4518 6750 4536 6768
rect 4518 6768 4536 6786
rect 4518 6786 4536 6804
rect 4518 6804 4536 6822
rect 4518 6822 4536 6840
rect 4518 6840 4536 6858
rect 4518 6858 4536 6876
rect 4518 6876 4536 6894
rect 4518 6894 4536 6912
rect 4518 6912 4536 6930
rect 4518 6930 4536 6948
rect 4518 6948 4536 6966
rect 4518 6966 4536 6984
rect 4518 6984 4536 7002
rect 4518 7002 4536 7020
rect 4518 7020 4536 7038
rect 4518 7038 4536 7056
rect 4518 7056 4536 7074
rect 4536 108 4554 126
rect 4536 126 4554 144
rect 4536 144 4554 162
rect 4536 162 4554 180
rect 4536 180 4554 198
rect 4536 198 4554 216
rect 4536 216 4554 234
rect 4536 234 4554 252
rect 4536 252 4554 270
rect 4536 270 4554 288
rect 4536 288 4554 306
rect 4536 306 4554 324
rect 4536 324 4554 342
rect 4536 342 4554 360
rect 4536 360 4554 378
rect 4536 378 4554 396
rect 4536 396 4554 414
rect 4536 414 4554 432
rect 4536 432 4554 450
rect 4536 450 4554 468
rect 4536 468 4554 486
rect 4536 486 4554 504
rect 4536 504 4554 522
rect 4536 522 4554 540
rect 4536 540 4554 558
rect 4536 558 4554 576
rect 4536 576 4554 594
rect 4536 594 4554 612
rect 4536 612 4554 630
rect 4536 630 4554 648
rect 4536 648 4554 666
rect 4536 666 4554 684
rect 4536 684 4554 702
rect 4536 702 4554 720
rect 4536 720 4554 738
rect 4536 738 4554 756
rect 4536 864 4554 882
rect 4536 882 4554 900
rect 4536 900 4554 918
rect 4536 918 4554 936
rect 4536 936 4554 954
rect 4536 954 4554 972
rect 4536 972 4554 990
rect 4536 990 4554 1008
rect 4536 1008 4554 1026
rect 4536 1026 4554 1044
rect 4536 1044 4554 1062
rect 4536 1062 4554 1080
rect 4536 1080 4554 1098
rect 4536 1098 4554 1116
rect 4536 1116 4554 1134
rect 4536 1134 4554 1152
rect 4536 1152 4554 1170
rect 4536 1170 4554 1188
rect 4536 1188 4554 1206
rect 4536 1206 4554 1224
rect 4536 1224 4554 1242
rect 4536 1242 4554 1260
rect 4536 1260 4554 1278
rect 4536 1278 4554 1296
rect 4536 1296 4554 1314
rect 4536 1314 4554 1332
rect 4536 1332 4554 1350
rect 4536 1350 4554 1368
rect 4536 1368 4554 1386
rect 4536 1386 4554 1404
rect 4536 1404 4554 1422
rect 4536 1422 4554 1440
rect 4536 1440 4554 1458
rect 4536 1458 4554 1476
rect 4536 1476 4554 1494
rect 4536 1494 4554 1512
rect 4536 1512 4554 1530
rect 4536 1530 4554 1548
rect 4536 1548 4554 1566
rect 4536 1566 4554 1584
rect 4536 1584 4554 1602
rect 4536 1602 4554 1620
rect 4536 1620 4554 1638
rect 4536 1638 4554 1656
rect 4536 1656 4554 1674
rect 4536 1674 4554 1692
rect 4536 1692 4554 1710
rect 4536 1710 4554 1728
rect 4536 1728 4554 1746
rect 4536 1746 4554 1764
rect 4536 1764 4554 1782
rect 4536 1782 4554 1800
rect 4536 1800 4554 1818
rect 4536 1818 4554 1836
rect 4536 1836 4554 1854
rect 4536 1854 4554 1872
rect 4536 1872 4554 1890
rect 4536 1890 4554 1908
rect 4536 1908 4554 1926
rect 4536 2160 4554 2178
rect 4536 2178 4554 2196
rect 4536 2196 4554 2214
rect 4536 2214 4554 2232
rect 4536 2232 4554 2250
rect 4536 2250 4554 2268
rect 4536 2268 4554 2286
rect 4536 2286 4554 2304
rect 4536 2304 4554 2322
rect 4536 2322 4554 2340
rect 4536 2340 4554 2358
rect 4536 2358 4554 2376
rect 4536 2376 4554 2394
rect 4536 2394 4554 2412
rect 4536 2412 4554 2430
rect 4536 2430 4554 2448
rect 4536 2448 4554 2466
rect 4536 2466 4554 2484
rect 4536 2484 4554 2502
rect 4536 2502 4554 2520
rect 4536 2520 4554 2538
rect 4536 2538 4554 2556
rect 4536 2556 4554 2574
rect 4536 2574 4554 2592
rect 4536 2592 4554 2610
rect 4536 2610 4554 2628
rect 4536 2628 4554 2646
rect 4536 2646 4554 2664
rect 4536 2664 4554 2682
rect 4536 2682 4554 2700
rect 4536 2700 4554 2718
rect 4536 2718 4554 2736
rect 4536 2736 4554 2754
rect 4536 2754 4554 2772
rect 4536 2772 4554 2790
rect 4536 2790 4554 2808
rect 4536 2808 4554 2826
rect 4536 2826 4554 2844
rect 4536 2844 4554 2862
rect 4536 2862 4554 2880
rect 4536 2880 4554 2898
rect 4536 2898 4554 2916
rect 4536 2916 4554 2934
rect 4536 2934 4554 2952
rect 4536 2952 4554 2970
rect 4536 2970 4554 2988
rect 4536 2988 4554 3006
rect 4536 3006 4554 3024
rect 4536 3024 4554 3042
rect 4536 3042 4554 3060
rect 4536 3060 4554 3078
rect 4536 3078 4554 3096
rect 4536 3096 4554 3114
rect 4536 3114 4554 3132
rect 4536 3132 4554 3150
rect 4536 3150 4554 3168
rect 4536 3168 4554 3186
rect 4536 3186 4554 3204
rect 4536 3204 4554 3222
rect 4536 3222 4554 3240
rect 4536 3240 4554 3258
rect 4536 3258 4554 3276
rect 4536 3276 4554 3294
rect 4536 3294 4554 3312
rect 4536 3312 4554 3330
rect 4536 3330 4554 3348
rect 4536 3348 4554 3366
rect 4536 3366 4554 3384
rect 4536 3384 4554 3402
rect 4536 3402 4554 3420
rect 4536 3420 4554 3438
rect 4536 3438 4554 3456
rect 4536 3456 4554 3474
rect 4536 3474 4554 3492
rect 4536 3492 4554 3510
rect 4536 3510 4554 3528
rect 4536 3528 4554 3546
rect 4536 3546 4554 3564
rect 4536 3564 4554 3582
rect 4536 3582 4554 3600
rect 4536 3600 4554 3618
rect 4536 3618 4554 3636
rect 4536 3636 4554 3654
rect 4536 3654 4554 3672
rect 4536 3672 4554 3690
rect 4536 3690 4554 3708
rect 4536 3708 4554 3726
rect 4536 3726 4554 3744
rect 4536 3744 4554 3762
rect 4536 3762 4554 3780
rect 4536 3780 4554 3798
rect 4536 3798 4554 3816
rect 4536 3816 4554 3834
rect 4536 4050 4554 4068
rect 4536 4068 4554 4086
rect 4536 4086 4554 4104
rect 4536 4104 4554 4122
rect 4536 4122 4554 4140
rect 4536 4140 4554 4158
rect 4536 4158 4554 4176
rect 4536 4176 4554 4194
rect 4536 4194 4554 4212
rect 4536 4212 4554 4230
rect 4536 4230 4554 4248
rect 4536 4248 4554 4266
rect 4536 4266 4554 4284
rect 4536 4284 4554 4302
rect 4536 4302 4554 4320
rect 4536 4320 4554 4338
rect 4536 4338 4554 4356
rect 4536 4356 4554 4374
rect 4536 4374 4554 4392
rect 4536 4392 4554 4410
rect 4536 4410 4554 4428
rect 4536 4428 4554 4446
rect 4536 4446 4554 4464
rect 4536 4464 4554 4482
rect 4536 4482 4554 4500
rect 4536 4500 4554 4518
rect 4536 4518 4554 4536
rect 4536 4536 4554 4554
rect 4536 4554 4554 4572
rect 4536 4572 4554 4590
rect 4536 4590 4554 4608
rect 4536 4608 4554 4626
rect 4536 4626 4554 4644
rect 4536 4644 4554 4662
rect 4536 4662 4554 4680
rect 4536 4680 4554 4698
rect 4536 4698 4554 4716
rect 4536 4716 4554 4734
rect 4536 4734 4554 4752
rect 4536 4752 4554 4770
rect 4536 4770 4554 4788
rect 4536 4788 4554 4806
rect 4536 4806 4554 4824
rect 4536 4824 4554 4842
rect 4536 4842 4554 4860
rect 4536 4860 4554 4878
rect 4536 4878 4554 4896
rect 4536 4896 4554 4914
rect 4536 4914 4554 4932
rect 4536 4932 4554 4950
rect 4536 4950 4554 4968
rect 4536 4968 4554 4986
rect 4536 4986 4554 5004
rect 4536 5004 4554 5022
rect 4536 5022 4554 5040
rect 4536 5040 4554 5058
rect 4536 5058 4554 5076
rect 4536 5076 4554 5094
rect 4536 5094 4554 5112
rect 4536 5112 4554 5130
rect 4536 5130 4554 5148
rect 4536 5148 4554 5166
rect 4536 5166 4554 5184
rect 4536 5184 4554 5202
rect 4536 5202 4554 5220
rect 4536 5220 4554 5238
rect 4536 5238 4554 5256
rect 4536 5256 4554 5274
rect 4536 5274 4554 5292
rect 4536 5292 4554 5310
rect 4536 5310 4554 5328
rect 4536 5328 4554 5346
rect 4536 5346 4554 5364
rect 4536 5364 4554 5382
rect 4536 5382 4554 5400
rect 4536 5400 4554 5418
rect 4536 5418 4554 5436
rect 4536 5436 4554 5454
rect 4536 5454 4554 5472
rect 4536 5472 4554 5490
rect 4536 5490 4554 5508
rect 4536 5508 4554 5526
rect 4536 5526 4554 5544
rect 4536 5544 4554 5562
rect 4536 5562 4554 5580
rect 4536 5580 4554 5598
rect 4536 5598 4554 5616
rect 4536 5616 4554 5634
rect 4536 5634 4554 5652
rect 4536 5652 4554 5670
rect 4536 5670 4554 5688
rect 4536 5688 4554 5706
rect 4536 5706 4554 5724
rect 4536 5724 4554 5742
rect 4536 5742 4554 5760
rect 4536 5760 4554 5778
rect 4536 5778 4554 5796
rect 4536 5796 4554 5814
rect 4536 5814 4554 5832
rect 4536 5832 4554 5850
rect 4536 5850 4554 5868
rect 4536 5868 4554 5886
rect 4536 5886 4554 5904
rect 4536 5904 4554 5922
rect 4536 5922 4554 5940
rect 4536 5940 4554 5958
rect 4536 5958 4554 5976
rect 4536 5976 4554 5994
rect 4536 5994 4554 6012
rect 4536 6012 4554 6030
rect 4536 6030 4554 6048
rect 4536 6048 4554 6066
rect 4536 6066 4554 6084
rect 4536 6084 4554 6102
rect 4536 6102 4554 6120
rect 4536 6120 4554 6138
rect 4536 6138 4554 6156
rect 4536 6156 4554 6174
rect 4536 6174 4554 6192
rect 4536 6192 4554 6210
rect 4536 6210 4554 6228
rect 4536 6228 4554 6246
rect 4536 6246 4554 6264
rect 4536 6264 4554 6282
rect 4536 6282 4554 6300
rect 4536 6300 4554 6318
rect 4536 6318 4554 6336
rect 4536 6336 4554 6354
rect 4536 6354 4554 6372
rect 4536 6372 4554 6390
rect 4536 6390 4554 6408
rect 4536 6408 4554 6426
rect 4536 6426 4554 6444
rect 4536 6444 4554 6462
rect 4536 6462 4554 6480
rect 4536 6480 4554 6498
rect 4536 6498 4554 6516
rect 4536 6516 4554 6534
rect 4536 6534 4554 6552
rect 4536 6552 4554 6570
rect 4536 6570 4554 6588
rect 4536 6588 4554 6606
rect 4536 6606 4554 6624
rect 4536 6624 4554 6642
rect 4536 6642 4554 6660
rect 4536 6660 4554 6678
rect 4536 6678 4554 6696
rect 4536 6696 4554 6714
rect 4536 6714 4554 6732
rect 4536 6732 4554 6750
rect 4536 6750 4554 6768
rect 4536 6768 4554 6786
rect 4536 6786 4554 6804
rect 4536 6804 4554 6822
rect 4536 6822 4554 6840
rect 4536 6840 4554 6858
rect 4536 6858 4554 6876
rect 4536 6876 4554 6894
rect 4536 6894 4554 6912
rect 4536 6912 4554 6930
rect 4536 6930 4554 6948
rect 4536 6948 4554 6966
rect 4536 6966 4554 6984
rect 4536 6984 4554 7002
rect 4536 7002 4554 7020
rect 4536 7020 4554 7038
rect 4536 7038 4554 7056
rect 4536 7056 4554 7074
rect 4536 7074 4554 7092
rect 4536 7092 4554 7110
rect 4554 108 4572 126
rect 4554 126 4572 144
rect 4554 144 4572 162
rect 4554 162 4572 180
rect 4554 180 4572 198
rect 4554 198 4572 216
rect 4554 216 4572 234
rect 4554 234 4572 252
rect 4554 252 4572 270
rect 4554 270 4572 288
rect 4554 288 4572 306
rect 4554 306 4572 324
rect 4554 324 4572 342
rect 4554 342 4572 360
rect 4554 360 4572 378
rect 4554 378 4572 396
rect 4554 396 4572 414
rect 4554 414 4572 432
rect 4554 432 4572 450
rect 4554 450 4572 468
rect 4554 468 4572 486
rect 4554 486 4572 504
rect 4554 504 4572 522
rect 4554 522 4572 540
rect 4554 540 4572 558
rect 4554 558 4572 576
rect 4554 576 4572 594
rect 4554 594 4572 612
rect 4554 612 4572 630
rect 4554 630 4572 648
rect 4554 648 4572 666
rect 4554 666 4572 684
rect 4554 684 4572 702
rect 4554 702 4572 720
rect 4554 720 4572 738
rect 4554 738 4572 756
rect 4554 864 4572 882
rect 4554 882 4572 900
rect 4554 900 4572 918
rect 4554 918 4572 936
rect 4554 936 4572 954
rect 4554 954 4572 972
rect 4554 972 4572 990
rect 4554 990 4572 1008
rect 4554 1008 4572 1026
rect 4554 1026 4572 1044
rect 4554 1044 4572 1062
rect 4554 1062 4572 1080
rect 4554 1080 4572 1098
rect 4554 1098 4572 1116
rect 4554 1116 4572 1134
rect 4554 1134 4572 1152
rect 4554 1152 4572 1170
rect 4554 1170 4572 1188
rect 4554 1188 4572 1206
rect 4554 1206 4572 1224
rect 4554 1224 4572 1242
rect 4554 1242 4572 1260
rect 4554 1260 4572 1278
rect 4554 1278 4572 1296
rect 4554 1296 4572 1314
rect 4554 1314 4572 1332
rect 4554 1332 4572 1350
rect 4554 1350 4572 1368
rect 4554 1368 4572 1386
rect 4554 1386 4572 1404
rect 4554 1404 4572 1422
rect 4554 1422 4572 1440
rect 4554 1440 4572 1458
rect 4554 1458 4572 1476
rect 4554 1476 4572 1494
rect 4554 1494 4572 1512
rect 4554 1512 4572 1530
rect 4554 1530 4572 1548
rect 4554 1548 4572 1566
rect 4554 1566 4572 1584
rect 4554 1584 4572 1602
rect 4554 1602 4572 1620
rect 4554 1620 4572 1638
rect 4554 1638 4572 1656
rect 4554 1656 4572 1674
rect 4554 1674 4572 1692
rect 4554 1692 4572 1710
rect 4554 1710 4572 1728
rect 4554 1728 4572 1746
rect 4554 1746 4572 1764
rect 4554 1764 4572 1782
rect 4554 1782 4572 1800
rect 4554 1800 4572 1818
rect 4554 1818 4572 1836
rect 4554 1836 4572 1854
rect 4554 1854 4572 1872
rect 4554 1872 4572 1890
rect 4554 1890 4572 1908
rect 4554 1908 4572 1926
rect 4554 1926 4572 1944
rect 4554 2178 4572 2196
rect 4554 2196 4572 2214
rect 4554 2214 4572 2232
rect 4554 2232 4572 2250
rect 4554 2250 4572 2268
rect 4554 2268 4572 2286
rect 4554 2286 4572 2304
rect 4554 2304 4572 2322
rect 4554 2322 4572 2340
rect 4554 2340 4572 2358
rect 4554 2358 4572 2376
rect 4554 2376 4572 2394
rect 4554 2394 4572 2412
rect 4554 2412 4572 2430
rect 4554 2430 4572 2448
rect 4554 2448 4572 2466
rect 4554 2466 4572 2484
rect 4554 2484 4572 2502
rect 4554 2502 4572 2520
rect 4554 2520 4572 2538
rect 4554 2538 4572 2556
rect 4554 2556 4572 2574
rect 4554 2574 4572 2592
rect 4554 2592 4572 2610
rect 4554 2610 4572 2628
rect 4554 2628 4572 2646
rect 4554 2646 4572 2664
rect 4554 2664 4572 2682
rect 4554 2682 4572 2700
rect 4554 2700 4572 2718
rect 4554 2718 4572 2736
rect 4554 2736 4572 2754
rect 4554 2754 4572 2772
rect 4554 2772 4572 2790
rect 4554 2790 4572 2808
rect 4554 2808 4572 2826
rect 4554 2826 4572 2844
rect 4554 2844 4572 2862
rect 4554 2862 4572 2880
rect 4554 2880 4572 2898
rect 4554 2898 4572 2916
rect 4554 2916 4572 2934
rect 4554 2934 4572 2952
rect 4554 2952 4572 2970
rect 4554 2970 4572 2988
rect 4554 2988 4572 3006
rect 4554 3006 4572 3024
rect 4554 3024 4572 3042
rect 4554 3042 4572 3060
rect 4554 3060 4572 3078
rect 4554 3078 4572 3096
rect 4554 3096 4572 3114
rect 4554 3114 4572 3132
rect 4554 3132 4572 3150
rect 4554 3150 4572 3168
rect 4554 3168 4572 3186
rect 4554 3186 4572 3204
rect 4554 3204 4572 3222
rect 4554 3222 4572 3240
rect 4554 3240 4572 3258
rect 4554 3258 4572 3276
rect 4554 3276 4572 3294
rect 4554 3294 4572 3312
rect 4554 3312 4572 3330
rect 4554 3330 4572 3348
rect 4554 3348 4572 3366
rect 4554 3366 4572 3384
rect 4554 3384 4572 3402
rect 4554 3402 4572 3420
rect 4554 3420 4572 3438
rect 4554 3438 4572 3456
rect 4554 3456 4572 3474
rect 4554 3474 4572 3492
rect 4554 3492 4572 3510
rect 4554 3510 4572 3528
rect 4554 3528 4572 3546
rect 4554 3546 4572 3564
rect 4554 3564 4572 3582
rect 4554 3582 4572 3600
rect 4554 3600 4572 3618
rect 4554 3618 4572 3636
rect 4554 3636 4572 3654
rect 4554 3654 4572 3672
rect 4554 3672 4572 3690
rect 4554 3690 4572 3708
rect 4554 3708 4572 3726
rect 4554 3726 4572 3744
rect 4554 3744 4572 3762
rect 4554 3762 4572 3780
rect 4554 3780 4572 3798
rect 4554 3798 4572 3816
rect 4554 3816 4572 3834
rect 4554 3834 4572 3852
rect 4554 3852 4572 3870
rect 4554 4068 4572 4086
rect 4554 4086 4572 4104
rect 4554 4104 4572 4122
rect 4554 4122 4572 4140
rect 4554 4140 4572 4158
rect 4554 4158 4572 4176
rect 4554 4176 4572 4194
rect 4554 4194 4572 4212
rect 4554 4212 4572 4230
rect 4554 4230 4572 4248
rect 4554 4248 4572 4266
rect 4554 4266 4572 4284
rect 4554 4284 4572 4302
rect 4554 4302 4572 4320
rect 4554 4320 4572 4338
rect 4554 4338 4572 4356
rect 4554 4356 4572 4374
rect 4554 4374 4572 4392
rect 4554 4392 4572 4410
rect 4554 4410 4572 4428
rect 4554 4428 4572 4446
rect 4554 4446 4572 4464
rect 4554 4464 4572 4482
rect 4554 4482 4572 4500
rect 4554 4500 4572 4518
rect 4554 4518 4572 4536
rect 4554 4536 4572 4554
rect 4554 4554 4572 4572
rect 4554 4572 4572 4590
rect 4554 4590 4572 4608
rect 4554 4608 4572 4626
rect 4554 4626 4572 4644
rect 4554 4644 4572 4662
rect 4554 4662 4572 4680
rect 4554 4680 4572 4698
rect 4554 4698 4572 4716
rect 4554 4716 4572 4734
rect 4554 4734 4572 4752
rect 4554 4752 4572 4770
rect 4554 4770 4572 4788
rect 4554 4788 4572 4806
rect 4554 4806 4572 4824
rect 4554 4824 4572 4842
rect 4554 4842 4572 4860
rect 4554 4860 4572 4878
rect 4554 4878 4572 4896
rect 4554 4896 4572 4914
rect 4554 4914 4572 4932
rect 4554 4932 4572 4950
rect 4554 4950 4572 4968
rect 4554 4968 4572 4986
rect 4554 4986 4572 5004
rect 4554 5004 4572 5022
rect 4554 5022 4572 5040
rect 4554 5040 4572 5058
rect 4554 5058 4572 5076
rect 4554 5076 4572 5094
rect 4554 5094 4572 5112
rect 4554 5112 4572 5130
rect 4554 5130 4572 5148
rect 4554 5148 4572 5166
rect 4554 5166 4572 5184
rect 4554 5184 4572 5202
rect 4554 5202 4572 5220
rect 4554 5220 4572 5238
rect 4554 5238 4572 5256
rect 4554 5256 4572 5274
rect 4554 5274 4572 5292
rect 4554 5292 4572 5310
rect 4554 5310 4572 5328
rect 4554 5328 4572 5346
rect 4554 5346 4572 5364
rect 4554 5364 4572 5382
rect 4554 5382 4572 5400
rect 4554 5400 4572 5418
rect 4554 5418 4572 5436
rect 4554 5436 4572 5454
rect 4554 5454 4572 5472
rect 4554 5472 4572 5490
rect 4554 5490 4572 5508
rect 4554 5508 4572 5526
rect 4554 5526 4572 5544
rect 4554 5544 4572 5562
rect 4554 5562 4572 5580
rect 4554 5580 4572 5598
rect 4554 5598 4572 5616
rect 4554 5616 4572 5634
rect 4554 5634 4572 5652
rect 4554 5652 4572 5670
rect 4554 5670 4572 5688
rect 4554 5688 4572 5706
rect 4554 5706 4572 5724
rect 4554 5724 4572 5742
rect 4554 5742 4572 5760
rect 4554 5760 4572 5778
rect 4554 5778 4572 5796
rect 4554 5796 4572 5814
rect 4554 5814 4572 5832
rect 4554 5832 4572 5850
rect 4554 5850 4572 5868
rect 4554 5868 4572 5886
rect 4554 5886 4572 5904
rect 4554 5904 4572 5922
rect 4554 5922 4572 5940
rect 4554 5940 4572 5958
rect 4554 5958 4572 5976
rect 4554 5976 4572 5994
rect 4554 5994 4572 6012
rect 4554 6012 4572 6030
rect 4554 6030 4572 6048
rect 4554 6048 4572 6066
rect 4554 6066 4572 6084
rect 4554 6084 4572 6102
rect 4554 6102 4572 6120
rect 4554 6120 4572 6138
rect 4554 6138 4572 6156
rect 4554 6156 4572 6174
rect 4554 6174 4572 6192
rect 4554 6192 4572 6210
rect 4554 6210 4572 6228
rect 4554 6228 4572 6246
rect 4554 6246 4572 6264
rect 4554 6264 4572 6282
rect 4554 6282 4572 6300
rect 4554 6300 4572 6318
rect 4554 6318 4572 6336
rect 4554 6336 4572 6354
rect 4554 6354 4572 6372
rect 4554 6372 4572 6390
rect 4554 6390 4572 6408
rect 4554 6408 4572 6426
rect 4554 6426 4572 6444
rect 4554 6444 4572 6462
rect 4554 6462 4572 6480
rect 4554 6480 4572 6498
rect 4554 6498 4572 6516
rect 4554 6516 4572 6534
rect 4554 6534 4572 6552
rect 4554 6552 4572 6570
rect 4554 6570 4572 6588
rect 4554 6588 4572 6606
rect 4554 6606 4572 6624
rect 4554 6624 4572 6642
rect 4554 6642 4572 6660
rect 4554 6660 4572 6678
rect 4554 6678 4572 6696
rect 4554 6696 4572 6714
rect 4554 6714 4572 6732
rect 4554 6732 4572 6750
rect 4554 6750 4572 6768
rect 4554 6768 4572 6786
rect 4554 6786 4572 6804
rect 4554 6804 4572 6822
rect 4554 6822 4572 6840
rect 4554 6840 4572 6858
rect 4554 6858 4572 6876
rect 4554 6876 4572 6894
rect 4554 6894 4572 6912
rect 4554 6912 4572 6930
rect 4554 6930 4572 6948
rect 4554 6948 4572 6966
rect 4554 6966 4572 6984
rect 4554 6984 4572 7002
rect 4554 7002 4572 7020
rect 4554 7020 4572 7038
rect 4554 7038 4572 7056
rect 4554 7056 4572 7074
rect 4554 7074 4572 7092
rect 4554 7092 4572 7110
rect 4554 7110 4572 7128
rect 4572 126 4590 144
rect 4572 144 4590 162
rect 4572 162 4590 180
rect 4572 180 4590 198
rect 4572 198 4590 216
rect 4572 216 4590 234
rect 4572 234 4590 252
rect 4572 252 4590 270
rect 4572 270 4590 288
rect 4572 288 4590 306
rect 4572 306 4590 324
rect 4572 324 4590 342
rect 4572 342 4590 360
rect 4572 360 4590 378
rect 4572 378 4590 396
rect 4572 396 4590 414
rect 4572 414 4590 432
rect 4572 432 4590 450
rect 4572 450 4590 468
rect 4572 468 4590 486
rect 4572 486 4590 504
rect 4572 504 4590 522
rect 4572 522 4590 540
rect 4572 540 4590 558
rect 4572 558 4590 576
rect 4572 576 4590 594
rect 4572 594 4590 612
rect 4572 612 4590 630
rect 4572 630 4590 648
rect 4572 648 4590 666
rect 4572 666 4590 684
rect 4572 684 4590 702
rect 4572 702 4590 720
rect 4572 720 4590 738
rect 4572 738 4590 756
rect 4572 864 4590 882
rect 4572 882 4590 900
rect 4572 900 4590 918
rect 4572 918 4590 936
rect 4572 936 4590 954
rect 4572 954 4590 972
rect 4572 972 4590 990
rect 4572 990 4590 1008
rect 4572 1008 4590 1026
rect 4572 1026 4590 1044
rect 4572 1044 4590 1062
rect 4572 1062 4590 1080
rect 4572 1080 4590 1098
rect 4572 1098 4590 1116
rect 4572 1116 4590 1134
rect 4572 1134 4590 1152
rect 4572 1152 4590 1170
rect 4572 1170 4590 1188
rect 4572 1188 4590 1206
rect 4572 1206 4590 1224
rect 4572 1224 4590 1242
rect 4572 1242 4590 1260
rect 4572 1260 4590 1278
rect 4572 1278 4590 1296
rect 4572 1296 4590 1314
rect 4572 1314 4590 1332
rect 4572 1332 4590 1350
rect 4572 1350 4590 1368
rect 4572 1368 4590 1386
rect 4572 1386 4590 1404
rect 4572 1404 4590 1422
rect 4572 1422 4590 1440
rect 4572 1440 4590 1458
rect 4572 1458 4590 1476
rect 4572 1476 4590 1494
rect 4572 1494 4590 1512
rect 4572 1512 4590 1530
rect 4572 1530 4590 1548
rect 4572 1548 4590 1566
rect 4572 1566 4590 1584
rect 4572 1584 4590 1602
rect 4572 1602 4590 1620
rect 4572 1620 4590 1638
rect 4572 1638 4590 1656
rect 4572 1656 4590 1674
rect 4572 1674 4590 1692
rect 4572 1692 4590 1710
rect 4572 1710 4590 1728
rect 4572 1728 4590 1746
rect 4572 1746 4590 1764
rect 4572 1764 4590 1782
rect 4572 1782 4590 1800
rect 4572 1800 4590 1818
rect 4572 1818 4590 1836
rect 4572 1836 4590 1854
rect 4572 1854 4590 1872
rect 4572 1872 4590 1890
rect 4572 1890 4590 1908
rect 4572 1908 4590 1926
rect 4572 1926 4590 1944
rect 4572 2178 4590 2196
rect 4572 2196 4590 2214
rect 4572 2214 4590 2232
rect 4572 2232 4590 2250
rect 4572 2250 4590 2268
rect 4572 2268 4590 2286
rect 4572 2286 4590 2304
rect 4572 2304 4590 2322
rect 4572 2322 4590 2340
rect 4572 2340 4590 2358
rect 4572 2358 4590 2376
rect 4572 2376 4590 2394
rect 4572 2394 4590 2412
rect 4572 2412 4590 2430
rect 4572 2430 4590 2448
rect 4572 2448 4590 2466
rect 4572 2466 4590 2484
rect 4572 2484 4590 2502
rect 4572 2502 4590 2520
rect 4572 2520 4590 2538
rect 4572 2538 4590 2556
rect 4572 2556 4590 2574
rect 4572 2574 4590 2592
rect 4572 2592 4590 2610
rect 4572 2610 4590 2628
rect 4572 2628 4590 2646
rect 4572 2646 4590 2664
rect 4572 2664 4590 2682
rect 4572 2682 4590 2700
rect 4572 2700 4590 2718
rect 4572 2718 4590 2736
rect 4572 2736 4590 2754
rect 4572 2754 4590 2772
rect 4572 2772 4590 2790
rect 4572 2790 4590 2808
rect 4572 2808 4590 2826
rect 4572 2826 4590 2844
rect 4572 2844 4590 2862
rect 4572 2862 4590 2880
rect 4572 2880 4590 2898
rect 4572 2898 4590 2916
rect 4572 2916 4590 2934
rect 4572 2934 4590 2952
rect 4572 2952 4590 2970
rect 4572 2970 4590 2988
rect 4572 2988 4590 3006
rect 4572 3006 4590 3024
rect 4572 3024 4590 3042
rect 4572 3042 4590 3060
rect 4572 3060 4590 3078
rect 4572 3078 4590 3096
rect 4572 3096 4590 3114
rect 4572 3114 4590 3132
rect 4572 3132 4590 3150
rect 4572 3150 4590 3168
rect 4572 3168 4590 3186
rect 4572 3186 4590 3204
rect 4572 3204 4590 3222
rect 4572 3222 4590 3240
rect 4572 3240 4590 3258
rect 4572 3258 4590 3276
rect 4572 3276 4590 3294
rect 4572 3294 4590 3312
rect 4572 3312 4590 3330
rect 4572 3330 4590 3348
rect 4572 3348 4590 3366
rect 4572 3366 4590 3384
rect 4572 3384 4590 3402
rect 4572 3402 4590 3420
rect 4572 3420 4590 3438
rect 4572 3438 4590 3456
rect 4572 3456 4590 3474
rect 4572 3474 4590 3492
rect 4572 3492 4590 3510
rect 4572 3510 4590 3528
rect 4572 3528 4590 3546
rect 4572 3546 4590 3564
rect 4572 3564 4590 3582
rect 4572 3582 4590 3600
rect 4572 3600 4590 3618
rect 4572 3618 4590 3636
rect 4572 3636 4590 3654
rect 4572 3654 4590 3672
rect 4572 3672 4590 3690
rect 4572 3690 4590 3708
rect 4572 3708 4590 3726
rect 4572 3726 4590 3744
rect 4572 3744 4590 3762
rect 4572 3762 4590 3780
rect 4572 3780 4590 3798
rect 4572 3798 4590 3816
rect 4572 3816 4590 3834
rect 4572 3834 4590 3852
rect 4572 3852 4590 3870
rect 4572 3870 4590 3888
rect 4572 4086 4590 4104
rect 4572 4104 4590 4122
rect 4572 4122 4590 4140
rect 4572 4140 4590 4158
rect 4572 4158 4590 4176
rect 4572 4176 4590 4194
rect 4572 4194 4590 4212
rect 4572 4212 4590 4230
rect 4572 4230 4590 4248
rect 4572 4248 4590 4266
rect 4572 4266 4590 4284
rect 4572 4284 4590 4302
rect 4572 4302 4590 4320
rect 4572 4320 4590 4338
rect 4572 4338 4590 4356
rect 4572 4356 4590 4374
rect 4572 4374 4590 4392
rect 4572 4392 4590 4410
rect 4572 4410 4590 4428
rect 4572 4428 4590 4446
rect 4572 4446 4590 4464
rect 4572 4464 4590 4482
rect 4572 4482 4590 4500
rect 4572 4500 4590 4518
rect 4572 4518 4590 4536
rect 4572 4536 4590 4554
rect 4572 4554 4590 4572
rect 4572 4572 4590 4590
rect 4572 4590 4590 4608
rect 4572 4608 4590 4626
rect 4572 4626 4590 4644
rect 4572 4644 4590 4662
rect 4572 4662 4590 4680
rect 4572 4680 4590 4698
rect 4572 4698 4590 4716
rect 4572 4716 4590 4734
rect 4572 4734 4590 4752
rect 4572 4752 4590 4770
rect 4572 4770 4590 4788
rect 4572 4788 4590 4806
rect 4572 4806 4590 4824
rect 4572 4824 4590 4842
rect 4572 4842 4590 4860
rect 4572 4860 4590 4878
rect 4572 4878 4590 4896
rect 4572 4896 4590 4914
rect 4572 4914 4590 4932
rect 4572 4932 4590 4950
rect 4572 4950 4590 4968
rect 4572 4968 4590 4986
rect 4572 4986 4590 5004
rect 4572 5004 4590 5022
rect 4572 5022 4590 5040
rect 4572 5040 4590 5058
rect 4572 5058 4590 5076
rect 4572 5076 4590 5094
rect 4572 5094 4590 5112
rect 4572 5112 4590 5130
rect 4572 5130 4590 5148
rect 4572 5148 4590 5166
rect 4572 5166 4590 5184
rect 4572 5184 4590 5202
rect 4572 5202 4590 5220
rect 4572 5220 4590 5238
rect 4572 5238 4590 5256
rect 4572 5256 4590 5274
rect 4572 5274 4590 5292
rect 4572 5292 4590 5310
rect 4572 5310 4590 5328
rect 4572 5328 4590 5346
rect 4572 5346 4590 5364
rect 4572 5364 4590 5382
rect 4572 5382 4590 5400
rect 4572 5400 4590 5418
rect 4572 5418 4590 5436
rect 4572 5436 4590 5454
rect 4572 5454 4590 5472
rect 4572 5472 4590 5490
rect 4572 5490 4590 5508
rect 4572 5508 4590 5526
rect 4572 5526 4590 5544
rect 4572 5544 4590 5562
rect 4572 5562 4590 5580
rect 4572 5580 4590 5598
rect 4572 5598 4590 5616
rect 4572 5616 4590 5634
rect 4572 5634 4590 5652
rect 4572 5652 4590 5670
rect 4572 5670 4590 5688
rect 4572 5688 4590 5706
rect 4572 5706 4590 5724
rect 4572 5724 4590 5742
rect 4572 5742 4590 5760
rect 4572 5760 4590 5778
rect 4572 5778 4590 5796
rect 4572 5796 4590 5814
rect 4572 5814 4590 5832
rect 4572 5832 4590 5850
rect 4572 5850 4590 5868
rect 4572 5868 4590 5886
rect 4572 5886 4590 5904
rect 4572 5904 4590 5922
rect 4572 5922 4590 5940
rect 4572 5940 4590 5958
rect 4572 5958 4590 5976
rect 4572 5976 4590 5994
rect 4572 5994 4590 6012
rect 4572 6012 4590 6030
rect 4572 6030 4590 6048
rect 4572 6048 4590 6066
rect 4572 6066 4590 6084
rect 4572 6084 4590 6102
rect 4572 6102 4590 6120
rect 4572 6120 4590 6138
rect 4572 6138 4590 6156
rect 4572 6156 4590 6174
rect 4572 6174 4590 6192
rect 4572 6192 4590 6210
rect 4572 6210 4590 6228
rect 4572 6228 4590 6246
rect 4572 6246 4590 6264
rect 4572 6264 4590 6282
rect 4572 6282 4590 6300
rect 4572 6300 4590 6318
rect 4572 6318 4590 6336
rect 4572 6336 4590 6354
rect 4572 6354 4590 6372
rect 4572 6372 4590 6390
rect 4572 6390 4590 6408
rect 4572 6408 4590 6426
rect 4572 6426 4590 6444
rect 4572 6444 4590 6462
rect 4572 6462 4590 6480
rect 4572 6480 4590 6498
rect 4572 6498 4590 6516
rect 4572 6516 4590 6534
rect 4572 6534 4590 6552
rect 4572 6552 4590 6570
rect 4572 6570 4590 6588
rect 4572 6588 4590 6606
rect 4572 6606 4590 6624
rect 4572 6624 4590 6642
rect 4572 6642 4590 6660
rect 4572 6660 4590 6678
rect 4572 6678 4590 6696
rect 4572 6696 4590 6714
rect 4572 6714 4590 6732
rect 4572 6732 4590 6750
rect 4572 6750 4590 6768
rect 4572 6768 4590 6786
rect 4572 6786 4590 6804
rect 4572 6804 4590 6822
rect 4572 6822 4590 6840
rect 4572 6840 4590 6858
rect 4572 6858 4590 6876
rect 4572 6876 4590 6894
rect 4572 6894 4590 6912
rect 4572 6912 4590 6930
rect 4572 6930 4590 6948
rect 4572 6948 4590 6966
rect 4572 6966 4590 6984
rect 4572 6984 4590 7002
rect 4572 7002 4590 7020
rect 4572 7020 4590 7038
rect 4572 7038 4590 7056
rect 4572 7056 4590 7074
rect 4572 7074 4590 7092
rect 4572 7092 4590 7110
rect 4572 7110 4590 7128
rect 4572 7128 4590 7146
rect 4572 7146 4590 7164
rect 4590 126 4608 144
rect 4590 144 4608 162
rect 4590 162 4608 180
rect 4590 180 4608 198
rect 4590 198 4608 216
rect 4590 216 4608 234
rect 4590 234 4608 252
rect 4590 252 4608 270
rect 4590 270 4608 288
rect 4590 288 4608 306
rect 4590 306 4608 324
rect 4590 324 4608 342
rect 4590 342 4608 360
rect 4590 360 4608 378
rect 4590 378 4608 396
rect 4590 396 4608 414
rect 4590 414 4608 432
rect 4590 432 4608 450
rect 4590 450 4608 468
rect 4590 468 4608 486
rect 4590 486 4608 504
rect 4590 504 4608 522
rect 4590 522 4608 540
rect 4590 540 4608 558
rect 4590 558 4608 576
rect 4590 576 4608 594
rect 4590 594 4608 612
rect 4590 612 4608 630
rect 4590 630 4608 648
rect 4590 648 4608 666
rect 4590 666 4608 684
rect 4590 684 4608 702
rect 4590 702 4608 720
rect 4590 720 4608 738
rect 4590 738 4608 756
rect 4590 864 4608 882
rect 4590 882 4608 900
rect 4590 900 4608 918
rect 4590 918 4608 936
rect 4590 936 4608 954
rect 4590 954 4608 972
rect 4590 972 4608 990
rect 4590 990 4608 1008
rect 4590 1008 4608 1026
rect 4590 1026 4608 1044
rect 4590 1044 4608 1062
rect 4590 1062 4608 1080
rect 4590 1080 4608 1098
rect 4590 1098 4608 1116
rect 4590 1116 4608 1134
rect 4590 1134 4608 1152
rect 4590 1152 4608 1170
rect 4590 1170 4608 1188
rect 4590 1188 4608 1206
rect 4590 1206 4608 1224
rect 4590 1224 4608 1242
rect 4590 1242 4608 1260
rect 4590 1260 4608 1278
rect 4590 1278 4608 1296
rect 4590 1296 4608 1314
rect 4590 1314 4608 1332
rect 4590 1332 4608 1350
rect 4590 1350 4608 1368
rect 4590 1368 4608 1386
rect 4590 1386 4608 1404
rect 4590 1404 4608 1422
rect 4590 1422 4608 1440
rect 4590 1440 4608 1458
rect 4590 1458 4608 1476
rect 4590 1476 4608 1494
rect 4590 1494 4608 1512
rect 4590 1512 4608 1530
rect 4590 1530 4608 1548
rect 4590 1548 4608 1566
rect 4590 1566 4608 1584
rect 4590 1584 4608 1602
rect 4590 1602 4608 1620
rect 4590 1620 4608 1638
rect 4590 1638 4608 1656
rect 4590 1656 4608 1674
rect 4590 1674 4608 1692
rect 4590 1692 4608 1710
rect 4590 1710 4608 1728
rect 4590 1728 4608 1746
rect 4590 1746 4608 1764
rect 4590 1764 4608 1782
rect 4590 1782 4608 1800
rect 4590 1800 4608 1818
rect 4590 1818 4608 1836
rect 4590 1836 4608 1854
rect 4590 1854 4608 1872
rect 4590 1872 4608 1890
rect 4590 1890 4608 1908
rect 4590 1908 4608 1926
rect 4590 1926 4608 1944
rect 4590 1944 4608 1962
rect 4590 2196 4608 2214
rect 4590 2214 4608 2232
rect 4590 2232 4608 2250
rect 4590 2250 4608 2268
rect 4590 2268 4608 2286
rect 4590 2286 4608 2304
rect 4590 2304 4608 2322
rect 4590 2322 4608 2340
rect 4590 2340 4608 2358
rect 4590 2358 4608 2376
rect 4590 2376 4608 2394
rect 4590 2394 4608 2412
rect 4590 2412 4608 2430
rect 4590 2430 4608 2448
rect 4590 2448 4608 2466
rect 4590 2466 4608 2484
rect 4590 2484 4608 2502
rect 4590 2502 4608 2520
rect 4590 2520 4608 2538
rect 4590 2538 4608 2556
rect 4590 2556 4608 2574
rect 4590 2574 4608 2592
rect 4590 2592 4608 2610
rect 4590 2610 4608 2628
rect 4590 2628 4608 2646
rect 4590 2646 4608 2664
rect 4590 2664 4608 2682
rect 4590 2682 4608 2700
rect 4590 2700 4608 2718
rect 4590 2718 4608 2736
rect 4590 2736 4608 2754
rect 4590 2754 4608 2772
rect 4590 2772 4608 2790
rect 4590 2790 4608 2808
rect 4590 2808 4608 2826
rect 4590 2826 4608 2844
rect 4590 2844 4608 2862
rect 4590 2862 4608 2880
rect 4590 2880 4608 2898
rect 4590 2898 4608 2916
rect 4590 2916 4608 2934
rect 4590 2934 4608 2952
rect 4590 2952 4608 2970
rect 4590 2970 4608 2988
rect 4590 2988 4608 3006
rect 4590 3006 4608 3024
rect 4590 3024 4608 3042
rect 4590 3042 4608 3060
rect 4590 3060 4608 3078
rect 4590 3078 4608 3096
rect 4590 3096 4608 3114
rect 4590 3114 4608 3132
rect 4590 3132 4608 3150
rect 4590 3150 4608 3168
rect 4590 3168 4608 3186
rect 4590 3186 4608 3204
rect 4590 3204 4608 3222
rect 4590 3222 4608 3240
rect 4590 3240 4608 3258
rect 4590 3258 4608 3276
rect 4590 3276 4608 3294
rect 4590 3294 4608 3312
rect 4590 3312 4608 3330
rect 4590 3330 4608 3348
rect 4590 3348 4608 3366
rect 4590 3366 4608 3384
rect 4590 3384 4608 3402
rect 4590 3402 4608 3420
rect 4590 3420 4608 3438
rect 4590 3438 4608 3456
rect 4590 3456 4608 3474
rect 4590 3474 4608 3492
rect 4590 3492 4608 3510
rect 4590 3510 4608 3528
rect 4590 3528 4608 3546
rect 4590 3546 4608 3564
rect 4590 3564 4608 3582
rect 4590 3582 4608 3600
rect 4590 3600 4608 3618
rect 4590 3618 4608 3636
rect 4590 3636 4608 3654
rect 4590 3654 4608 3672
rect 4590 3672 4608 3690
rect 4590 3690 4608 3708
rect 4590 3708 4608 3726
rect 4590 3726 4608 3744
rect 4590 3744 4608 3762
rect 4590 3762 4608 3780
rect 4590 3780 4608 3798
rect 4590 3798 4608 3816
rect 4590 3816 4608 3834
rect 4590 3834 4608 3852
rect 4590 3852 4608 3870
rect 4590 3870 4608 3888
rect 4590 3888 4608 3906
rect 4590 4104 4608 4122
rect 4590 4122 4608 4140
rect 4590 4140 4608 4158
rect 4590 4158 4608 4176
rect 4590 4176 4608 4194
rect 4590 4194 4608 4212
rect 4590 4212 4608 4230
rect 4590 4230 4608 4248
rect 4590 4248 4608 4266
rect 4590 4266 4608 4284
rect 4590 4284 4608 4302
rect 4590 4302 4608 4320
rect 4590 4320 4608 4338
rect 4590 4338 4608 4356
rect 4590 4356 4608 4374
rect 4590 4374 4608 4392
rect 4590 4392 4608 4410
rect 4590 4410 4608 4428
rect 4590 4428 4608 4446
rect 4590 4446 4608 4464
rect 4590 4464 4608 4482
rect 4590 4482 4608 4500
rect 4590 4500 4608 4518
rect 4590 4518 4608 4536
rect 4590 4536 4608 4554
rect 4590 4554 4608 4572
rect 4590 4572 4608 4590
rect 4590 4590 4608 4608
rect 4590 4608 4608 4626
rect 4590 4626 4608 4644
rect 4590 4644 4608 4662
rect 4590 4662 4608 4680
rect 4590 4680 4608 4698
rect 4590 4698 4608 4716
rect 4590 4716 4608 4734
rect 4590 4734 4608 4752
rect 4590 4752 4608 4770
rect 4590 4770 4608 4788
rect 4590 4788 4608 4806
rect 4590 4806 4608 4824
rect 4590 4824 4608 4842
rect 4590 4842 4608 4860
rect 4590 4860 4608 4878
rect 4590 4878 4608 4896
rect 4590 4896 4608 4914
rect 4590 4914 4608 4932
rect 4590 4932 4608 4950
rect 4590 4950 4608 4968
rect 4590 4968 4608 4986
rect 4590 4986 4608 5004
rect 4590 5004 4608 5022
rect 4590 5022 4608 5040
rect 4590 5040 4608 5058
rect 4590 5058 4608 5076
rect 4590 5076 4608 5094
rect 4590 5094 4608 5112
rect 4590 5112 4608 5130
rect 4590 5130 4608 5148
rect 4590 5148 4608 5166
rect 4590 5166 4608 5184
rect 4590 5184 4608 5202
rect 4590 5202 4608 5220
rect 4590 5220 4608 5238
rect 4590 5238 4608 5256
rect 4590 5256 4608 5274
rect 4590 5274 4608 5292
rect 4590 5292 4608 5310
rect 4590 5310 4608 5328
rect 4590 5328 4608 5346
rect 4590 5346 4608 5364
rect 4590 5364 4608 5382
rect 4590 5382 4608 5400
rect 4590 5400 4608 5418
rect 4590 5418 4608 5436
rect 4590 5436 4608 5454
rect 4590 5454 4608 5472
rect 4590 5472 4608 5490
rect 4590 5490 4608 5508
rect 4590 5508 4608 5526
rect 4590 5526 4608 5544
rect 4590 5544 4608 5562
rect 4590 5562 4608 5580
rect 4590 5580 4608 5598
rect 4590 5598 4608 5616
rect 4590 5616 4608 5634
rect 4590 5634 4608 5652
rect 4590 5652 4608 5670
rect 4590 5670 4608 5688
rect 4590 5688 4608 5706
rect 4590 5706 4608 5724
rect 4590 5724 4608 5742
rect 4590 5742 4608 5760
rect 4590 5760 4608 5778
rect 4590 5778 4608 5796
rect 4590 5796 4608 5814
rect 4590 5814 4608 5832
rect 4590 5832 4608 5850
rect 4590 5850 4608 5868
rect 4590 5868 4608 5886
rect 4590 5886 4608 5904
rect 4590 5904 4608 5922
rect 4590 5922 4608 5940
rect 4590 5940 4608 5958
rect 4590 5958 4608 5976
rect 4590 5976 4608 5994
rect 4590 5994 4608 6012
rect 4590 6012 4608 6030
rect 4590 6030 4608 6048
rect 4590 6048 4608 6066
rect 4590 6066 4608 6084
rect 4590 6084 4608 6102
rect 4590 6102 4608 6120
rect 4590 6120 4608 6138
rect 4590 6138 4608 6156
rect 4590 6156 4608 6174
rect 4590 6174 4608 6192
rect 4590 6192 4608 6210
rect 4590 6210 4608 6228
rect 4590 6228 4608 6246
rect 4590 6246 4608 6264
rect 4590 6264 4608 6282
rect 4590 6282 4608 6300
rect 4590 6300 4608 6318
rect 4590 6318 4608 6336
rect 4590 6336 4608 6354
rect 4590 6354 4608 6372
rect 4590 6372 4608 6390
rect 4590 6390 4608 6408
rect 4590 6408 4608 6426
rect 4590 6426 4608 6444
rect 4590 6444 4608 6462
rect 4590 6462 4608 6480
rect 4590 6480 4608 6498
rect 4590 6498 4608 6516
rect 4590 6516 4608 6534
rect 4590 6534 4608 6552
rect 4590 6552 4608 6570
rect 4590 6570 4608 6588
rect 4590 6588 4608 6606
rect 4590 6606 4608 6624
rect 4590 6624 4608 6642
rect 4590 6642 4608 6660
rect 4590 6660 4608 6678
rect 4590 6678 4608 6696
rect 4590 6696 4608 6714
rect 4590 6714 4608 6732
rect 4590 6732 4608 6750
rect 4590 6750 4608 6768
rect 4590 6768 4608 6786
rect 4590 6786 4608 6804
rect 4590 6804 4608 6822
rect 4590 6822 4608 6840
rect 4590 6840 4608 6858
rect 4590 6858 4608 6876
rect 4590 6876 4608 6894
rect 4590 6894 4608 6912
rect 4590 6912 4608 6930
rect 4590 6930 4608 6948
rect 4590 6948 4608 6966
rect 4590 6966 4608 6984
rect 4590 6984 4608 7002
rect 4590 7002 4608 7020
rect 4590 7020 4608 7038
rect 4590 7038 4608 7056
rect 4590 7056 4608 7074
rect 4590 7074 4608 7092
rect 4590 7092 4608 7110
rect 4590 7110 4608 7128
rect 4590 7128 4608 7146
rect 4590 7146 4608 7164
rect 4590 7164 4608 7182
rect 4590 7182 4608 7200
rect 4608 126 4626 144
rect 4608 144 4626 162
rect 4608 162 4626 180
rect 4608 180 4626 198
rect 4608 198 4626 216
rect 4608 216 4626 234
rect 4608 234 4626 252
rect 4608 252 4626 270
rect 4608 270 4626 288
rect 4608 288 4626 306
rect 4608 306 4626 324
rect 4608 324 4626 342
rect 4608 342 4626 360
rect 4608 360 4626 378
rect 4608 378 4626 396
rect 4608 396 4626 414
rect 4608 414 4626 432
rect 4608 432 4626 450
rect 4608 450 4626 468
rect 4608 468 4626 486
rect 4608 486 4626 504
rect 4608 504 4626 522
rect 4608 522 4626 540
rect 4608 540 4626 558
rect 4608 558 4626 576
rect 4608 576 4626 594
rect 4608 594 4626 612
rect 4608 612 4626 630
rect 4608 630 4626 648
rect 4608 648 4626 666
rect 4608 666 4626 684
rect 4608 684 4626 702
rect 4608 702 4626 720
rect 4608 720 4626 738
rect 4608 738 4626 756
rect 4608 864 4626 882
rect 4608 882 4626 900
rect 4608 900 4626 918
rect 4608 918 4626 936
rect 4608 936 4626 954
rect 4608 954 4626 972
rect 4608 972 4626 990
rect 4608 990 4626 1008
rect 4608 1008 4626 1026
rect 4608 1026 4626 1044
rect 4608 1044 4626 1062
rect 4608 1062 4626 1080
rect 4608 1080 4626 1098
rect 4608 1098 4626 1116
rect 4608 1116 4626 1134
rect 4608 1134 4626 1152
rect 4608 1152 4626 1170
rect 4608 1170 4626 1188
rect 4608 1188 4626 1206
rect 4608 1206 4626 1224
rect 4608 1224 4626 1242
rect 4608 1242 4626 1260
rect 4608 1260 4626 1278
rect 4608 1278 4626 1296
rect 4608 1296 4626 1314
rect 4608 1314 4626 1332
rect 4608 1332 4626 1350
rect 4608 1350 4626 1368
rect 4608 1368 4626 1386
rect 4608 1386 4626 1404
rect 4608 1404 4626 1422
rect 4608 1422 4626 1440
rect 4608 1440 4626 1458
rect 4608 1458 4626 1476
rect 4608 1476 4626 1494
rect 4608 1494 4626 1512
rect 4608 1512 4626 1530
rect 4608 1530 4626 1548
rect 4608 1548 4626 1566
rect 4608 1566 4626 1584
rect 4608 1584 4626 1602
rect 4608 1602 4626 1620
rect 4608 1620 4626 1638
rect 4608 1638 4626 1656
rect 4608 1656 4626 1674
rect 4608 1674 4626 1692
rect 4608 1692 4626 1710
rect 4608 1710 4626 1728
rect 4608 1728 4626 1746
rect 4608 1746 4626 1764
rect 4608 1764 4626 1782
rect 4608 1782 4626 1800
rect 4608 1800 4626 1818
rect 4608 1818 4626 1836
rect 4608 1836 4626 1854
rect 4608 1854 4626 1872
rect 4608 1872 4626 1890
rect 4608 1890 4626 1908
rect 4608 1908 4626 1926
rect 4608 1926 4626 1944
rect 4608 1944 4626 1962
rect 4608 1962 4626 1980
rect 4608 2214 4626 2232
rect 4608 2232 4626 2250
rect 4608 2250 4626 2268
rect 4608 2268 4626 2286
rect 4608 2286 4626 2304
rect 4608 2304 4626 2322
rect 4608 2322 4626 2340
rect 4608 2340 4626 2358
rect 4608 2358 4626 2376
rect 4608 2376 4626 2394
rect 4608 2394 4626 2412
rect 4608 2412 4626 2430
rect 4608 2430 4626 2448
rect 4608 2448 4626 2466
rect 4608 2466 4626 2484
rect 4608 2484 4626 2502
rect 4608 2502 4626 2520
rect 4608 2520 4626 2538
rect 4608 2538 4626 2556
rect 4608 2556 4626 2574
rect 4608 2574 4626 2592
rect 4608 2592 4626 2610
rect 4608 2610 4626 2628
rect 4608 2628 4626 2646
rect 4608 2646 4626 2664
rect 4608 2664 4626 2682
rect 4608 2682 4626 2700
rect 4608 2700 4626 2718
rect 4608 2718 4626 2736
rect 4608 2736 4626 2754
rect 4608 2754 4626 2772
rect 4608 2772 4626 2790
rect 4608 2790 4626 2808
rect 4608 2808 4626 2826
rect 4608 2826 4626 2844
rect 4608 2844 4626 2862
rect 4608 2862 4626 2880
rect 4608 2880 4626 2898
rect 4608 2898 4626 2916
rect 4608 2916 4626 2934
rect 4608 2934 4626 2952
rect 4608 2952 4626 2970
rect 4608 2970 4626 2988
rect 4608 2988 4626 3006
rect 4608 3006 4626 3024
rect 4608 3024 4626 3042
rect 4608 3042 4626 3060
rect 4608 3060 4626 3078
rect 4608 3078 4626 3096
rect 4608 3096 4626 3114
rect 4608 3114 4626 3132
rect 4608 3132 4626 3150
rect 4608 3150 4626 3168
rect 4608 3168 4626 3186
rect 4608 3186 4626 3204
rect 4608 3204 4626 3222
rect 4608 3222 4626 3240
rect 4608 3240 4626 3258
rect 4608 3258 4626 3276
rect 4608 3276 4626 3294
rect 4608 3294 4626 3312
rect 4608 3312 4626 3330
rect 4608 3330 4626 3348
rect 4608 3348 4626 3366
rect 4608 3366 4626 3384
rect 4608 3384 4626 3402
rect 4608 3402 4626 3420
rect 4608 3420 4626 3438
rect 4608 3438 4626 3456
rect 4608 3456 4626 3474
rect 4608 3474 4626 3492
rect 4608 3492 4626 3510
rect 4608 3510 4626 3528
rect 4608 3528 4626 3546
rect 4608 3546 4626 3564
rect 4608 3564 4626 3582
rect 4608 3582 4626 3600
rect 4608 3600 4626 3618
rect 4608 3618 4626 3636
rect 4608 3636 4626 3654
rect 4608 3654 4626 3672
rect 4608 3672 4626 3690
rect 4608 3690 4626 3708
rect 4608 3708 4626 3726
rect 4608 3726 4626 3744
rect 4608 3744 4626 3762
rect 4608 3762 4626 3780
rect 4608 3780 4626 3798
rect 4608 3798 4626 3816
rect 4608 3816 4626 3834
rect 4608 3834 4626 3852
rect 4608 3852 4626 3870
rect 4608 3870 4626 3888
rect 4608 3888 4626 3906
rect 4608 3906 4626 3924
rect 4608 4140 4626 4158
rect 4608 4158 4626 4176
rect 4608 4176 4626 4194
rect 4608 4194 4626 4212
rect 4608 4212 4626 4230
rect 4608 4230 4626 4248
rect 4608 4248 4626 4266
rect 4608 4266 4626 4284
rect 4608 4284 4626 4302
rect 4608 4302 4626 4320
rect 4608 4320 4626 4338
rect 4608 4338 4626 4356
rect 4608 4356 4626 4374
rect 4608 4374 4626 4392
rect 4608 4392 4626 4410
rect 4608 4410 4626 4428
rect 4608 4428 4626 4446
rect 4608 4446 4626 4464
rect 4608 4464 4626 4482
rect 4608 4482 4626 4500
rect 4608 4500 4626 4518
rect 4608 4518 4626 4536
rect 4608 4536 4626 4554
rect 4608 4554 4626 4572
rect 4608 4572 4626 4590
rect 4608 4590 4626 4608
rect 4608 4608 4626 4626
rect 4608 4626 4626 4644
rect 4608 4644 4626 4662
rect 4608 4662 4626 4680
rect 4608 4680 4626 4698
rect 4608 4698 4626 4716
rect 4608 4716 4626 4734
rect 4608 4734 4626 4752
rect 4608 4752 4626 4770
rect 4608 4770 4626 4788
rect 4608 4788 4626 4806
rect 4608 4806 4626 4824
rect 4608 4824 4626 4842
rect 4608 4842 4626 4860
rect 4608 4860 4626 4878
rect 4608 4878 4626 4896
rect 4608 4896 4626 4914
rect 4608 4914 4626 4932
rect 4608 4932 4626 4950
rect 4608 4950 4626 4968
rect 4608 4968 4626 4986
rect 4608 4986 4626 5004
rect 4608 5004 4626 5022
rect 4608 5022 4626 5040
rect 4608 5040 4626 5058
rect 4608 5058 4626 5076
rect 4608 5076 4626 5094
rect 4608 5094 4626 5112
rect 4608 5112 4626 5130
rect 4608 5130 4626 5148
rect 4608 5148 4626 5166
rect 4608 5166 4626 5184
rect 4608 5184 4626 5202
rect 4608 5202 4626 5220
rect 4608 5220 4626 5238
rect 4608 5238 4626 5256
rect 4608 5256 4626 5274
rect 4608 5274 4626 5292
rect 4608 5292 4626 5310
rect 4608 5310 4626 5328
rect 4608 5328 4626 5346
rect 4608 5346 4626 5364
rect 4608 5364 4626 5382
rect 4608 5382 4626 5400
rect 4608 5400 4626 5418
rect 4608 5418 4626 5436
rect 4608 5436 4626 5454
rect 4608 5454 4626 5472
rect 4608 5472 4626 5490
rect 4608 5490 4626 5508
rect 4608 5508 4626 5526
rect 4608 5526 4626 5544
rect 4608 5544 4626 5562
rect 4608 5562 4626 5580
rect 4608 5580 4626 5598
rect 4608 5598 4626 5616
rect 4608 5616 4626 5634
rect 4608 5634 4626 5652
rect 4608 5652 4626 5670
rect 4608 5670 4626 5688
rect 4608 5688 4626 5706
rect 4608 5706 4626 5724
rect 4608 5724 4626 5742
rect 4608 5742 4626 5760
rect 4608 5760 4626 5778
rect 4608 5778 4626 5796
rect 4608 5796 4626 5814
rect 4608 5814 4626 5832
rect 4608 5832 4626 5850
rect 4608 5850 4626 5868
rect 4608 5868 4626 5886
rect 4608 5886 4626 5904
rect 4608 5904 4626 5922
rect 4608 5922 4626 5940
rect 4608 5940 4626 5958
rect 4608 5958 4626 5976
rect 4608 5976 4626 5994
rect 4608 5994 4626 6012
rect 4608 6012 4626 6030
rect 4608 6030 4626 6048
rect 4608 6048 4626 6066
rect 4608 6066 4626 6084
rect 4608 6084 4626 6102
rect 4608 6102 4626 6120
rect 4608 6120 4626 6138
rect 4608 6138 4626 6156
rect 4608 6156 4626 6174
rect 4608 6174 4626 6192
rect 4608 6192 4626 6210
rect 4608 6210 4626 6228
rect 4608 6228 4626 6246
rect 4608 6246 4626 6264
rect 4608 6264 4626 6282
rect 4608 6282 4626 6300
rect 4608 6300 4626 6318
rect 4608 6318 4626 6336
rect 4608 6336 4626 6354
rect 4608 6354 4626 6372
rect 4608 6372 4626 6390
rect 4608 6390 4626 6408
rect 4608 6408 4626 6426
rect 4608 6426 4626 6444
rect 4608 6444 4626 6462
rect 4608 6462 4626 6480
rect 4608 6480 4626 6498
rect 4608 6498 4626 6516
rect 4608 6516 4626 6534
rect 4608 6534 4626 6552
rect 4608 6552 4626 6570
rect 4608 6570 4626 6588
rect 4608 6588 4626 6606
rect 4608 6606 4626 6624
rect 4608 6624 4626 6642
rect 4608 6642 4626 6660
rect 4608 6660 4626 6678
rect 4608 6678 4626 6696
rect 4608 6696 4626 6714
rect 4608 6714 4626 6732
rect 4608 6732 4626 6750
rect 4608 6750 4626 6768
rect 4608 6768 4626 6786
rect 4608 6786 4626 6804
rect 4608 6804 4626 6822
rect 4608 6822 4626 6840
rect 4608 6840 4626 6858
rect 4608 6858 4626 6876
rect 4608 6876 4626 6894
rect 4608 6894 4626 6912
rect 4608 6912 4626 6930
rect 4608 6930 4626 6948
rect 4608 6948 4626 6966
rect 4608 6966 4626 6984
rect 4608 6984 4626 7002
rect 4608 7002 4626 7020
rect 4608 7020 4626 7038
rect 4608 7038 4626 7056
rect 4608 7056 4626 7074
rect 4608 7074 4626 7092
rect 4608 7092 4626 7110
rect 4608 7110 4626 7128
rect 4608 7128 4626 7146
rect 4608 7146 4626 7164
rect 4608 7164 4626 7182
rect 4608 7182 4626 7200
rect 4608 7200 4626 7218
rect 4626 144 4644 162
rect 4626 162 4644 180
rect 4626 180 4644 198
rect 4626 198 4644 216
rect 4626 216 4644 234
rect 4626 234 4644 252
rect 4626 252 4644 270
rect 4626 270 4644 288
rect 4626 288 4644 306
rect 4626 306 4644 324
rect 4626 324 4644 342
rect 4626 342 4644 360
rect 4626 360 4644 378
rect 4626 378 4644 396
rect 4626 396 4644 414
rect 4626 414 4644 432
rect 4626 432 4644 450
rect 4626 450 4644 468
rect 4626 468 4644 486
rect 4626 486 4644 504
rect 4626 504 4644 522
rect 4626 522 4644 540
rect 4626 540 4644 558
rect 4626 558 4644 576
rect 4626 576 4644 594
rect 4626 594 4644 612
rect 4626 612 4644 630
rect 4626 630 4644 648
rect 4626 648 4644 666
rect 4626 666 4644 684
rect 4626 684 4644 702
rect 4626 702 4644 720
rect 4626 720 4644 738
rect 4626 738 4644 756
rect 4626 864 4644 882
rect 4626 882 4644 900
rect 4626 900 4644 918
rect 4626 918 4644 936
rect 4626 936 4644 954
rect 4626 954 4644 972
rect 4626 972 4644 990
rect 4626 990 4644 1008
rect 4626 1008 4644 1026
rect 4626 1026 4644 1044
rect 4626 1044 4644 1062
rect 4626 1062 4644 1080
rect 4626 1080 4644 1098
rect 4626 1098 4644 1116
rect 4626 1116 4644 1134
rect 4626 1134 4644 1152
rect 4626 1152 4644 1170
rect 4626 1170 4644 1188
rect 4626 1188 4644 1206
rect 4626 1206 4644 1224
rect 4626 1224 4644 1242
rect 4626 1242 4644 1260
rect 4626 1260 4644 1278
rect 4626 1278 4644 1296
rect 4626 1296 4644 1314
rect 4626 1314 4644 1332
rect 4626 1332 4644 1350
rect 4626 1350 4644 1368
rect 4626 1368 4644 1386
rect 4626 1386 4644 1404
rect 4626 1404 4644 1422
rect 4626 1422 4644 1440
rect 4626 1440 4644 1458
rect 4626 1458 4644 1476
rect 4626 1476 4644 1494
rect 4626 1494 4644 1512
rect 4626 1512 4644 1530
rect 4626 1530 4644 1548
rect 4626 1548 4644 1566
rect 4626 1566 4644 1584
rect 4626 1584 4644 1602
rect 4626 1602 4644 1620
rect 4626 1620 4644 1638
rect 4626 1638 4644 1656
rect 4626 1656 4644 1674
rect 4626 1674 4644 1692
rect 4626 1692 4644 1710
rect 4626 1710 4644 1728
rect 4626 1728 4644 1746
rect 4626 1746 4644 1764
rect 4626 1764 4644 1782
rect 4626 1782 4644 1800
rect 4626 1800 4644 1818
rect 4626 1818 4644 1836
rect 4626 1836 4644 1854
rect 4626 1854 4644 1872
rect 4626 1872 4644 1890
rect 4626 1890 4644 1908
rect 4626 1908 4644 1926
rect 4626 1926 4644 1944
rect 4626 1944 4644 1962
rect 4626 1962 4644 1980
rect 4626 2214 4644 2232
rect 4626 2232 4644 2250
rect 4626 2250 4644 2268
rect 4626 2268 4644 2286
rect 4626 2286 4644 2304
rect 4626 2304 4644 2322
rect 4626 2322 4644 2340
rect 4626 2340 4644 2358
rect 4626 2358 4644 2376
rect 4626 2376 4644 2394
rect 4626 2394 4644 2412
rect 4626 2412 4644 2430
rect 4626 2430 4644 2448
rect 4626 2448 4644 2466
rect 4626 2466 4644 2484
rect 4626 2484 4644 2502
rect 4626 2502 4644 2520
rect 4626 2520 4644 2538
rect 4626 2538 4644 2556
rect 4626 2556 4644 2574
rect 4626 2574 4644 2592
rect 4626 2592 4644 2610
rect 4626 2610 4644 2628
rect 4626 2628 4644 2646
rect 4626 2646 4644 2664
rect 4626 2664 4644 2682
rect 4626 2682 4644 2700
rect 4626 2700 4644 2718
rect 4626 2718 4644 2736
rect 4626 2736 4644 2754
rect 4626 2754 4644 2772
rect 4626 2772 4644 2790
rect 4626 2790 4644 2808
rect 4626 2808 4644 2826
rect 4626 2826 4644 2844
rect 4626 2844 4644 2862
rect 4626 2862 4644 2880
rect 4626 2880 4644 2898
rect 4626 2898 4644 2916
rect 4626 2916 4644 2934
rect 4626 2934 4644 2952
rect 4626 2952 4644 2970
rect 4626 2970 4644 2988
rect 4626 2988 4644 3006
rect 4626 3006 4644 3024
rect 4626 3024 4644 3042
rect 4626 3042 4644 3060
rect 4626 3060 4644 3078
rect 4626 3078 4644 3096
rect 4626 3096 4644 3114
rect 4626 3114 4644 3132
rect 4626 3132 4644 3150
rect 4626 3150 4644 3168
rect 4626 3168 4644 3186
rect 4626 3186 4644 3204
rect 4626 3204 4644 3222
rect 4626 3222 4644 3240
rect 4626 3240 4644 3258
rect 4626 3258 4644 3276
rect 4626 3276 4644 3294
rect 4626 3294 4644 3312
rect 4626 3312 4644 3330
rect 4626 3330 4644 3348
rect 4626 3348 4644 3366
rect 4626 3366 4644 3384
rect 4626 3384 4644 3402
rect 4626 3402 4644 3420
rect 4626 3420 4644 3438
rect 4626 3438 4644 3456
rect 4626 3456 4644 3474
rect 4626 3474 4644 3492
rect 4626 3492 4644 3510
rect 4626 3510 4644 3528
rect 4626 3528 4644 3546
rect 4626 3546 4644 3564
rect 4626 3564 4644 3582
rect 4626 3582 4644 3600
rect 4626 3600 4644 3618
rect 4626 3618 4644 3636
rect 4626 3636 4644 3654
rect 4626 3654 4644 3672
rect 4626 3672 4644 3690
rect 4626 3690 4644 3708
rect 4626 3708 4644 3726
rect 4626 3726 4644 3744
rect 4626 3744 4644 3762
rect 4626 3762 4644 3780
rect 4626 3780 4644 3798
rect 4626 3798 4644 3816
rect 4626 3816 4644 3834
rect 4626 3834 4644 3852
rect 4626 3852 4644 3870
rect 4626 3870 4644 3888
rect 4626 3888 4644 3906
rect 4626 3906 4644 3924
rect 4626 3924 4644 3942
rect 4626 3942 4644 3960
rect 4626 4158 4644 4176
rect 4626 4176 4644 4194
rect 4626 4194 4644 4212
rect 4626 4212 4644 4230
rect 4626 4230 4644 4248
rect 4626 4248 4644 4266
rect 4626 4266 4644 4284
rect 4626 4284 4644 4302
rect 4626 4302 4644 4320
rect 4626 4320 4644 4338
rect 4626 4338 4644 4356
rect 4626 4356 4644 4374
rect 4626 4374 4644 4392
rect 4626 4392 4644 4410
rect 4626 4410 4644 4428
rect 4626 4428 4644 4446
rect 4626 4446 4644 4464
rect 4626 4464 4644 4482
rect 4626 4482 4644 4500
rect 4626 4500 4644 4518
rect 4626 4518 4644 4536
rect 4626 4536 4644 4554
rect 4626 4554 4644 4572
rect 4626 4572 4644 4590
rect 4626 4590 4644 4608
rect 4626 4608 4644 4626
rect 4626 4626 4644 4644
rect 4626 4644 4644 4662
rect 4626 4662 4644 4680
rect 4626 4680 4644 4698
rect 4626 4698 4644 4716
rect 4626 4716 4644 4734
rect 4626 4734 4644 4752
rect 4626 4752 4644 4770
rect 4626 4770 4644 4788
rect 4626 4788 4644 4806
rect 4626 4806 4644 4824
rect 4626 4824 4644 4842
rect 4626 4842 4644 4860
rect 4626 4860 4644 4878
rect 4626 4878 4644 4896
rect 4626 4896 4644 4914
rect 4626 4914 4644 4932
rect 4626 4932 4644 4950
rect 4626 4950 4644 4968
rect 4626 4968 4644 4986
rect 4626 4986 4644 5004
rect 4626 5004 4644 5022
rect 4626 5022 4644 5040
rect 4626 5040 4644 5058
rect 4626 5058 4644 5076
rect 4626 5076 4644 5094
rect 4626 5094 4644 5112
rect 4626 5112 4644 5130
rect 4626 5130 4644 5148
rect 4626 5148 4644 5166
rect 4626 5166 4644 5184
rect 4626 5184 4644 5202
rect 4626 5202 4644 5220
rect 4626 5220 4644 5238
rect 4626 5238 4644 5256
rect 4626 5256 4644 5274
rect 4626 5274 4644 5292
rect 4626 5292 4644 5310
rect 4626 5310 4644 5328
rect 4626 5328 4644 5346
rect 4626 5346 4644 5364
rect 4626 5364 4644 5382
rect 4626 5382 4644 5400
rect 4626 5400 4644 5418
rect 4626 5418 4644 5436
rect 4626 5436 4644 5454
rect 4626 5454 4644 5472
rect 4626 5472 4644 5490
rect 4626 5490 4644 5508
rect 4626 5508 4644 5526
rect 4626 5526 4644 5544
rect 4626 5544 4644 5562
rect 4626 5562 4644 5580
rect 4626 5580 4644 5598
rect 4626 5598 4644 5616
rect 4626 5616 4644 5634
rect 4626 5634 4644 5652
rect 4626 5652 4644 5670
rect 4626 5670 4644 5688
rect 4626 5688 4644 5706
rect 4626 5706 4644 5724
rect 4626 5724 4644 5742
rect 4626 5742 4644 5760
rect 4626 5760 4644 5778
rect 4626 5778 4644 5796
rect 4626 5796 4644 5814
rect 4626 5814 4644 5832
rect 4626 5832 4644 5850
rect 4626 5850 4644 5868
rect 4626 5868 4644 5886
rect 4626 5886 4644 5904
rect 4626 5904 4644 5922
rect 4626 5922 4644 5940
rect 4626 5940 4644 5958
rect 4626 5958 4644 5976
rect 4626 5976 4644 5994
rect 4626 5994 4644 6012
rect 4626 6012 4644 6030
rect 4626 6030 4644 6048
rect 4626 6048 4644 6066
rect 4626 6066 4644 6084
rect 4626 6084 4644 6102
rect 4626 6102 4644 6120
rect 4626 6120 4644 6138
rect 4626 6138 4644 6156
rect 4626 6156 4644 6174
rect 4626 6174 4644 6192
rect 4626 6192 4644 6210
rect 4626 6210 4644 6228
rect 4626 6228 4644 6246
rect 4626 6246 4644 6264
rect 4626 6264 4644 6282
rect 4626 6282 4644 6300
rect 4626 6300 4644 6318
rect 4626 6318 4644 6336
rect 4626 6336 4644 6354
rect 4626 6354 4644 6372
rect 4626 6372 4644 6390
rect 4626 6390 4644 6408
rect 4626 6408 4644 6426
rect 4626 6426 4644 6444
rect 4626 6444 4644 6462
rect 4626 6462 4644 6480
rect 4626 6480 4644 6498
rect 4626 6498 4644 6516
rect 4626 6516 4644 6534
rect 4626 6534 4644 6552
rect 4626 6552 4644 6570
rect 4626 6570 4644 6588
rect 4626 6588 4644 6606
rect 4626 6606 4644 6624
rect 4626 6624 4644 6642
rect 4626 6642 4644 6660
rect 4626 6660 4644 6678
rect 4626 6678 4644 6696
rect 4626 6696 4644 6714
rect 4626 6714 4644 6732
rect 4626 6732 4644 6750
rect 4626 6750 4644 6768
rect 4626 6768 4644 6786
rect 4626 6786 4644 6804
rect 4626 6804 4644 6822
rect 4626 6822 4644 6840
rect 4626 6840 4644 6858
rect 4626 6858 4644 6876
rect 4626 6876 4644 6894
rect 4626 6894 4644 6912
rect 4626 6912 4644 6930
rect 4626 6930 4644 6948
rect 4626 6948 4644 6966
rect 4626 6966 4644 6984
rect 4626 6984 4644 7002
rect 4626 7002 4644 7020
rect 4626 7020 4644 7038
rect 4626 7038 4644 7056
rect 4626 7056 4644 7074
rect 4626 7074 4644 7092
rect 4626 7092 4644 7110
rect 4626 7110 4644 7128
rect 4626 7128 4644 7146
rect 4626 7146 4644 7164
rect 4626 7164 4644 7182
rect 4626 7182 4644 7200
rect 4626 7200 4644 7218
rect 4626 7218 4644 7236
rect 4626 7236 4644 7254
rect 4644 144 4662 162
rect 4644 162 4662 180
rect 4644 180 4662 198
rect 4644 198 4662 216
rect 4644 216 4662 234
rect 4644 234 4662 252
rect 4644 252 4662 270
rect 4644 270 4662 288
rect 4644 288 4662 306
rect 4644 306 4662 324
rect 4644 324 4662 342
rect 4644 342 4662 360
rect 4644 360 4662 378
rect 4644 378 4662 396
rect 4644 396 4662 414
rect 4644 414 4662 432
rect 4644 432 4662 450
rect 4644 450 4662 468
rect 4644 468 4662 486
rect 4644 486 4662 504
rect 4644 504 4662 522
rect 4644 522 4662 540
rect 4644 540 4662 558
rect 4644 558 4662 576
rect 4644 576 4662 594
rect 4644 594 4662 612
rect 4644 612 4662 630
rect 4644 630 4662 648
rect 4644 648 4662 666
rect 4644 666 4662 684
rect 4644 684 4662 702
rect 4644 702 4662 720
rect 4644 720 4662 738
rect 4644 738 4662 756
rect 4644 864 4662 882
rect 4644 882 4662 900
rect 4644 900 4662 918
rect 4644 918 4662 936
rect 4644 936 4662 954
rect 4644 954 4662 972
rect 4644 972 4662 990
rect 4644 990 4662 1008
rect 4644 1008 4662 1026
rect 4644 1026 4662 1044
rect 4644 1044 4662 1062
rect 4644 1062 4662 1080
rect 4644 1080 4662 1098
rect 4644 1098 4662 1116
rect 4644 1116 4662 1134
rect 4644 1134 4662 1152
rect 4644 1152 4662 1170
rect 4644 1170 4662 1188
rect 4644 1188 4662 1206
rect 4644 1206 4662 1224
rect 4644 1224 4662 1242
rect 4644 1242 4662 1260
rect 4644 1260 4662 1278
rect 4644 1278 4662 1296
rect 4644 1296 4662 1314
rect 4644 1314 4662 1332
rect 4644 1332 4662 1350
rect 4644 1350 4662 1368
rect 4644 1368 4662 1386
rect 4644 1386 4662 1404
rect 4644 1404 4662 1422
rect 4644 1422 4662 1440
rect 4644 1440 4662 1458
rect 4644 1458 4662 1476
rect 4644 1476 4662 1494
rect 4644 1494 4662 1512
rect 4644 1512 4662 1530
rect 4644 1530 4662 1548
rect 4644 1548 4662 1566
rect 4644 1566 4662 1584
rect 4644 1584 4662 1602
rect 4644 1602 4662 1620
rect 4644 1620 4662 1638
rect 4644 1638 4662 1656
rect 4644 1656 4662 1674
rect 4644 1674 4662 1692
rect 4644 1692 4662 1710
rect 4644 1710 4662 1728
rect 4644 1728 4662 1746
rect 4644 1746 4662 1764
rect 4644 1764 4662 1782
rect 4644 1782 4662 1800
rect 4644 1800 4662 1818
rect 4644 1818 4662 1836
rect 4644 1836 4662 1854
rect 4644 1854 4662 1872
rect 4644 1872 4662 1890
rect 4644 1890 4662 1908
rect 4644 1908 4662 1926
rect 4644 1926 4662 1944
rect 4644 1944 4662 1962
rect 4644 1962 4662 1980
rect 4644 1980 4662 1998
rect 4644 2232 4662 2250
rect 4644 2250 4662 2268
rect 4644 2268 4662 2286
rect 4644 2286 4662 2304
rect 4644 2304 4662 2322
rect 4644 2322 4662 2340
rect 4644 2340 4662 2358
rect 4644 2358 4662 2376
rect 4644 2376 4662 2394
rect 4644 2394 4662 2412
rect 4644 2412 4662 2430
rect 4644 2430 4662 2448
rect 4644 2448 4662 2466
rect 4644 2466 4662 2484
rect 4644 2484 4662 2502
rect 4644 2502 4662 2520
rect 4644 2520 4662 2538
rect 4644 2538 4662 2556
rect 4644 2556 4662 2574
rect 4644 2574 4662 2592
rect 4644 2592 4662 2610
rect 4644 2610 4662 2628
rect 4644 2628 4662 2646
rect 4644 2646 4662 2664
rect 4644 2664 4662 2682
rect 4644 2682 4662 2700
rect 4644 2700 4662 2718
rect 4644 2718 4662 2736
rect 4644 2736 4662 2754
rect 4644 2754 4662 2772
rect 4644 2772 4662 2790
rect 4644 2790 4662 2808
rect 4644 2808 4662 2826
rect 4644 2826 4662 2844
rect 4644 2844 4662 2862
rect 4644 2862 4662 2880
rect 4644 2880 4662 2898
rect 4644 2898 4662 2916
rect 4644 2916 4662 2934
rect 4644 2934 4662 2952
rect 4644 2952 4662 2970
rect 4644 2970 4662 2988
rect 4644 2988 4662 3006
rect 4644 3006 4662 3024
rect 4644 3024 4662 3042
rect 4644 3042 4662 3060
rect 4644 3060 4662 3078
rect 4644 3078 4662 3096
rect 4644 3096 4662 3114
rect 4644 3114 4662 3132
rect 4644 3132 4662 3150
rect 4644 3150 4662 3168
rect 4644 3168 4662 3186
rect 4644 3186 4662 3204
rect 4644 3204 4662 3222
rect 4644 3222 4662 3240
rect 4644 3240 4662 3258
rect 4644 3258 4662 3276
rect 4644 3276 4662 3294
rect 4644 3294 4662 3312
rect 4644 3312 4662 3330
rect 4644 3330 4662 3348
rect 4644 3348 4662 3366
rect 4644 3366 4662 3384
rect 4644 3384 4662 3402
rect 4644 3402 4662 3420
rect 4644 3420 4662 3438
rect 4644 3438 4662 3456
rect 4644 3456 4662 3474
rect 4644 3474 4662 3492
rect 4644 3492 4662 3510
rect 4644 3510 4662 3528
rect 4644 3528 4662 3546
rect 4644 3546 4662 3564
rect 4644 3564 4662 3582
rect 4644 3582 4662 3600
rect 4644 3600 4662 3618
rect 4644 3618 4662 3636
rect 4644 3636 4662 3654
rect 4644 3654 4662 3672
rect 4644 3672 4662 3690
rect 4644 3690 4662 3708
rect 4644 3708 4662 3726
rect 4644 3726 4662 3744
rect 4644 3744 4662 3762
rect 4644 3762 4662 3780
rect 4644 3780 4662 3798
rect 4644 3798 4662 3816
rect 4644 3816 4662 3834
rect 4644 3834 4662 3852
rect 4644 3852 4662 3870
rect 4644 3870 4662 3888
rect 4644 3888 4662 3906
rect 4644 3906 4662 3924
rect 4644 3924 4662 3942
rect 4644 3942 4662 3960
rect 4644 3960 4662 3978
rect 4644 4176 4662 4194
rect 4644 4194 4662 4212
rect 4644 4212 4662 4230
rect 4644 4230 4662 4248
rect 4644 4248 4662 4266
rect 4644 4266 4662 4284
rect 4644 4284 4662 4302
rect 4644 4302 4662 4320
rect 4644 4320 4662 4338
rect 4644 4338 4662 4356
rect 4644 4356 4662 4374
rect 4644 4374 4662 4392
rect 4644 4392 4662 4410
rect 4644 4410 4662 4428
rect 4644 4428 4662 4446
rect 4644 4446 4662 4464
rect 4644 4464 4662 4482
rect 4644 4482 4662 4500
rect 4644 4500 4662 4518
rect 4644 4518 4662 4536
rect 4644 4536 4662 4554
rect 4644 4554 4662 4572
rect 4644 4572 4662 4590
rect 4644 4590 4662 4608
rect 4644 4608 4662 4626
rect 4644 4626 4662 4644
rect 4644 4644 4662 4662
rect 4644 4662 4662 4680
rect 4644 4680 4662 4698
rect 4644 4698 4662 4716
rect 4644 4716 4662 4734
rect 4644 4734 4662 4752
rect 4644 4752 4662 4770
rect 4644 4770 4662 4788
rect 4644 4788 4662 4806
rect 4644 4806 4662 4824
rect 4644 4824 4662 4842
rect 4644 4842 4662 4860
rect 4644 4860 4662 4878
rect 4644 4878 4662 4896
rect 4644 4896 4662 4914
rect 4644 4914 4662 4932
rect 4644 4932 4662 4950
rect 4644 4950 4662 4968
rect 4644 4968 4662 4986
rect 4644 4986 4662 5004
rect 4644 5004 4662 5022
rect 4644 5022 4662 5040
rect 4644 5040 4662 5058
rect 4644 5058 4662 5076
rect 4644 5076 4662 5094
rect 4644 5094 4662 5112
rect 4644 5112 4662 5130
rect 4644 5130 4662 5148
rect 4644 5148 4662 5166
rect 4644 5166 4662 5184
rect 4644 5184 4662 5202
rect 4644 5202 4662 5220
rect 4644 5220 4662 5238
rect 4644 5238 4662 5256
rect 4644 5256 4662 5274
rect 4644 5274 4662 5292
rect 4644 5292 4662 5310
rect 4644 5310 4662 5328
rect 4644 5328 4662 5346
rect 4644 5346 4662 5364
rect 4644 5364 4662 5382
rect 4644 5382 4662 5400
rect 4644 5400 4662 5418
rect 4644 5418 4662 5436
rect 4644 5436 4662 5454
rect 4644 5454 4662 5472
rect 4644 5472 4662 5490
rect 4644 5490 4662 5508
rect 4644 5508 4662 5526
rect 4644 5526 4662 5544
rect 4644 5544 4662 5562
rect 4644 5562 4662 5580
rect 4644 5580 4662 5598
rect 4644 5598 4662 5616
rect 4644 5616 4662 5634
rect 4644 5634 4662 5652
rect 4644 5652 4662 5670
rect 4644 5670 4662 5688
rect 4644 5688 4662 5706
rect 4644 5706 4662 5724
rect 4644 5724 4662 5742
rect 4644 5742 4662 5760
rect 4644 5760 4662 5778
rect 4644 5778 4662 5796
rect 4644 5796 4662 5814
rect 4644 5814 4662 5832
rect 4644 5832 4662 5850
rect 4644 5850 4662 5868
rect 4644 5868 4662 5886
rect 4644 5886 4662 5904
rect 4644 5904 4662 5922
rect 4644 5922 4662 5940
rect 4644 5940 4662 5958
rect 4644 5958 4662 5976
rect 4644 5976 4662 5994
rect 4644 5994 4662 6012
rect 4644 6012 4662 6030
rect 4644 6030 4662 6048
rect 4644 6048 4662 6066
rect 4644 6066 4662 6084
rect 4644 6084 4662 6102
rect 4644 6102 4662 6120
rect 4644 6120 4662 6138
rect 4644 6138 4662 6156
rect 4644 6156 4662 6174
rect 4644 6174 4662 6192
rect 4644 6192 4662 6210
rect 4644 6210 4662 6228
rect 4644 6228 4662 6246
rect 4644 6246 4662 6264
rect 4644 6264 4662 6282
rect 4644 6282 4662 6300
rect 4644 6300 4662 6318
rect 4644 6318 4662 6336
rect 4644 6336 4662 6354
rect 4644 6354 4662 6372
rect 4644 6372 4662 6390
rect 4644 6390 4662 6408
rect 4644 6408 4662 6426
rect 4644 6426 4662 6444
rect 4644 6444 4662 6462
rect 4644 6462 4662 6480
rect 4644 6480 4662 6498
rect 4644 6498 4662 6516
rect 4644 6516 4662 6534
rect 4644 6534 4662 6552
rect 4644 6552 4662 6570
rect 4644 6570 4662 6588
rect 4644 6588 4662 6606
rect 4644 6606 4662 6624
rect 4644 6624 4662 6642
rect 4644 6642 4662 6660
rect 4644 6660 4662 6678
rect 4644 6678 4662 6696
rect 4644 6696 4662 6714
rect 4644 6714 4662 6732
rect 4644 6732 4662 6750
rect 4644 6750 4662 6768
rect 4644 6768 4662 6786
rect 4644 6786 4662 6804
rect 4644 6804 4662 6822
rect 4644 6822 4662 6840
rect 4644 6840 4662 6858
rect 4644 6858 4662 6876
rect 4644 6876 4662 6894
rect 4644 6894 4662 6912
rect 4644 6912 4662 6930
rect 4644 6930 4662 6948
rect 4644 6948 4662 6966
rect 4644 6966 4662 6984
rect 4644 6984 4662 7002
rect 4644 7002 4662 7020
rect 4644 7020 4662 7038
rect 4644 7038 4662 7056
rect 4644 7056 4662 7074
rect 4644 7074 4662 7092
rect 4644 7092 4662 7110
rect 4644 7110 4662 7128
rect 4644 7128 4662 7146
rect 4644 7146 4662 7164
rect 4644 7164 4662 7182
rect 4644 7182 4662 7200
rect 4644 7200 4662 7218
rect 4644 7218 4662 7236
rect 4644 7236 4662 7254
rect 4644 7254 4662 7272
rect 4644 7272 4662 7290
rect 4662 144 4680 162
rect 4662 162 4680 180
rect 4662 180 4680 198
rect 4662 198 4680 216
rect 4662 216 4680 234
rect 4662 234 4680 252
rect 4662 252 4680 270
rect 4662 270 4680 288
rect 4662 288 4680 306
rect 4662 306 4680 324
rect 4662 324 4680 342
rect 4662 342 4680 360
rect 4662 360 4680 378
rect 4662 378 4680 396
rect 4662 396 4680 414
rect 4662 414 4680 432
rect 4662 432 4680 450
rect 4662 450 4680 468
rect 4662 468 4680 486
rect 4662 486 4680 504
rect 4662 504 4680 522
rect 4662 522 4680 540
rect 4662 540 4680 558
rect 4662 558 4680 576
rect 4662 576 4680 594
rect 4662 594 4680 612
rect 4662 612 4680 630
rect 4662 630 4680 648
rect 4662 648 4680 666
rect 4662 666 4680 684
rect 4662 684 4680 702
rect 4662 702 4680 720
rect 4662 720 4680 738
rect 4662 738 4680 756
rect 4662 864 4680 882
rect 4662 882 4680 900
rect 4662 900 4680 918
rect 4662 918 4680 936
rect 4662 936 4680 954
rect 4662 954 4680 972
rect 4662 972 4680 990
rect 4662 990 4680 1008
rect 4662 1008 4680 1026
rect 4662 1026 4680 1044
rect 4662 1044 4680 1062
rect 4662 1062 4680 1080
rect 4662 1080 4680 1098
rect 4662 1098 4680 1116
rect 4662 1116 4680 1134
rect 4662 1134 4680 1152
rect 4662 1152 4680 1170
rect 4662 1170 4680 1188
rect 4662 1188 4680 1206
rect 4662 1206 4680 1224
rect 4662 1224 4680 1242
rect 4662 1242 4680 1260
rect 4662 1260 4680 1278
rect 4662 1278 4680 1296
rect 4662 1296 4680 1314
rect 4662 1314 4680 1332
rect 4662 1332 4680 1350
rect 4662 1350 4680 1368
rect 4662 1368 4680 1386
rect 4662 1386 4680 1404
rect 4662 1404 4680 1422
rect 4662 1422 4680 1440
rect 4662 1440 4680 1458
rect 4662 1458 4680 1476
rect 4662 1476 4680 1494
rect 4662 1494 4680 1512
rect 4662 1512 4680 1530
rect 4662 1530 4680 1548
rect 4662 1548 4680 1566
rect 4662 1566 4680 1584
rect 4662 1584 4680 1602
rect 4662 1602 4680 1620
rect 4662 1620 4680 1638
rect 4662 1638 4680 1656
rect 4662 1656 4680 1674
rect 4662 1674 4680 1692
rect 4662 1692 4680 1710
rect 4662 1710 4680 1728
rect 4662 1728 4680 1746
rect 4662 1746 4680 1764
rect 4662 1764 4680 1782
rect 4662 1782 4680 1800
rect 4662 1800 4680 1818
rect 4662 1818 4680 1836
rect 4662 1836 4680 1854
rect 4662 1854 4680 1872
rect 4662 1872 4680 1890
rect 4662 1890 4680 1908
rect 4662 1908 4680 1926
rect 4662 1926 4680 1944
rect 4662 1944 4680 1962
rect 4662 1962 4680 1980
rect 4662 1980 4680 1998
rect 4662 1998 4680 2016
rect 4662 2232 4680 2250
rect 4662 2250 4680 2268
rect 4662 2268 4680 2286
rect 4662 2286 4680 2304
rect 4662 2304 4680 2322
rect 4662 2322 4680 2340
rect 4662 2340 4680 2358
rect 4662 2358 4680 2376
rect 4662 2376 4680 2394
rect 4662 2394 4680 2412
rect 4662 2412 4680 2430
rect 4662 2430 4680 2448
rect 4662 2448 4680 2466
rect 4662 2466 4680 2484
rect 4662 2484 4680 2502
rect 4662 2502 4680 2520
rect 4662 2520 4680 2538
rect 4662 2538 4680 2556
rect 4662 2556 4680 2574
rect 4662 2574 4680 2592
rect 4662 2592 4680 2610
rect 4662 2610 4680 2628
rect 4662 2628 4680 2646
rect 4662 2646 4680 2664
rect 4662 2664 4680 2682
rect 4662 2682 4680 2700
rect 4662 2700 4680 2718
rect 4662 2718 4680 2736
rect 4662 2736 4680 2754
rect 4662 2754 4680 2772
rect 4662 2772 4680 2790
rect 4662 2790 4680 2808
rect 4662 2808 4680 2826
rect 4662 2826 4680 2844
rect 4662 2844 4680 2862
rect 4662 2862 4680 2880
rect 4662 2880 4680 2898
rect 4662 2898 4680 2916
rect 4662 2916 4680 2934
rect 4662 2934 4680 2952
rect 4662 2952 4680 2970
rect 4662 2970 4680 2988
rect 4662 2988 4680 3006
rect 4662 3006 4680 3024
rect 4662 3024 4680 3042
rect 4662 3042 4680 3060
rect 4662 3060 4680 3078
rect 4662 3078 4680 3096
rect 4662 3096 4680 3114
rect 4662 3114 4680 3132
rect 4662 3132 4680 3150
rect 4662 3150 4680 3168
rect 4662 3168 4680 3186
rect 4662 3186 4680 3204
rect 4662 3204 4680 3222
rect 4662 3222 4680 3240
rect 4662 3240 4680 3258
rect 4662 3258 4680 3276
rect 4662 3276 4680 3294
rect 4662 3294 4680 3312
rect 4662 3312 4680 3330
rect 4662 3330 4680 3348
rect 4662 3348 4680 3366
rect 4662 3366 4680 3384
rect 4662 3384 4680 3402
rect 4662 3402 4680 3420
rect 4662 3420 4680 3438
rect 4662 3438 4680 3456
rect 4662 3456 4680 3474
rect 4662 3474 4680 3492
rect 4662 3492 4680 3510
rect 4662 3510 4680 3528
rect 4662 3528 4680 3546
rect 4662 3546 4680 3564
rect 4662 3564 4680 3582
rect 4662 3582 4680 3600
rect 4662 3600 4680 3618
rect 4662 3618 4680 3636
rect 4662 3636 4680 3654
rect 4662 3654 4680 3672
rect 4662 3672 4680 3690
rect 4662 3690 4680 3708
rect 4662 3708 4680 3726
rect 4662 3726 4680 3744
rect 4662 3744 4680 3762
rect 4662 3762 4680 3780
rect 4662 3780 4680 3798
rect 4662 3798 4680 3816
rect 4662 3816 4680 3834
rect 4662 3834 4680 3852
rect 4662 3852 4680 3870
rect 4662 3870 4680 3888
rect 4662 3888 4680 3906
rect 4662 3906 4680 3924
rect 4662 3924 4680 3942
rect 4662 3942 4680 3960
rect 4662 3960 4680 3978
rect 4662 3978 4680 3996
rect 4662 4194 4680 4212
rect 4662 4212 4680 4230
rect 4662 4230 4680 4248
rect 4662 4248 4680 4266
rect 4662 4266 4680 4284
rect 4662 4284 4680 4302
rect 4662 4302 4680 4320
rect 4662 4320 4680 4338
rect 4662 4338 4680 4356
rect 4662 4356 4680 4374
rect 4662 4374 4680 4392
rect 4662 4392 4680 4410
rect 4662 4410 4680 4428
rect 4662 4428 4680 4446
rect 4662 4446 4680 4464
rect 4662 4464 4680 4482
rect 4662 4482 4680 4500
rect 4662 4500 4680 4518
rect 4662 4518 4680 4536
rect 4662 4536 4680 4554
rect 4662 4554 4680 4572
rect 4662 4572 4680 4590
rect 4662 4590 4680 4608
rect 4662 4608 4680 4626
rect 4662 4626 4680 4644
rect 4662 4644 4680 4662
rect 4662 4662 4680 4680
rect 4662 4680 4680 4698
rect 4662 4698 4680 4716
rect 4662 4716 4680 4734
rect 4662 4734 4680 4752
rect 4662 4752 4680 4770
rect 4662 4770 4680 4788
rect 4662 4788 4680 4806
rect 4662 4806 4680 4824
rect 4662 4824 4680 4842
rect 4662 4842 4680 4860
rect 4662 4860 4680 4878
rect 4662 4878 4680 4896
rect 4662 4896 4680 4914
rect 4662 4914 4680 4932
rect 4662 4932 4680 4950
rect 4662 4950 4680 4968
rect 4662 4968 4680 4986
rect 4662 4986 4680 5004
rect 4662 5004 4680 5022
rect 4662 5022 4680 5040
rect 4662 5040 4680 5058
rect 4662 5058 4680 5076
rect 4662 5076 4680 5094
rect 4662 5094 4680 5112
rect 4662 5112 4680 5130
rect 4662 5130 4680 5148
rect 4662 5148 4680 5166
rect 4662 5166 4680 5184
rect 4662 5184 4680 5202
rect 4662 5202 4680 5220
rect 4662 5220 4680 5238
rect 4662 5238 4680 5256
rect 4662 5256 4680 5274
rect 4662 5274 4680 5292
rect 4662 5292 4680 5310
rect 4662 5310 4680 5328
rect 4662 5328 4680 5346
rect 4662 5346 4680 5364
rect 4662 5364 4680 5382
rect 4662 5382 4680 5400
rect 4662 5400 4680 5418
rect 4662 5418 4680 5436
rect 4662 5436 4680 5454
rect 4662 5454 4680 5472
rect 4662 5472 4680 5490
rect 4662 5490 4680 5508
rect 4662 5508 4680 5526
rect 4662 5526 4680 5544
rect 4662 5544 4680 5562
rect 4662 5562 4680 5580
rect 4662 5580 4680 5598
rect 4662 5598 4680 5616
rect 4662 5616 4680 5634
rect 4662 5634 4680 5652
rect 4662 5652 4680 5670
rect 4662 5670 4680 5688
rect 4662 5688 4680 5706
rect 4662 5706 4680 5724
rect 4662 5724 4680 5742
rect 4662 5742 4680 5760
rect 4662 5760 4680 5778
rect 4662 5778 4680 5796
rect 4662 5796 4680 5814
rect 4662 5814 4680 5832
rect 4662 5832 4680 5850
rect 4662 5850 4680 5868
rect 4662 5868 4680 5886
rect 4662 5886 4680 5904
rect 4662 5904 4680 5922
rect 4662 5922 4680 5940
rect 4662 5940 4680 5958
rect 4662 5958 4680 5976
rect 4662 5976 4680 5994
rect 4662 5994 4680 6012
rect 4662 6012 4680 6030
rect 4662 6030 4680 6048
rect 4662 6048 4680 6066
rect 4662 6066 4680 6084
rect 4662 6084 4680 6102
rect 4662 6102 4680 6120
rect 4662 6120 4680 6138
rect 4662 6138 4680 6156
rect 4662 6156 4680 6174
rect 4662 6174 4680 6192
rect 4662 6192 4680 6210
rect 4662 6210 4680 6228
rect 4662 6228 4680 6246
rect 4662 6246 4680 6264
rect 4662 6264 4680 6282
rect 4662 6282 4680 6300
rect 4662 6300 4680 6318
rect 4662 6318 4680 6336
rect 4662 6336 4680 6354
rect 4662 6354 4680 6372
rect 4662 6372 4680 6390
rect 4662 6390 4680 6408
rect 4662 6408 4680 6426
rect 4662 6426 4680 6444
rect 4662 6444 4680 6462
rect 4662 6462 4680 6480
rect 4662 6480 4680 6498
rect 4662 6498 4680 6516
rect 4662 6516 4680 6534
rect 4662 6534 4680 6552
rect 4662 6552 4680 6570
rect 4662 6570 4680 6588
rect 4662 6588 4680 6606
rect 4662 6606 4680 6624
rect 4662 6624 4680 6642
rect 4662 6642 4680 6660
rect 4662 6660 4680 6678
rect 4662 6678 4680 6696
rect 4662 6696 4680 6714
rect 4662 6714 4680 6732
rect 4662 6732 4680 6750
rect 4662 6750 4680 6768
rect 4662 6768 4680 6786
rect 4662 6786 4680 6804
rect 4662 6804 4680 6822
rect 4662 6822 4680 6840
rect 4662 6840 4680 6858
rect 4662 6858 4680 6876
rect 4662 6876 4680 6894
rect 4662 6894 4680 6912
rect 4662 6912 4680 6930
rect 4662 6930 4680 6948
rect 4662 6948 4680 6966
rect 4662 6966 4680 6984
rect 4662 6984 4680 7002
rect 4662 7002 4680 7020
rect 4662 7020 4680 7038
rect 4662 7038 4680 7056
rect 4662 7056 4680 7074
rect 4662 7074 4680 7092
rect 4662 7092 4680 7110
rect 4662 7110 4680 7128
rect 4662 7128 4680 7146
rect 4662 7146 4680 7164
rect 4662 7164 4680 7182
rect 4662 7182 4680 7200
rect 4662 7200 4680 7218
rect 4662 7218 4680 7236
rect 4662 7236 4680 7254
rect 4662 7254 4680 7272
rect 4662 7272 4680 7290
rect 4662 7290 4680 7308
rect 4680 144 4698 162
rect 4680 162 4698 180
rect 4680 180 4698 198
rect 4680 198 4698 216
rect 4680 216 4698 234
rect 4680 234 4698 252
rect 4680 252 4698 270
rect 4680 270 4698 288
rect 4680 288 4698 306
rect 4680 306 4698 324
rect 4680 324 4698 342
rect 4680 342 4698 360
rect 4680 360 4698 378
rect 4680 378 4698 396
rect 4680 396 4698 414
rect 4680 414 4698 432
rect 4680 432 4698 450
rect 4680 450 4698 468
rect 4680 468 4698 486
rect 4680 486 4698 504
rect 4680 504 4698 522
rect 4680 522 4698 540
rect 4680 540 4698 558
rect 4680 558 4698 576
rect 4680 576 4698 594
rect 4680 594 4698 612
rect 4680 612 4698 630
rect 4680 630 4698 648
rect 4680 648 4698 666
rect 4680 666 4698 684
rect 4680 684 4698 702
rect 4680 702 4698 720
rect 4680 720 4698 738
rect 4680 738 4698 756
rect 4680 864 4698 882
rect 4680 882 4698 900
rect 4680 900 4698 918
rect 4680 918 4698 936
rect 4680 936 4698 954
rect 4680 954 4698 972
rect 4680 972 4698 990
rect 4680 990 4698 1008
rect 4680 1008 4698 1026
rect 4680 1026 4698 1044
rect 4680 1044 4698 1062
rect 4680 1062 4698 1080
rect 4680 1080 4698 1098
rect 4680 1098 4698 1116
rect 4680 1116 4698 1134
rect 4680 1134 4698 1152
rect 4680 1152 4698 1170
rect 4680 1170 4698 1188
rect 4680 1188 4698 1206
rect 4680 1206 4698 1224
rect 4680 1224 4698 1242
rect 4680 1242 4698 1260
rect 4680 1260 4698 1278
rect 4680 1278 4698 1296
rect 4680 1296 4698 1314
rect 4680 1314 4698 1332
rect 4680 1332 4698 1350
rect 4680 1350 4698 1368
rect 4680 1368 4698 1386
rect 4680 1386 4698 1404
rect 4680 1404 4698 1422
rect 4680 1422 4698 1440
rect 4680 1440 4698 1458
rect 4680 1458 4698 1476
rect 4680 1476 4698 1494
rect 4680 1494 4698 1512
rect 4680 1512 4698 1530
rect 4680 1530 4698 1548
rect 4680 1548 4698 1566
rect 4680 1566 4698 1584
rect 4680 1584 4698 1602
rect 4680 1602 4698 1620
rect 4680 1620 4698 1638
rect 4680 1638 4698 1656
rect 4680 1656 4698 1674
rect 4680 1674 4698 1692
rect 4680 1692 4698 1710
rect 4680 1710 4698 1728
rect 4680 1728 4698 1746
rect 4680 1746 4698 1764
rect 4680 1764 4698 1782
rect 4680 1782 4698 1800
rect 4680 1800 4698 1818
rect 4680 1818 4698 1836
rect 4680 1836 4698 1854
rect 4680 1854 4698 1872
rect 4680 1872 4698 1890
rect 4680 1890 4698 1908
rect 4680 1908 4698 1926
rect 4680 1926 4698 1944
rect 4680 1944 4698 1962
rect 4680 1962 4698 1980
rect 4680 1980 4698 1998
rect 4680 1998 4698 2016
rect 4680 2250 4698 2268
rect 4680 2268 4698 2286
rect 4680 2286 4698 2304
rect 4680 2304 4698 2322
rect 4680 2322 4698 2340
rect 4680 2340 4698 2358
rect 4680 2358 4698 2376
rect 4680 2376 4698 2394
rect 4680 2394 4698 2412
rect 4680 2412 4698 2430
rect 4680 2430 4698 2448
rect 4680 2448 4698 2466
rect 4680 2466 4698 2484
rect 4680 2484 4698 2502
rect 4680 2502 4698 2520
rect 4680 2520 4698 2538
rect 4680 2538 4698 2556
rect 4680 2556 4698 2574
rect 4680 2574 4698 2592
rect 4680 2592 4698 2610
rect 4680 2610 4698 2628
rect 4680 2628 4698 2646
rect 4680 2646 4698 2664
rect 4680 2664 4698 2682
rect 4680 2682 4698 2700
rect 4680 2700 4698 2718
rect 4680 2718 4698 2736
rect 4680 2736 4698 2754
rect 4680 2754 4698 2772
rect 4680 2772 4698 2790
rect 4680 2790 4698 2808
rect 4680 2808 4698 2826
rect 4680 2826 4698 2844
rect 4680 2844 4698 2862
rect 4680 2862 4698 2880
rect 4680 2880 4698 2898
rect 4680 2898 4698 2916
rect 4680 2916 4698 2934
rect 4680 2934 4698 2952
rect 4680 2952 4698 2970
rect 4680 2970 4698 2988
rect 4680 2988 4698 3006
rect 4680 3006 4698 3024
rect 4680 3024 4698 3042
rect 4680 3042 4698 3060
rect 4680 3060 4698 3078
rect 4680 3078 4698 3096
rect 4680 3096 4698 3114
rect 4680 3114 4698 3132
rect 4680 3132 4698 3150
rect 4680 3150 4698 3168
rect 4680 3168 4698 3186
rect 4680 3186 4698 3204
rect 4680 3204 4698 3222
rect 4680 3222 4698 3240
rect 4680 3240 4698 3258
rect 4680 3258 4698 3276
rect 4680 3276 4698 3294
rect 4680 3294 4698 3312
rect 4680 3312 4698 3330
rect 4680 3330 4698 3348
rect 4680 3348 4698 3366
rect 4680 3366 4698 3384
rect 4680 3384 4698 3402
rect 4680 3402 4698 3420
rect 4680 3420 4698 3438
rect 4680 3438 4698 3456
rect 4680 3456 4698 3474
rect 4680 3474 4698 3492
rect 4680 3492 4698 3510
rect 4680 3510 4698 3528
rect 4680 3528 4698 3546
rect 4680 3546 4698 3564
rect 4680 3564 4698 3582
rect 4680 3582 4698 3600
rect 4680 3600 4698 3618
rect 4680 3618 4698 3636
rect 4680 3636 4698 3654
rect 4680 3654 4698 3672
rect 4680 3672 4698 3690
rect 4680 3690 4698 3708
rect 4680 3708 4698 3726
rect 4680 3726 4698 3744
rect 4680 3744 4698 3762
rect 4680 3762 4698 3780
rect 4680 3780 4698 3798
rect 4680 3798 4698 3816
rect 4680 3816 4698 3834
rect 4680 3834 4698 3852
rect 4680 3852 4698 3870
rect 4680 3870 4698 3888
rect 4680 3888 4698 3906
rect 4680 3906 4698 3924
rect 4680 3924 4698 3942
rect 4680 3942 4698 3960
rect 4680 3960 4698 3978
rect 4680 3978 4698 3996
rect 4680 3996 4698 4014
rect 4680 4212 4698 4230
rect 4680 4230 4698 4248
rect 4680 4248 4698 4266
rect 4680 4266 4698 4284
rect 4680 4284 4698 4302
rect 4680 4302 4698 4320
rect 4680 4320 4698 4338
rect 4680 4338 4698 4356
rect 4680 4356 4698 4374
rect 4680 4374 4698 4392
rect 4680 4392 4698 4410
rect 4680 4410 4698 4428
rect 4680 4428 4698 4446
rect 4680 4446 4698 4464
rect 4680 4464 4698 4482
rect 4680 4482 4698 4500
rect 4680 4500 4698 4518
rect 4680 4518 4698 4536
rect 4680 4536 4698 4554
rect 4680 4554 4698 4572
rect 4680 4572 4698 4590
rect 4680 4590 4698 4608
rect 4680 4608 4698 4626
rect 4680 4626 4698 4644
rect 4680 4644 4698 4662
rect 4680 4662 4698 4680
rect 4680 4680 4698 4698
rect 4680 4698 4698 4716
rect 4680 4716 4698 4734
rect 4680 4734 4698 4752
rect 4680 4752 4698 4770
rect 4680 4770 4698 4788
rect 4680 4788 4698 4806
rect 4680 4806 4698 4824
rect 4680 4824 4698 4842
rect 4680 4842 4698 4860
rect 4680 4860 4698 4878
rect 4680 4878 4698 4896
rect 4680 4896 4698 4914
rect 4680 4914 4698 4932
rect 4680 4932 4698 4950
rect 4680 4950 4698 4968
rect 4680 4968 4698 4986
rect 4680 4986 4698 5004
rect 4680 5004 4698 5022
rect 4680 5022 4698 5040
rect 4680 5040 4698 5058
rect 4680 5058 4698 5076
rect 4680 5076 4698 5094
rect 4680 5094 4698 5112
rect 4680 5112 4698 5130
rect 4680 5130 4698 5148
rect 4680 5148 4698 5166
rect 4680 5166 4698 5184
rect 4680 5184 4698 5202
rect 4680 5202 4698 5220
rect 4680 5220 4698 5238
rect 4680 5238 4698 5256
rect 4680 5256 4698 5274
rect 4680 5274 4698 5292
rect 4680 5292 4698 5310
rect 4680 5310 4698 5328
rect 4680 5328 4698 5346
rect 4680 5346 4698 5364
rect 4680 5364 4698 5382
rect 4680 5382 4698 5400
rect 4680 5400 4698 5418
rect 4680 5418 4698 5436
rect 4680 5436 4698 5454
rect 4680 5454 4698 5472
rect 4680 5472 4698 5490
rect 4680 5490 4698 5508
rect 4680 5508 4698 5526
rect 4680 5526 4698 5544
rect 4680 5544 4698 5562
rect 4680 5562 4698 5580
rect 4680 5580 4698 5598
rect 4680 5598 4698 5616
rect 4680 5616 4698 5634
rect 4680 5634 4698 5652
rect 4680 5652 4698 5670
rect 4680 5670 4698 5688
rect 4680 5688 4698 5706
rect 4680 5706 4698 5724
rect 4680 5724 4698 5742
rect 4680 5742 4698 5760
rect 4680 5760 4698 5778
rect 4680 5778 4698 5796
rect 4680 5796 4698 5814
rect 4680 5814 4698 5832
rect 4680 5832 4698 5850
rect 4680 5850 4698 5868
rect 4680 5868 4698 5886
rect 4680 5886 4698 5904
rect 4680 5904 4698 5922
rect 4680 5922 4698 5940
rect 4680 5940 4698 5958
rect 4680 5958 4698 5976
rect 4680 5976 4698 5994
rect 4680 5994 4698 6012
rect 4680 6012 4698 6030
rect 4680 6030 4698 6048
rect 4680 6048 4698 6066
rect 4680 6066 4698 6084
rect 4680 6084 4698 6102
rect 4680 6102 4698 6120
rect 4680 6120 4698 6138
rect 4680 6138 4698 6156
rect 4680 6156 4698 6174
rect 4680 6174 4698 6192
rect 4680 6192 4698 6210
rect 4680 6210 4698 6228
rect 4680 6228 4698 6246
rect 4680 6246 4698 6264
rect 4680 6264 4698 6282
rect 4680 6282 4698 6300
rect 4680 6300 4698 6318
rect 4680 6318 4698 6336
rect 4680 6336 4698 6354
rect 4680 6354 4698 6372
rect 4680 6372 4698 6390
rect 4680 6390 4698 6408
rect 4680 6408 4698 6426
rect 4680 6426 4698 6444
rect 4680 6444 4698 6462
rect 4680 6462 4698 6480
rect 4680 6480 4698 6498
rect 4680 6498 4698 6516
rect 4680 6516 4698 6534
rect 4680 6534 4698 6552
rect 4680 6552 4698 6570
rect 4680 6570 4698 6588
rect 4680 6588 4698 6606
rect 4680 6606 4698 6624
rect 4680 6624 4698 6642
rect 4680 6642 4698 6660
rect 4680 6660 4698 6678
rect 4680 6678 4698 6696
rect 4680 6696 4698 6714
rect 4680 6714 4698 6732
rect 4680 6732 4698 6750
rect 4680 6750 4698 6768
rect 4680 6768 4698 6786
rect 4680 6786 4698 6804
rect 4680 6804 4698 6822
rect 4680 6822 4698 6840
rect 4680 6840 4698 6858
rect 4680 6858 4698 6876
rect 4680 6876 4698 6894
rect 4680 6894 4698 6912
rect 4680 6912 4698 6930
rect 4680 6930 4698 6948
rect 4680 6948 4698 6966
rect 4680 6966 4698 6984
rect 4680 6984 4698 7002
rect 4680 7002 4698 7020
rect 4680 7020 4698 7038
rect 4680 7038 4698 7056
rect 4680 7056 4698 7074
rect 4680 7074 4698 7092
rect 4680 7092 4698 7110
rect 4680 7110 4698 7128
rect 4680 7128 4698 7146
rect 4680 7146 4698 7164
rect 4680 7164 4698 7182
rect 4680 7182 4698 7200
rect 4680 7200 4698 7218
rect 4680 7218 4698 7236
rect 4680 7236 4698 7254
rect 4680 7254 4698 7272
rect 4680 7272 4698 7290
rect 4680 7290 4698 7308
rect 4680 7308 4698 7326
rect 4680 7326 4698 7344
rect 4698 162 4716 180
rect 4698 180 4716 198
rect 4698 198 4716 216
rect 4698 216 4716 234
rect 4698 234 4716 252
rect 4698 252 4716 270
rect 4698 270 4716 288
rect 4698 288 4716 306
rect 4698 306 4716 324
rect 4698 324 4716 342
rect 4698 342 4716 360
rect 4698 360 4716 378
rect 4698 378 4716 396
rect 4698 396 4716 414
rect 4698 414 4716 432
rect 4698 432 4716 450
rect 4698 450 4716 468
rect 4698 468 4716 486
rect 4698 486 4716 504
rect 4698 504 4716 522
rect 4698 522 4716 540
rect 4698 540 4716 558
rect 4698 558 4716 576
rect 4698 576 4716 594
rect 4698 594 4716 612
rect 4698 612 4716 630
rect 4698 630 4716 648
rect 4698 648 4716 666
rect 4698 666 4716 684
rect 4698 684 4716 702
rect 4698 702 4716 720
rect 4698 720 4716 738
rect 4698 738 4716 756
rect 4698 864 4716 882
rect 4698 882 4716 900
rect 4698 900 4716 918
rect 4698 918 4716 936
rect 4698 936 4716 954
rect 4698 954 4716 972
rect 4698 972 4716 990
rect 4698 990 4716 1008
rect 4698 1008 4716 1026
rect 4698 1026 4716 1044
rect 4698 1044 4716 1062
rect 4698 1062 4716 1080
rect 4698 1080 4716 1098
rect 4698 1098 4716 1116
rect 4698 1116 4716 1134
rect 4698 1134 4716 1152
rect 4698 1152 4716 1170
rect 4698 1170 4716 1188
rect 4698 1188 4716 1206
rect 4698 1206 4716 1224
rect 4698 1224 4716 1242
rect 4698 1242 4716 1260
rect 4698 1260 4716 1278
rect 4698 1278 4716 1296
rect 4698 1296 4716 1314
rect 4698 1314 4716 1332
rect 4698 1332 4716 1350
rect 4698 1350 4716 1368
rect 4698 1368 4716 1386
rect 4698 1386 4716 1404
rect 4698 1404 4716 1422
rect 4698 1422 4716 1440
rect 4698 1440 4716 1458
rect 4698 1458 4716 1476
rect 4698 1476 4716 1494
rect 4698 1494 4716 1512
rect 4698 1512 4716 1530
rect 4698 1530 4716 1548
rect 4698 1548 4716 1566
rect 4698 1566 4716 1584
rect 4698 1584 4716 1602
rect 4698 1602 4716 1620
rect 4698 1620 4716 1638
rect 4698 1638 4716 1656
rect 4698 1656 4716 1674
rect 4698 1674 4716 1692
rect 4698 1692 4716 1710
rect 4698 1710 4716 1728
rect 4698 1728 4716 1746
rect 4698 1746 4716 1764
rect 4698 1764 4716 1782
rect 4698 1782 4716 1800
rect 4698 1800 4716 1818
rect 4698 1818 4716 1836
rect 4698 1836 4716 1854
rect 4698 1854 4716 1872
rect 4698 1872 4716 1890
rect 4698 1890 4716 1908
rect 4698 1908 4716 1926
rect 4698 1926 4716 1944
rect 4698 1944 4716 1962
rect 4698 1962 4716 1980
rect 4698 1980 4716 1998
rect 4698 1998 4716 2016
rect 4698 2016 4716 2034
rect 4698 2268 4716 2286
rect 4698 2286 4716 2304
rect 4698 2304 4716 2322
rect 4698 2322 4716 2340
rect 4698 2340 4716 2358
rect 4698 2358 4716 2376
rect 4698 2376 4716 2394
rect 4698 2394 4716 2412
rect 4698 2412 4716 2430
rect 4698 2430 4716 2448
rect 4698 2448 4716 2466
rect 4698 2466 4716 2484
rect 4698 2484 4716 2502
rect 4698 2502 4716 2520
rect 4698 2520 4716 2538
rect 4698 2538 4716 2556
rect 4698 2556 4716 2574
rect 4698 2574 4716 2592
rect 4698 2592 4716 2610
rect 4698 2610 4716 2628
rect 4698 2628 4716 2646
rect 4698 2646 4716 2664
rect 4698 2664 4716 2682
rect 4698 2682 4716 2700
rect 4698 2700 4716 2718
rect 4698 2718 4716 2736
rect 4698 2736 4716 2754
rect 4698 2754 4716 2772
rect 4698 2772 4716 2790
rect 4698 2790 4716 2808
rect 4698 2808 4716 2826
rect 4698 2826 4716 2844
rect 4698 2844 4716 2862
rect 4698 2862 4716 2880
rect 4698 2880 4716 2898
rect 4698 2898 4716 2916
rect 4698 2916 4716 2934
rect 4698 2934 4716 2952
rect 4698 2952 4716 2970
rect 4698 2970 4716 2988
rect 4698 2988 4716 3006
rect 4698 3006 4716 3024
rect 4698 3024 4716 3042
rect 4698 3042 4716 3060
rect 4698 3060 4716 3078
rect 4698 3078 4716 3096
rect 4698 3096 4716 3114
rect 4698 3114 4716 3132
rect 4698 3132 4716 3150
rect 4698 3150 4716 3168
rect 4698 3168 4716 3186
rect 4698 3186 4716 3204
rect 4698 3204 4716 3222
rect 4698 3222 4716 3240
rect 4698 3240 4716 3258
rect 4698 3258 4716 3276
rect 4698 3276 4716 3294
rect 4698 3294 4716 3312
rect 4698 3312 4716 3330
rect 4698 3330 4716 3348
rect 4698 3348 4716 3366
rect 4698 3366 4716 3384
rect 4698 3384 4716 3402
rect 4698 3402 4716 3420
rect 4698 3420 4716 3438
rect 4698 3438 4716 3456
rect 4698 3456 4716 3474
rect 4698 3474 4716 3492
rect 4698 3492 4716 3510
rect 4698 3510 4716 3528
rect 4698 3528 4716 3546
rect 4698 3546 4716 3564
rect 4698 3564 4716 3582
rect 4698 3582 4716 3600
rect 4698 3600 4716 3618
rect 4698 3618 4716 3636
rect 4698 3636 4716 3654
rect 4698 3654 4716 3672
rect 4698 3672 4716 3690
rect 4698 3690 4716 3708
rect 4698 3708 4716 3726
rect 4698 3726 4716 3744
rect 4698 3744 4716 3762
rect 4698 3762 4716 3780
rect 4698 3780 4716 3798
rect 4698 3798 4716 3816
rect 4698 3816 4716 3834
rect 4698 3834 4716 3852
rect 4698 3852 4716 3870
rect 4698 3870 4716 3888
rect 4698 3888 4716 3906
rect 4698 3906 4716 3924
rect 4698 3924 4716 3942
rect 4698 3942 4716 3960
rect 4698 3960 4716 3978
rect 4698 3978 4716 3996
rect 4698 3996 4716 4014
rect 4698 4014 4716 4032
rect 4698 4248 4716 4266
rect 4698 4266 4716 4284
rect 4698 4284 4716 4302
rect 4698 4302 4716 4320
rect 4698 4320 4716 4338
rect 4698 4338 4716 4356
rect 4698 4356 4716 4374
rect 4698 4374 4716 4392
rect 4698 4392 4716 4410
rect 4698 4410 4716 4428
rect 4698 4428 4716 4446
rect 4698 4446 4716 4464
rect 4698 4464 4716 4482
rect 4698 4482 4716 4500
rect 4698 4500 4716 4518
rect 4698 4518 4716 4536
rect 4698 4536 4716 4554
rect 4698 4554 4716 4572
rect 4698 4572 4716 4590
rect 4698 4590 4716 4608
rect 4698 4608 4716 4626
rect 4698 4626 4716 4644
rect 4698 4644 4716 4662
rect 4698 4662 4716 4680
rect 4698 4680 4716 4698
rect 4698 4698 4716 4716
rect 4698 4716 4716 4734
rect 4698 4734 4716 4752
rect 4698 4752 4716 4770
rect 4698 4770 4716 4788
rect 4698 4788 4716 4806
rect 4698 4806 4716 4824
rect 4698 4824 4716 4842
rect 4698 4842 4716 4860
rect 4698 4860 4716 4878
rect 4698 4878 4716 4896
rect 4698 4896 4716 4914
rect 4698 4914 4716 4932
rect 4698 4932 4716 4950
rect 4698 4950 4716 4968
rect 4698 4968 4716 4986
rect 4698 4986 4716 5004
rect 4698 5004 4716 5022
rect 4698 5022 4716 5040
rect 4698 5040 4716 5058
rect 4698 5058 4716 5076
rect 4698 5076 4716 5094
rect 4698 5094 4716 5112
rect 4698 5112 4716 5130
rect 4698 5130 4716 5148
rect 4698 5148 4716 5166
rect 4698 5166 4716 5184
rect 4698 5184 4716 5202
rect 4698 5202 4716 5220
rect 4698 5220 4716 5238
rect 4698 5238 4716 5256
rect 4698 5256 4716 5274
rect 4698 5274 4716 5292
rect 4698 5292 4716 5310
rect 4698 5310 4716 5328
rect 4698 5328 4716 5346
rect 4698 5346 4716 5364
rect 4698 5364 4716 5382
rect 4698 5382 4716 5400
rect 4698 5400 4716 5418
rect 4698 5418 4716 5436
rect 4698 5436 4716 5454
rect 4698 5454 4716 5472
rect 4698 5472 4716 5490
rect 4698 5490 4716 5508
rect 4698 5508 4716 5526
rect 4698 5526 4716 5544
rect 4698 5544 4716 5562
rect 4698 5562 4716 5580
rect 4698 5580 4716 5598
rect 4698 5598 4716 5616
rect 4698 5616 4716 5634
rect 4698 5634 4716 5652
rect 4698 5652 4716 5670
rect 4698 5670 4716 5688
rect 4698 5688 4716 5706
rect 4698 5706 4716 5724
rect 4698 5724 4716 5742
rect 4698 5742 4716 5760
rect 4698 5760 4716 5778
rect 4698 5778 4716 5796
rect 4698 5796 4716 5814
rect 4698 5814 4716 5832
rect 4698 5832 4716 5850
rect 4698 5850 4716 5868
rect 4698 5868 4716 5886
rect 4698 5886 4716 5904
rect 4698 5904 4716 5922
rect 4698 5922 4716 5940
rect 4698 5940 4716 5958
rect 4698 5958 4716 5976
rect 4698 5976 4716 5994
rect 4698 5994 4716 6012
rect 4698 6012 4716 6030
rect 4698 6030 4716 6048
rect 4698 6048 4716 6066
rect 4698 6066 4716 6084
rect 4698 6084 4716 6102
rect 4698 6102 4716 6120
rect 4698 6120 4716 6138
rect 4698 6138 4716 6156
rect 4698 6156 4716 6174
rect 4698 6174 4716 6192
rect 4698 6192 4716 6210
rect 4698 6210 4716 6228
rect 4698 6228 4716 6246
rect 4698 6246 4716 6264
rect 4698 6264 4716 6282
rect 4698 6282 4716 6300
rect 4698 6300 4716 6318
rect 4698 6318 4716 6336
rect 4698 6336 4716 6354
rect 4698 6354 4716 6372
rect 4698 6372 4716 6390
rect 4698 6390 4716 6408
rect 4698 6408 4716 6426
rect 4698 6426 4716 6444
rect 4698 6444 4716 6462
rect 4698 6462 4716 6480
rect 4698 6480 4716 6498
rect 4698 6498 4716 6516
rect 4698 6516 4716 6534
rect 4698 6534 4716 6552
rect 4698 6552 4716 6570
rect 4698 6570 4716 6588
rect 4698 6588 4716 6606
rect 4698 6606 4716 6624
rect 4698 6624 4716 6642
rect 4698 6642 4716 6660
rect 4698 6660 4716 6678
rect 4698 6678 4716 6696
rect 4698 6696 4716 6714
rect 4698 6714 4716 6732
rect 4698 6732 4716 6750
rect 4698 6750 4716 6768
rect 4698 6768 4716 6786
rect 4698 6786 4716 6804
rect 4698 6804 4716 6822
rect 4698 6822 4716 6840
rect 4698 6840 4716 6858
rect 4698 6858 4716 6876
rect 4698 6876 4716 6894
rect 4698 6894 4716 6912
rect 4698 6912 4716 6930
rect 4698 6930 4716 6948
rect 4698 6948 4716 6966
rect 4698 6966 4716 6984
rect 4698 6984 4716 7002
rect 4698 7002 4716 7020
rect 4698 7020 4716 7038
rect 4698 7038 4716 7056
rect 4698 7056 4716 7074
rect 4698 7074 4716 7092
rect 4698 7092 4716 7110
rect 4698 7110 4716 7128
rect 4698 7128 4716 7146
rect 4698 7146 4716 7164
rect 4698 7164 4716 7182
rect 4698 7182 4716 7200
rect 4698 7200 4716 7218
rect 4698 7218 4716 7236
rect 4698 7236 4716 7254
rect 4698 7254 4716 7272
rect 4698 7272 4716 7290
rect 4698 7290 4716 7308
rect 4698 7308 4716 7326
rect 4698 7326 4716 7344
rect 4698 7344 4716 7362
rect 4698 7362 4716 7380
rect 4716 162 4734 180
rect 4716 180 4734 198
rect 4716 198 4734 216
rect 4716 216 4734 234
rect 4716 234 4734 252
rect 4716 252 4734 270
rect 4716 270 4734 288
rect 4716 288 4734 306
rect 4716 306 4734 324
rect 4716 324 4734 342
rect 4716 342 4734 360
rect 4716 360 4734 378
rect 4716 378 4734 396
rect 4716 396 4734 414
rect 4716 414 4734 432
rect 4716 432 4734 450
rect 4716 450 4734 468
rect 4716 468 4734 486
rect 4716 486 4734 504
rect 4716 504 4734 522
rect 4716 522 4734 540
rect 4716 540 4734 558
rect 4716 558 4734 576
rect 4716 576 4734 594
rect 4716 594 4734 612
rect 4716 612 4734 630
rect 4716 630 4734 648
rect 4716 648 4734 666
rect 4716 666 4734 684
rect 4716 684 4734 702
rect 4716 702 4734 720
rect 4716 720 4734 738
rect 4716 738 4734 756
rect 4716 864 4734 882
rect 4716 882 4734 900
rect 4716 900 4734 918
rect 4716 918 4734 936
rect 4716 936 4734 954
rect 4716 954 4734 972
rect 4716 972 4734 990
rect 4716 990 4734 1008
rect 4716 1008 4734 1026
rect 4716 1026 4734 1044
rect 4716 1044 4734 1062
rect 4716 1062 4734 1080
rect 4716 1080 4734 1098
rect 4716 1098 4734 1116
rect 4716 1116 4734 1134
rect 4716 1134 4734 1152
rect 4716 1152 4734 1170
rect 4716 1170 4734 1188
rect 4716 1188 4734 1206
rect 4716 1206 4734 1224
rect 4716 1224 4734 1242
rect 4716 1242 4734 1260
rect 4716 1260 4734 1278
rect 4716 1278 4734 1296
rect 4716 1296 4734 1314
rect 4716 1314 4734 1332
rect 4716 1332 4734 1350
rect 4716 1350 4734 1368
rect 4716 1368 4734 1386
rect 4716 1386 4734 1404
rect 4716 1404 4734 1422
rect 4716 1422 4734 1440
rect 4716 1440 4734 1458
rect 4716 1458 4734 1476
rect 4716 1476 4734 1494
rect 4716 1494 4734 1512
rect 4716 1512 4734 1530
rect 4716 1530 4734 1548
rect 4716 1548 4734 1566
rect 4716 1566 4734 1584
rect 4716 1584 4734 1602
rect 4716 1602 4734 1620
rect 4716 1620 4734 1638
rect 4716 1638 4734 1656
rect 4716 1656 4734 1674
rect 4716 1674 4734 1692
rect 4716 1692 4734 1710
rect 4716 1710 4734 1728
rect 4716 1728 4734 1746
rect 4716 1746 4734 1764
rect 4716 1764 4734 1782
rect 4716 1782 4734 1800
rect 4716 1800 4734 1818
rect 4716 1818 4734 1836
rect 4716 1836 4734 1854
rect 4716 1854 4734 1872
rect 4716 1872 4734 1890
rect 4716 1890 4734 1908
rect 4716 1908 4734 1926
rect 4716 1926 4734 1944
rect 4716 1944 4734 1962
rect 4716 1962 4734 1980
rect 4716 1980 4734 1998
rect 4716 1998 4734 2016
rect 4716 2016 4734 2034
rect 4716 2034 4734 2052
rect 4716 2268 4734 2286
rect 4716 2286 4734 2304
rect 4716 2304 4734 2322
rect 4716 2322 4734 2340
rect 4716 2340 4734 2358
rect 4716 2358 4734 2376
rect 4716 2376 4734 2394
rect 4716 2394 4734 2412
rect 4716 2412 4734 2430
rect 4716 2430 4734 2448
rect 4716 2448 4734 2466
rect 4716 2466 4734 2484
rect 4716 2484 4734 2502
rect 4716 2502 4734 2520
rect 4716 2520 4734 2538
rect 4716 2538 4734 2556
rect 4716 2556 4734 2574
rect 4716 2574 4734 2592
rect 4716 2592 4734 2610
rect 4716 2610 4734 2628
rect 4716 2628 4734 2646
rect 4716 2646 4734 2664
rect 4716 2664 4734 2682
rect 4716 2682 4734 2700
rect 4716 2700 4734 2718
rect 4716 2718 4734 2736
rect 4716 2736 4734 2754
rect 4716 2754 4734 2772
rect 4716 2772 4734 2790
rect 4716 2790 4734 2808
rect 4716 2808 4734 2826
rect 4716 2826 4734 2844
rect 4716 2844 4734 2862
rect 4716 2862 4734 2880
rect 4716 2880 4734 2898
rect 4716 2898 4734 2916
rect 4716 2916 4734 2934
rect 4716 2934 4734 2952
rect 4716 2952 4734 2970
rect 4716 2970 4734 2988
rect 4716 2988 4734 3006
rect 4716 3006 4734 3024
rect 4716 3024 4734 3042
rect 4716 3042 4734 3060
rect 4716 3060 4734 3078
rect 4716 3078 4734 3096
rect 4716 3096 4734 3114
rect 4716 3114 4734 3132
rect 4716 3132 4734 3150
rect 4716 3150 4734 3168
rect 4716 3168 4734 3186
rect 4716 3186 4734 3204
rect 4716 3204 4734 3222
rect 4716 3222 4734 3240
rect 4716 3240 4734 3258
rect 4716 3258 4734 3276
rect 4716 3276 4734 3294
rect 4716 3294 4734 3312
rect 4716 3312 4734 3330
rect 4716 3330 4734 3348
rect 4716 3348 4734 3366
rect 4716 3366 4734 3384
rect 4716 3384 4734 3402
rect 4716 3402 4734 3420
rect 4716 3420 4734 3438
rect 4716 3438 4734 3456
rect 4716 3456 4734 3474
rect 4716 3474 4734 3492
rect 4716 3492 4734 3510
rect 4716 3510 4734 3528
rect 4716 3528 4734 3546
rect 4716 3546 4734 3564
rect 4716 3564 4734 3582
rect 4716 3582 4734 3600
rect 4716 3600 4734 3618
rect 4716 3618 4734 3636
rect 4716 3636 4734 3654
rect 4716 3654 4734 3672
rect 4716 3672 4734 3690
rect 4716 3690 4734 3708
rect 4716 3708 4734 3726
rect 4716 3726 4734 3744
rect 4716 3744 4734 3762
rect 4716 3762 4734 3780
rect 4716 3780 4734 3798
rect 4716 3798 4734 3816
rect 4716 3816 4734 3834
rect 4716 3834 4734 3852
rect 4716 3852 4734 3870
rect 4716 3870 4734 3888
rect 4716 3888 4734 3906
rect 4716 3906 4734 3924
rect 4716 3924 4734 3942
rect 4716 3942 4734 3960
rect 4716 3960 4734 3978
rect 4716 3978 4734 3996
rect 4716 3996 4734 4014
rect 4716 4014 4734 4032
rect 4716 4032 4734 4050
rect 4716 4050 4734 4068
rect 4716 4266 4734 4284
rect 4716 4284 4734 4302
rect 4716 4302 4734 4320
rect 4716 4320 4734 4338
rect 4716 4338 4734 4356
rect 4716 4356 4734 4374
rect 4716 4374 4734 4392
rect 4716 4392 4734 4410
rect 4716 4410 4734 4428
rect 4716 4428 4734 4446
rect 4716 4446 4734 4464
rect 4716 4464 4734 4482
rect 4716 4482 4734 4500
rect 4716 4500 4734 4518
rect 4716 4518 4734 4536
rect 4716 4536 4734 4554
rect 4716 4554 4734 4572
rect 4716 4572 4734 4590
rect 4716 4590 4734 4608
rect 4716 4608 4734 4626
rect 4716 4626 4734 4644
rect 4716 4644 4734 4662
rect 4716 4662 4734 4680
rect 4716 4680 4734 4698
rect 4716 4698 4734 4716
rect 4716 4716 4734 4734
rect 4716 4734 4734 4752
rect 4716 4752 4734 4770
rect 4716 4770 4734 4788
rect 4716 4788 4734 4806
rect 4716 4806 4734 4824
rect 4716 4824 4734 4842
rect 4716 4842 4734 4860
rect 4716 4860 4734 4878
rect 4716 4878 4734 4896
rect 4716 4896 4734 4914
rect 4716 4914 4734 4932
rect 4716 4932 4734 4950
rect 4716 4950 4734 4968
rect 4716 4968 4734 4986
rect 4716 4986 4734 5004
rect 4716 5004 4734 5022
rect 4716 5022 4734 5040
rect 4716 5040 4734 5058
rect 4716 5058 4734 5076
rect 4716 5076 4734 5094
rect 4716 5094 4734 5112
rect 4716 5112 4734 5130
rect 4716 5130 4734 5148
rect 4716 5148 4734 5166
rect 4716 5166 4734 5184
rect 4716 5184 4734 5202
rect 4716 5202 4734 5220
rect 4716 5220 4734 5238
rect 4716 5238 4734 5256
rect 4716 5256 4734 5274
rect 4716 5274 4734 5292
rect 4716 5292 4734 5310
rect 4716 5310 4734 5328
rect 4716 5328 4734 5346
rect 4716 5346 4734 5364
rect 4716 5364 4734 5382
rect 4716 5382 4734 5400
rect 4716 5400 4734 5418
rect 4716 5418 4734 5436
rect 4716 5436 4734 5454
rect 4716 5454 4734 5472
rect 4716 5472 4734 5490
rect 4716 5490 4734 5508
rect 4716 5508 4734 5526
rect 4716 5526 4734 5544
rect 4716 5544 4734 5562
rect 4716 5562 4734 5580
rect 4716 5580 4734 5598
rect 4716 5598 4734 5616
rect 4716 5616 4734 5634
rect 4716 5634 4734 5652
rect 4716 5652 4734 5670
rect 4716 5670 4734 5688
rect 4716 5688 4734 5706
rect 4716 5706 4734 5724
rect 4716 5724 4734 5742
rect 4716 5742 4734 5760
rect 4716 5760 4734 5778
rect 4716 5778 4734 5796
rect 4716 5796 4734 5814
rect 4716 5814 4734 5832
rect 4716 5832 4734 5850
rect 4716 5850 4734 5868
rect 4716 5868 4734 5886
rect 4716 5886 4734 5904
rect 4716 5904 4734 5922
rect 4716 5922 4734 5940
rect 4716 5940 4734 5958
rect 4716 5958 4734 5976
rect 4716 5976 4734 5994
rect 4716 5994 4734 6012
rect 4716 6012 4734 6030
rect 4716 6030 4734 6048
rect 4716 6048 4734 6066
rect 4716 6066 4734 6084
rect 4716 6084 4734 6102
rect 4716 6102 4734 6120
rect 4716 6120 4734 6138
rect 4716 6138 4734 6156
rect 4716 6156 4734 6174
rect 4716 6174 4734 6192
rect 4716 6192 4734 6210
rect 4716 6210 4734 6228
rect 4716 6228 4734 6246
rect 4716 6246 4734 6264
rect 4716 6264 4734 6282
rect 4716 6282 4734 6300
rect 4716 6300 4734 6318
rect 4716 6318 4734 6336
rect 4716 6336 4734 6354
rect 4716 6354 4734 6372
rect 4716 6372 4734 6390
rect 4716 6390 4734 6408
rect 4716 6408 4734 6426
rect 4716 6426 4734 6444
rect 4716 6444 4734 6462
rect 4716 6462 4734 6480
rect 4716 6480 4734 6498
rect 4716 6498 4734 6516
rect 4716 6516 4734 6534
rect 4716 6534 4734 6552
rect 4716 6552 4734 6570
rect 4716 6570 4734 6588
rect 4716 6588 4734 6606
rect 4716 6606 4734 6624
rect 4716 6624 4734 6642
rect 4716 6642 4734 6660
rect 4716 6660 4734 6678
rect 4716 6678 4734 6696
rect 4716 6696 4734 6714
rect 4716 6714 4734 6732
rect 4716 6732 4734 6750
rect 4716 6750 4734 6768
rect 4716 6768 4734 6786
rect 4716 6786 4734 6804
rect 4716 6804 4734 6822
rect 4716 6822 4734 6840
rect 4716 6840 4734 6858
rect 4716 6858 4734 6876
rect 4716 6876 4734 6894
rect 4716 6894 4734 6912
rect 4716 6912 4734 6930
rect 4716 6930 4734 6948
rect 4716 6948 4734 6966
rect 4716 6966 4734 6984
rect 4716 6984 4734 7002
rect 4716 7002 4734 7020
rect 4716 7020 4734 7038
rect 4716 7038 4734 7056
rect 4716 7056 4734 7074
rect 4716 7074 4734 7092
rect 4716 7092 4734 7110
rect 4716 7110 4734 7128
rect 4716 7128 4734 7146
rect 4716 7146 4734 7164
rect 4716 7164 4734 7182
rect 4716 7182 4734 7200
rect 4716 7200 4734 7218
rect 4716 7218 4734 7236
rect 4716 7236 4734 7254
rect 4716 7254 4734 7272
rect 4716 7272 4734 7290
rect 4716 7290 4734 7308
rect 4716 7308 4734 7326
rect 4716 7326 4734 7344
rect 4716 7344 4734 7362
rect 4716 7362 4734 7380
rect 4716 7380 4734 7398
rect 4734 162 4752 180
rect 4734 180 4752 198
rect 4734 198 4752 216
rect 4734 216 4752 234
rect 4734 234 4752 252
rect 4734 252 4752 270
rect 4734 270 4752 288
rect 4734 288 4752 306
rect 4734 306 4752 324
rect 4734 324 4752 342
rect 4734 342 4752 360
rect 4734 360 4752 378
rect 4734 378 4752 396
rect 4734 396 4752 414
rect 4734 414 4752 432
rect 4734 432 4752 450
rect 4734 450 4752 468
rect 4734 468 4752 486
rect 4734 486 4752 504
rect 4734 504 4752 522
rect 4734 522 4752 540
rect 4734 540 4752 558
rect 4734 558 4752 576
rect 4734 576 4752 594
rect 4734 594 4752 612
rect 4734 612 4752 630
rect 4734 630 4752 648
rect 4734 648 4752 666
rect 4734 666 4752 684
rect 4734 684 4752 702
rect 4734 702 4752 720
rect 4734 720 4752 738
rect 4734 738 4752 756
rect 4734 864 4752 882
rect 4734 882 4752 900
rect 4734 900 4752 918
rect 4734 918 4752 936
rect 4734 936 4752 954
rect 4734 954 4752 972
rect 4734 972 4752 990
rect 4734 990 4752 1008
rect 4734 1008 4752 1026
rect 4734 1026 4752 1044
rect 4734 1044 4752 1062
rect 4734 1062 4752 1080
rect 4734 1080 4752 1098
rect 4734 1098 4752 1116
rect 4734 1116 4752 1134
rect 4734 1134 4752 1152
rect 4734 1152 4752 1170
rect 4734 1170 4752 1188
rect 4734 1188 4752 1206
rect 4734 1206 4752 1224
rect 4734 1224 4752 1242
rect 4734 1242 4752 1260
rect 4734 1260 4752 1278
rect 4734 1278 4752 1296
rect 4734 1296 4752 1314
rect 4734 1314 4752 1332
rect 4734 1332 4752 1350
rect 4734 1350 4752 1368
rect 4734 1368 4752 1386
rect 4734 1386 4752 1404
rect 4734 1404 4752 1422
rect 4734 1422 4752 1440
rect 4734 1440 4752 1458
rect 4734 1458 4752 1476
rect 4734 1476 4752 1494
rect 4734 1494 4752 1512
rect 4734 1512 4752 1530
rect 4734 1530 4752 1548
rect 4734 1548 4752 1566
rect 4734 1566 4752 1584
rect 4734 1584 4752 1602
rect 4734 1602 4752 1620
rect 4734 1620 4752 1638
rect 4734 1638 4752 1656
rect 4734 1656 4752 1674
rect 4734 1674 4752 1692
rect 4734 1692 4752 1710
rect 4734 1710 4752 1728
rect 4734 1728 4752 1746
rect 4734 1746 4752 1764
rect 4734 1764 4752 1782
rect 4734 1782 4752 1800
rect 4734 1800 4752 1818
rect 4734 1818 4752 1836
rect 4734 1836 4752 1854
rect 4734 1854 4752 1872
rect 4734 1872 4752 1890
rect 4734 1890 4752 1908
rect 4734 1908 4752 1926
rect 4734 1926 4752 1944
rect 4734 1944 4752 1962
rect 4734 1962 4752 1980
rect 4734 1980 4752 1998
rect 4734 1998 4752 2016
rect 4734 2016 4752 2034
rect 4734 2034 4752 2052
rect 4734 2286 4752 2304
rect 4734 2304 4752 2322
rect 4734 2322 4752 2340
rect 4734 2340 4752 2358
rect 4734 2358 4752 2376
rect 4734 2376 4752 2394
rect 4734 2394 4752 2412
rect 4734 2412 4752 2430
rect 4734 2430 4752 2448
rect 4734 2448 4752 2466
rect 4734 2466 4752 2484
rect 4734 2484 4752 2502
rect 4734 2502 4752 2520
rect 4734 2520 4752 2538
rect 4734 2538 4752 2556
rect 4734 2556 4752 2574
rect 4734 2574 4752 2592
rect 4734 2592 4752 2610
rect 4734 2610 4752 2628
rect 4734 2628 4752 2646
rect 4734 2646 4752 2664
rect 4734 2664 4752 2682
rect 4734 2682 4752 2700
rect 4734 2700 4752 2718
rect 4734 2718 4752 2736
rect 4734 2736 4752 2754
rect 4734 2754 4752 2772
rect 4734 2772 4752 2790
rect 4734 2790 4752 2808
rect 4734 2808 4752 2826
rect 4734 2826 4752 2844
rect 4734 2844 4752 2862
rect 4734 2862 4752 2880
rect 4734 2880 4752 2898
rect 4734 2898 4752 2916
rect 4734 2916 4752 2934
rect 4734 2934 4752 2952
rect 4734 2952 4752 2970
rect 4734 2970 4752 2988
rect 4734 2988 4752 3006
rect 4734 3006 4752 3024
rect 4734 3024 4752 3042
rect 4734 3042 4752 3060
rect 4734 3060 4752 3078
rect 4734 3078 4752 3096
rect 4734 3096 4752 3114
rect 4734 3114 4752 3132
rect 4734 3132 4752 3150
rect 4734 3150 4752 3168
rect 4734 3168 4752 3186
rect 4734 3186 4752 3204
rect 4734 3204 4752 3222
rect 4734 3222 4752 3240
rect 4734 3240 4752 3258
rect 4734 3258 4752 3276
rect 4734 3276 4752 3294
rect 4734 3294 4752 3312
rect 4734 3312 4752 3330
rect 4734 3330 4752 3348
rect 4734 3348 4752 3366
rect 4734 3366 4752 3384
rect 4734 3384 4752 3402
rect 4734 3402 4752 3420
rect 4734 3420 4752 3438
rect 4734 3438 4752 3456
rect 4734 3456 4752 3474
rect 4734 3474 4752 3492
rect 4734 3492 4752 3510
rect 4734 3510 4752 3528
rect 4734 3528 4752 3546
rect 4734 3546 4752 3564
rect 4734 3564 4752 3582
rect 4734 3582 4752 3600
rect 4734 3600 4752 3618
rect 4734 3618 4752 3636
rect 4734 3636 4752 3654
rect 4734 3654 4752 3672
rect 4734 3672 4752 3690
rect 4734 3690 4752 3708
rect 4734 3708 4752 3726
rect 4734 3726 4752 3744
rect 4734 3744 4752 3762
rect 4734 3762 4752 3780
rect 4734 3780 4752 3798
rect 4734 3798 4752 3816
rect 4734 3816 4752 3834
rect 4734 3834 4752 3852
rect 4734 3852 4752 3870
rect 4734 3870 4752 3888
rect 4734 3888 4752 3906
rect 4734 3906 4752 3924
rect 4734 3924 4752 3942
rect 4734 3942 4752 3960
rect 4734 3960 4752 3978
rect 4734 3978 4752 3996
rect 4734 3996 4752 4014
rect 4734 4014 4752 4032
rect 4734 4032 4752 4050
rect 4734 4050 4752 4068
rect 4734 4068 4752 4086
rect 4734 4284 4752 4302
rect 4734 4302 4752 4320
rect 4734 4320 4752 4338
rect 4734 4338 4752 4356
rect 4734 4356 4752 4374
rect 4734 4374 4752 4392
rect 4734 4392 4752 4410
rect 4734 4410 4752 4428
rect 4734 4428 4752 4446
rect 4734 4446 4752 4464
rect 4734 4464 4752 4482
rect 4734 4482 4752 4500
rect 4734 4500 4752 4518
rect 4734 4518 4752 4536
rect 4734 4536 4752 4554
rect 4734 4554 4752 4572
rect 4734 4572 4752 4590
rect 4734 4590 4752 4608
rect 4734 4608 4752 4626
rect 4734 4626 4752 4644
rect 4734 4644 4752 4662
rect 4734 4662 4752 4680
rect 4734 4680 4752 4698
rect 4734 4698 4752 4716
rect 4734 4716 4752 4734
rect 4734 4734 4752 4752
rect 4734 4752 4752 4770
rect 4734 4770 4752 4788
rect 4734 4788 4752 4806
rect 4734 4806 4752 4824
rect 4734 4824 4752 4842
rect 4734 4842 4752 4860
rect 4734 4860 4752 4878
rect 4734 4878 4752 4896
rect 4734 4896 4752 4914
rect 4734 4914 4752 4932
rect 4734 4932 4752 4950
rect 4734 4950 4752 4968
rect 4734 4968 4752 4986
rect 4734 4986 4752 5004
rect 4734 5004 4752 5022
rect 4734 5022 4752 5040
rect 4734 5040 4752 5058
rect 4734 5058 4752 5076
rect 4734 5076 4752 5094
rect 4734 5094 4752 5112
rect 4734 5112 4752 5130
rect 4734 5130 4752 5148
rect 4734 5148 4752 5166
rect 4734 5166 4752 5184
rect 4734 5184 4752 5202
rect 4734 5202 4752 5220
rect 4734 5220 4752 5238
rect 4734 5238 4752 5256
rect 4734 5256 4752 5274
rect 4734 5274 4752 5292
rect 4734 5292 4752 5310
rect 4734 5310 4752 5328
rect 4734 5328 4752 5346
rect 4734 5346 4752 5364
rect 4734 5364 4752 5382
rect 4734 5382 4752 5400
rect 4734 5400 4752 5418
rect 4734 5418 4752 5436
rect 4734 5436 4752 5454
rect 4734 5454 4752 5472
rect 4734 5472 4752 5490
rect 4734 5490 4752 5508
rect 4734 5508 4752 5526
rect 4734 5526 4752 5544
rect 4734 5544 4752 5562
rect 4734 5562 4752 5580
rect 4734 5580 4752 5598
rect 4734 5598 4752 5616
rect 4734 5616 4752 5634
rect 4734 5634 4752 5652
rect 4734 5652 4752 5670
rect 4734 5670 4752 5688
rect 4734 5688 4752 5706
rect 4734 5706 4752 5724
rect 4734 5724 4752 5742
rect 4734 5742 4752 5760
rect 4734 5760 4752 5778
rect 4734 5778 4752 5796
rect 4734 5796 4752 5814
rect 4734 5814 4752 5832
rect 4734 5832 4752 5850
rect 4734 5850 4752 5868
rect 4734 5868 4752 5886
rect 4734 5886 4752 5904
rect 4734 5904 4752 5922
rect 4734 5922 4752 5940
rect 4734 5940 4752 5958
rect 4734 5958 4752 5976
rect 4734 5976 4752 5994
rect 4734 5994 4752 6012
rect 4734 6012 4752 6030
rect 4734 6030 4752 6048
rect 4734 6048 4752 6066
rect 4734 6066 4752 6084
rect 4734 6084 4752 6102
rect 4734 6102 4752 6120
rect 4734 6120 4752 6138
rect 4734 6138 4752 6156
rect 4734 6156 4752 6174
rect 4734 6174 4752 6192
rect 4734 6192 4752 6210
rect 4734 6210 4752 6228
rect 4734 6228 4752 6246
rect 4734 6246 4752 6264
rect 4734 6264 4752 6282
rect 4734 6282 4752 6300
rect 4734 6300 4752 6318
rect 4734 6318 4752 6336
rect 4734 6336 4752 6354
rect 4734 6354 4752 6372
rect 4734 6372 4752 6390
rect 4734 6390 4752 6408
rect 4734 6408 4752 6426
rect 4734 6426 4752 6444
rect 4734 6444 4752 6462
rect 4734 6462 4752 6480
rect 4734 6480 4752 6498
rect 4734 6498 4752 6516
rect 4734 6516 4752 6534
rect 4734 6534 4752 6552
rect 4734 6552 4752 6570
rect 4734 6570 4752 6588
rect 4734 6588 4752 6606
rect 4734 6606 4752 6624
rect 4734 6624 4752 6642
rect 4734 6642 4752 6660
rect 4734 6660 4752 6678
rect 4734 6678 4752 6696
rect 4734 6696 4752 6714
rect 4734 6714 4752 6732
rect 4734 6732 4752 6750
rect 4734 6750 4752 6768
rect 4734 6768 4752 6786
rect 4734 6786 4752 6804
rect 4734 6804 4752 6822
rect 4734 6822 4752 6840
rect 4734 6840 4752 6858
rect 4734 6858 4752 6876
rect 4734 6876 4752 6894
rect 4734 6894 4752 6912
rect 4734 6912 4752 6930
rect 4734 6930 4752 6948
rect 4734 6948 4752 6966
rect 4734 6966 4752 6984
rect 4734 6984 4752 7002
rect 4734 7002 4752 7020
rect 4734 7020 4752 7038
rect 4734 7038 4752 7056
rect 4734 7056 4752 7074
rect 4734 7074 4752 7092
rect 4734 7092 4752 7110
rect 4734 7110 4752 7128
rect 4734 7128 4752 7146
rect 4734 7146 4752 7164
rect 4734 7164 4752 7182
rect 4734 7182 4752 7200
rect 4734 7200 4752 7218
rect 4734 7218 4752 7236
rect 4734 7236 4752 7254
rect 4734 7254 4752 7272
rect 4734 7272 4752 7290
rect 4734 7290 4752 7308
rect 4734 7308 4752 7326
rect 4734 7326 4752 7344
rect 4734 7344 4752 7362
rect 4734 7362 4752 7380
rect 4734 7380 4752 7398
rect 4734 7398 4752 7416
rect 4734 7416 4752 7434
rect 4752 180 4770 198
rect 4752 198 4770 216
rect 4752 216 4770 234
rect 4752 234 4770 252
rect 4752 252 4770 270
rect 4752 270 4770 288
rect 4752 288 4770 306
rect 4752 306 4770 324
rect 4752 324 4770 342
rect 4752 342 4770 360
rect 4752 360 4770 378
rect 4752 378 4770 396
rect 4752 396 4770 414
rect 4752 414 4770 432
rect 4752 432 4770 450
rect 4752 450 4770 468
rect 4752 468 4770 486
rect 4752 486 4770 504
rect 4752 504 4770 522
rect 4752 522 4770 540
rect 4752 540 4770 558
rect 4752 558 4770 576
rect 4752 576 4770 594
rect 4752 594 4770 612
rect 4752 612 4770 630
rect 4752 630 4770 648
rect 4752 648 4770 666
rect 4752 666 4770 684
rect 4752 684 4770 702
rect 4752 702 4770 720
rect 4752 720 4770 738
rect 4752 738 4770 756
rect 4752 864 4770 882
rect 4752 882 4770 900
rect 4752 900 4770 918
rect 4752 918 4770 936
rect 4752 936 4770 954
rect 4752 954 4770 972
rect 4752 972 4770 990
rect 4752 990 4770 1008
rect 4752 1008 4770 1026
rect 4752 1026 4770 1044
rect 4752 1044 4770 1062
rect 4752 1062 4770 1080
rect 4752 1080 4770 1098
rect 4752 1098 4770 1116
rect 4752 1116 4770 1134
rect 4752 1134 4770 1152
rect 4752 1152 4770 1170
rect 4752 1170 4770 1188
rect 4752 1188 4770 1206
rect 4752 1206 4770 1224
rect 4752 1224 4770 1242
rect 4752 1242 4770 1260
rect 4752 1260 4770 1278
rect 4752 1278 4770 1296
rect 4752 1296 4770 1314
rect 4752 1314 4770 1332
rect 4752 1332 4770 1350
rect 4752 1350 4770 1368
rect 4752 1368 4770 1386
rect 4752 1386 4770 1404
rect 4752 1404 4770 1422
rect 4752 1422 4770 1440
rect 4752 1440 4770 1458
rect 4752 1458 4770 1476
rect 4752 1476 4770 1494
rect 4752 1494 4770 1512
rect 4752 1512 4770 1530
rect 4752 1530 4770 1548
rect 4752 1548 4770 1566
rect 4752 1566 4770 1584
rect 4752 1584 4770 1602
rect 4752 1602 4770 1620
rect 4752 1620 4770 1638
rect 4752 1638 4770 1656
rect 4752 1656 4770 1674
rect 4752 1674 4770 1692
rect 4752 1692 4770 1710
rect 4752 1710 4770 1728
rect 4752 1728 4770 1746
rect 4752 1746 4770 1764
rect 4752 1764 4770 1782
rect 4752 1782 4770 1800
rect 4752 1800 4770 1818
rect 4752 1818 4770 1836
rect 4752 1836 4770 1854
rect 4752 1854 4770 1872
rect 4752 1872 4770 1890
rect 4752 1890 4770 1908
rect 4752 1908 4770 1926
rect 4752 1926 4770 1944
rect 4752 1944 4770 1962
rect 4752 1962 4770 1980
rect 4752 1980 4770 1998
rect 4752 1998 4770 2016
rect 4752 2016 4770 2034
rect 4752 2034 4770 2052
rect 4752 2052 4770 2070
rect 4752 2304 4770 2322
rect 4752 2322 4770 2340
rect 4752 2340 4770 2358
rect 4752 2358 4770 2376
rect 4752 2376 4770 2394
rect 4752 2394 4770 2412
rect 4752 2412 4770 2430
rect 4752 2430 4770 2448
rect 4752 2448 4770 2466
rect 4752 2466 4770 2484
rect 4752 2484 4770 2502
rect 4752 2502 4770 2520
rect 4752 2520 4770 2538
rect 4752 2538 4770 2556
rect 4752 2556 4770 2574
rect 4752 2574 4770 2592
rect 4752 2592 4770 2610
rect 4752 2610 4770 2628
rect 4752 2628 4770 2646
rect 4752 2646 4770 2664
rect 4752 2664 4770 2682
rect 4752 2682 4770 2700
rect 4752 2700 4770 2718
rect 4752 2718 4770 2736
rect 4752 2736 4770 2754
rect 4752 2754 4770 2772
rect 4752 2772 4770 2790
rect 4752 2790 4770 2808
rect 4752 2808 4770 2826
rect 4752 2826 4770 2844
rect 4752 2844 4770 2862
rect 4752 2862 4770 2880
rect 4752 2880 4770 2898
rect 4752 2898 4770 2916
rect 4752 2916 4770 2934
rect 4752 2934 4770 2952
rect 4752 2952 4770 2970
rect 4752 2970 4770 2988
rect 4752 2988 4770 3006
rect 4752 3006 4770 3024
rect 4752 3024 4770 3042
rect 4752 3042 4770 3060
rect 4752 3060 4770 3078
rect 4752 3078 4770 3096
rect 4752 3096 4770 3114
rect 4752 3114 4770 3132
rect 4752 3132 4770 3150
rect 4752 3150 4770 3168
rect 4752 3168 4770 3186
rect 4752 3186 4770 3204
rect 4752 3204 4770 3222
rect 4752 3222 4770 3240
rect 4752 3240 4770 3258
rect 4752 3258 4770 3276
rect 4752 3276 4770 3294
rect 4752 3294 4770 3312
rect 4752 3312 4770 3330
rect 4752 3330 4770 3348
rect 4752 3348 4770 3366
rect 4752 3366 4770 3384
rect 4752 3384 4770 3402
rect 4752 3402 4770 3420
rect 4752 3420 4770 3438
rect 4752 3438 4770 3456
rect 4752 3456 4770 3474
rect 4752 3474 4770 3492
rect 4752 3492 4770 3510
rect 4752 3510 4770 3528
rect 4752 3528 4770 3546
rect 4752 3546 4770 3564
rect 4752 3564 4770 3582
rect 4752 3582 4770 3600
rect 4752 3600 4770 3618
rect 4752 3618 4770 3636
rect 4752 3636 4770 3654
rect 4752 3654 4770 3672
rect 4752 3672 4770 3690
rect 4752 3690 4770 3708
rect 4752 3708 4770 3726
rect 4752 3726 4770 3744
rect 4752 3744 4770 3762
rect 4752 3762 4770 3780
rect 4752 3780 4770 3798
rect 4752 3798 4770 3816
rect 4752 3816 4770 3834
rect 4752 3834 4770 3852
rect 4752 3852 4770 3870
rect 4752 3870 4770 3888
rect 4752 3888 4770 3906
rect 4752 3906 4770 3924
rect 4752 3924 4770 3942
rect 4752 3942 4770 3960
rect 4752 3960 4770 3978
rect 4752 3978 4770 3996
rect 4752 3996 4770 4014
rect 4752 4014 4770 4032
rect 4752 4032 4770 4050
rect 4752 4050 4770 4068
rect 4752 4068 4770 4086
rect 4752 4086 4770 4104
rect 4752 4302 4770 4320
rect 4752 4320 4770 4338
rect 4752 4338 4770 4356
rect 4752 4356 4770 4374
rect 4752 4374 4770 4392
rect 4752 4392 4770 4410
rect 4752 4410 4770 4428
rect 4752 4428 4770 4446
rect 4752 4446 4770 4464
rect 4752 4464 4770 4482
rect 4752 4482 4770 4500
rect 4752 4500 4770 4518
rect 4752 4518 4770 4536
rect 4752 4536 4770 4554
rect 4752 4554 4770 4572
rect 4752 4572 4770 4590
rect 4752 4590 4770 4608
rect 4752 4608 4770 4626
rect 4752 4626 4770 4644
rect 4752 4644 4770 4662
rect 4752 4662 4770 4680
rect 4752 4680 4770 4698
rect 4752 4698 4770 4716
rect 4752 4716 4770 4734
rect 4752 4734 4770 4752
rect 4752 4752 4770 4770
rect 4752 4770 4770 4788
rect 4752 4788 4770 4806
rect 4752 4806 4770 4824
rect 4752 4824 4770 4842
rect 4752 4842 4770 4860
rect 4752 4860 4770 4878
rect 4752 4878 4770 4896
rect 4752 4896 4770 4914
rect 4752 4914 4770 4932
rect 4752 4932 4770 4950
rect 4752 4950 4770 4968
rect 4752 4968 4770 4986
rect 4752 4986 4770 5004
rect 4752 5004 4770 5022
rect 4752 5022 4770 5040
rect 4752 5040 4770 5058
rect 4752 5058 4770 5076
rect 4752 5076 4770 5094
rect 4752 5094 4770 5112
rect 4752 5112 4770 5130
rect 4752 5130 4770 5148
rect 4752 5148 4770 5166
rect 4752 5166 4770 5184
rect 4752 5184 4770 5202
rect 4752 5202 4770 5220
rect 4752 5220 4770 5238
rect 4752 5238 4770 5256
rect 4752 5256 4770 5274
rect 4752 5274 4770 5292
rect 4752 5292 4770 5310
rect 4752 5310 4770 5328
rect 4752 5328 4770 5346
rect 4752 5346 4770 5364
rect 4752 5364 4770 5382
rect 4752 5382 4770 5400
rect 4752 5400 4770 5418
rect 4752 5418 4770 5436
rect 4752 5436 4770 5454
rect 4752 5454 4770 5472
rect 4752 5472 4770 5490
rect 4752 5490 4770 5508
rect 4752 5508 4770 5526
rect 4752 5526 4770 5544
rect 4752 5544 4770 5562
rect 4752 5562 4770 5580
rect 4752 5580 4770 5598
rect 4752 5598 4770 5616
rect 4752 5616 4770 5634
rect 4752 5634 4770 5652
rect 4752 5652 4770 5670
rect 4752 5670 4770 5688
rect 4752 5688 4770 5706
rect 4752 5706 4770 5724
rect 4752 5724 4770 5742
rect 4752 5742 4770 5760
rect 4752 5760 4770 5778
rect 4752 5778 4770 5796
rect 4752 5796 4770 5814
rect 4752 5814 4770 5832
rect 4752 5832 4770 5850
rect 4752 5850 4770 5868
rect 4752 5868 4770 5886
rect 4752 5886 4770 5904
rect 4752 5904 4770 5922
rect 4752 5922 4770 5940
rect 4752 5940 4770 5958
rect 4752 5958 4770 5976
rect 4752 5976 4770 5994
rect 4752 5994 4770 6012
rect 4752 6012 4770 6030
rect 4752 6030 4770 6048
rect 4752 6048 4770 6066
rect 4752 6066 4770 6084
rect 4752 6084 4770 6102
rect 4752 6102 4770 6120
rect 4752 6120 4770 6138
rect 4752 6138 4770 6156
rect 4752 6156 4770 6174
rect 4752 6174 4770 6192
rect 4752 6192 4770 6210
rect 4752 6210 4770 6228
rect 4752 6228 4770 6246
rect 4752 6246 4770 6264
rect 4752 6264 4770 6282
rect 4752 6282 4770 6300
rect 4752 6300 4770 6318
rect 4752 6318 4770 6336
rect 4752 6336 4770 6354
rect 4752 6354 4770 6372
rect 4752 6372 4770 6390
rect 4752 6390 4770 6408
rect 4752 6408 4770 6426
rect 4752 6426 4770 6444
rect 4752 6444 4770 6462
rect 4752 6462 4770 6480
rect 4752 6480 4770 6498
rect 4752 6498 4770 6516
rect 4752 6516 4770 6534
rect 4752 6534 4770 6552
rect 4752 6552 4770 6570
rect 4752 6570 4770 6588
rect 4752 6588 4770 6606
rect 4752 6606 4770 6624
rect 4752 6624 4770 6642
rect 4752 6642 4770 6660
rect 4752 6660 4770 6678
rect 4752 6678 4770 6696
rect 4752 6696 4770 6714
rect 4752 6714 4770 6732
rect 4752 6732 4770 6750
rect 4752 6750 4770 6768
rect 4752 6768 4770 6786
rect 4752 6786 4770 6804
rect 4752 6804 4770 6822
rect 4752 6822 4770 6840
rect 4752 6840 4770 6858
rect 4752 6858 4770 6876
rect 4752 6876 4770 6894
rect 4752 6894 4770 6912
rect 4752 6912 4770 6930
rect 4752 6930 4770 6948
rect 4752 6948 4770 6966
rect 4752 6966 4770 6984
rect 4752 6984 4770 7002
rect 4752 7002 4770 7020
rect 4752 7020 4770 7038
rect 4752 7038 4770 7056
rect 4752 7056 4770 7074
rect 4752 7074 4770 7092
rect 4752 7092 4770 7110
rect 4752 7110 4770 7128
rect 4752 7128 4770 7146
rect 4752 7146 4770 7164
rect 4752 7164 4770 7182
rect 4752 7182 4770 7200
rect 4752 7200 4770 7218
rect 4752 7218 4770 7236
rect 4752 7236 4770 7254
rect 4752 7254 4770 7272
rect 4752 7272 4770 7290
rect 4752 7290 4770 7308
rect 4752 7308 4770 7326
rect 4752 7326 4770 7344
rect 4752 7344 4770 7362
rect 4752 7362 4770 7380
rect 4752 7380 4770 7398
rect 4752 7398 4770 7416
rect 4752 7416 4770 7434
rect 4752 7434 4770 7452
rect 4770 180 4788 198
rect 4770 198 4788 216
rect 4770 216 4788 234
rect 4770 234 4788 252
rect 4770 252 4788 270
rect 4770 270 4788 288
rect 4770 288 4788 306
rect 4770 306 4788 324
rect 4770 324 4788 342
rect 4770 342 4788 360
rect 4770 360 4788 378
rect 4770 378 4788 396
rect 4770 396 4788 414
rect 4770 414 4788 432
rect 4770 432 4788 450
rect 4770 450 4788 468
rect 4770 468 4788 486
rect 4770 486 4788 504
rect 4770 504 4788 522
rect 4770 522 4788 540
rect 4770 540 4788 558
rect 4770 558 4788 576
rect 4770 576 4788 594
rect 4770 594 4788 612
rect 4770 612 4788 630
rect 4770 630 4788 648
rect 4770 648 4788 666
rect 4770 666 4788 684
rect 4770 684 4788 702
rect 4770 702 4788 720
rect 4770 720 4788 738
rect 4770 738 4788 756
rect 4770 864 4788 882
rect 4770 882 4788 900
rect 4770 900 4788 918
rect 4770 918 4788 936
rect 4770 936 4788 954
rect 4770 954 4788 972
rect 4770 972 4788 990
rect 4770 990 4788 1008
rect 4770 1008 4788 1026
rect 4770 1026 4788 1044
rect 4770 1044 4788 1062
rect 4770 1062 4788 1080
rect 4770 1080 4788 1098
rect 4770 1098 4788 1116
rect 4770 1116 4788 1134
rect 4770 1134 4788 1152
rect 4770 1152 4788 1170
rect 4770 1170 4788 1188
rect 4770 1188 4788 1206
rect 4770 1206 4788 1224
rect 4770 1224 4788 1242
rect 4770 1242 4788 1260
rect 4770 1260 4788 1278
rect 4770 1278 4788 1296
rect 4770 1296 4788 1314
rect 4770 1314 4788 1332
rect 4770 1332 4788 1350
rect 4770 1350 4788 1368
rect 4770 1368 4788 1386
rect 4770 1386 4788 1404
rect 4770 1404 4788 1422
rect 4770 1422 4788 1440
rect 4770 1440 4788 1458
rect 4770 1458 4788 1476
rect 4770 1476 4788 1494
rect 4770 1494 4788 1512
rect 4770 1512 4788 1530
rect 4770 1530 4788 1548
rect 4770 1548 4788 1566
rect 4770 1566 4788 1584
rect 4770 1584 4788 1602
rect 4770 1602 4788 1620
rect 4770 1620 4788 1638
rect 4770 1638 4788 1656
rect 4770 1656 4788 1674
rect 4770 1674 4788 1692
rect 4770 1692 4788 1710
rect 4770 1710 4788 1728
rect 4770 1728 4788 1746
rect 4770 1746 4788 1764
rect 4770 1764 4788 1782
rect 4770 1782 4788 1800
rect 4770 1800 4788 1818
rect 4770 1818 4788 1836
rect 4770 1836 4788 1854
rect 4770 1854 4788 1872
rect 4770 1872 4788 1890
rect 4770 1890 4788 1908
rect 4770 1908 4788 1926
rect 4770 1926 4788 1944
rect 4770 1944 4788 1962
rect 4770 1962 4788 1980
rect 4770 1980 4788 1998
rect 4770 1998 4788 2016
rect 4770 2016 4788 2034
rect 4770 2034 4788 2052
rect 4770 2052 4788 2070
rect 4770 2070 4788 2088
rect 4770 2304 4788 2322
rect 4770 2322 4788 2340
rect 4770 2340 4788 2358
rect 4770 2358 4788 2376
rect 4770 2376 4788 2394
rect 4770 2394 4788 2412
rect 4770 2412 4788 2430
rect 4770 2430 4788 2448
rect 4770 2448 4788 2466
rect 4770 2466 4788 2484
rect 4770 2484 4788 2502
rect 4770 2502 4788 2520
rect 4770 2520 4788 2538
rect 4770 2538 4788 2556
rect 4770 2556 4788 2574
rect 4770 2574 4788 2592
rect 4770 2592 4788 2610
rect 4770 2610 4788 2628
rect 4770 2628 4788 2646
rect 4770 2646 4788 2664
rect 4770 2664 4788 2682
rect 4770 2682 4788 2700
rect 4770 2700 4788 2718
rect 4770 2718 4788 2736
rect 4770 2736 4788 2754
rect 4770 2754 4788 2772
rect 4770 2772 4788 2790
rect 4770 2790 4788 2808
rect 4770 2808 4788 2826
rect 4770 2826 4788 2844
rect 4770 2844 4788 2862
rect 4770 2862 4788 2880
rect 4770 2880 4788 2898
rect 4770 2898 4788 2916
rect 4770 2916 4788 2934
rect 4770 2934 4788 2952
rect 4770 2952 4788 2970
rect 4770 2970 4788 2988
rect 4770 2988 4788 3006
rect 4770 3006 4788 3024
rect 4770 3024 4788 3042
rect 4770 3042 4788 3060
rect 4770 3060 4788 3078
rect 4770 3078 4788 3096
rect 4770 3096 4788 3114
rect 4770 3114 4788 3132
rect 4770 3132 4788 3150
rect 4770 3150 4788 3168
rect 4770 3168 4788 3186
rect 4770 3186 4788 3204
rect 4770 3204 4788 3222
rect 4770 3222 4788 3240
rect 4770 3240 4788 3258
rect 4770 3258 4788 3276
rect 4770 3276 4788 3294
rect 4770 3294 4788 3312
rect 4770 3312 4788 3330
rect 4770 3330 4788 3348
rect 4770 3348 4788 3366
rect 4770 3366 4788 3384
rect 4770 3384 4788 3402
rect 4770 3402 4788 3420
rect 4770 3420 4788 3438
rect 4770 3438 4788 3456
rect 4770 3456 4788 3474
rect 4770 3474 4788 3492
rect 4770 3492 4788 3510
rect 4770 3510 4788 3528
rect 4770 3528 4788 3546
rect 4770 3546 4788 3564
rect 4770 3564 4788 3582
rect 4770 3582 4788 3600
rect 4770 3600 4788 3618
rect 4770 3618 4788 3636
rect 4770 3636 4788 3654
rect 4770 3654 4788 3672
rect 4770 3672 4788 3690
rect 4770 3690 4788 3708
rect 4770 3708 4788 3726
rect 4770 3726 4788 3744
rect 4770 3744 4788 3762
rect 4770 3762 4788 3780
rect 4770 3780 4788 3798
rect 4770 3798 4788 3816
rect 4770 3816 4788 3834
rect 4770 3834 4788 3852
rect 4770 3852 4788 3870
rect 4770 3870 4788 3888
rect 4770 3888 4788 3906
rect 4770 3906 4788 3924
rect 4770 3924 4788 3942
rect 4770 3942 4788 3960
rect 4770 3960 4788 3978
rect 4770 3978 4788 3996
rect 4770 3996 4788 4014
rect 4770 4014 4788 4032
rect 4770 4032 4788 4050
rect 4770 4050 4788 4068
rect 4770 4068 4788 4086
rect 4770 4086 4788 4104
rect 4770 4104 4788 4122
rect 4770 4320 4788 4338
rect 4770 4338 4788 4356
rect 4770 4356 4788 4374
rect 4770 4374 4788 4392
rect 4770 4392 4788 4410
rect 4770 4410 4788 4428
rect 4770 4428 4788 4446
rect 4770 4446 4788 4464
rect 4770 4464 4788 4482
rect 4770 4482 4788 4500
rect 4770 4500 4788 4518
rect 4770 4518 4788 4536
rect 4770 4536 4788 4554
rect 4770 4554 4788 4572
rect 4770 4572 4788 4590
rect 4770 4590 4788 4608
rect 4770 4608 4788 4626
rect 4770 4626 4788 4644
rect 4770 4644 4788 4662
rect 4770 4662 4788 4680
rect 4770 4680 4788 4698
rect 4770 4698 4788 4716
rect 4770 4716 4788 4734
rect 4770 4734 4788 4752
rect 4770 4752 4788 4770
rect 4770 4770 4788 4788
rect 4770 4788 4788 4806
rect 4770 4806 4788 4824
rect 4770 4824 4788 4842
rect 4770 4842 4788 4860
rect 4770 4860 4788 4878
rect 4770 4878 4788 4896
rect 4770 4896 4788 4914
rect 4770 4914 4788 4932
rect 4770 4932 4788 4950
rect 4770 4950 4788 4968
rect 4770 4968 4788 4986
rect 4770 4986 4788 5004
rect 4770 5004 4788 5022
rect 4770 5022 4788 5040
rect 4770 5040 4788 5058
rect 4770 5058 4788 5076
rect 4770 5076 4788 5094
rect 4770 5094 4788 5112
rect 4770 5112 4788 5130
rect 4770 5130 4788 5148
rect 4770 5148 4788 5166
rect 4770 5166 4788 5184
rect 4770 5184 4788 5202
rect 4770 5202 4788 5220
rect 4770 5220 4788 5238
rect 4770 5238 4788 5256
rect 4770 5256 4788 5274
rect 4770 5274 4788 5292
rect 4770 5292 4788 5310
rect 4770 5310 4788 5328
rect 4770 5328 4788 5346
rect 4770 5346 4788 5364
rect 4770 5364 4788 5382
rect 4770 5382 4788 5400
rect 4770 5400 4788 5418
rect 4770 5418 4788 5436
rect 4770 5436 4788 5454
rect 4770 5454 4788 5472
rect 4770 5472 4788 5490
rect 4770 5490 4788 5508
rect 4770 5508 4788 5526
rect 4770 5526 4788 5544
rect 4770 5544 4788 5562
rect 4770 5562 4788 5580
rect 4770 5580 4788 5598
rect 4770 5598 4788 5616
rect 4770 5616 4788 5634
rect 4770 5634 4788 5652
rect 4770 5652 4788 5670
rect 4770 5670 4788 5688
rect 4770 5688 4788 5706
rect 4770 5706 4788 5724
rect 4770 5724 4788 5742
rect 4770 5742 4788 5760
rect 4770 5760 4788 5778
rect 4770 5778 4788 5796
rect 4770 5796 4788 5814
rect 4770 5814 4788 5832
rect 4770 5832 4788 5850
rect 4770 5850 4788 5868
rect 4770 5868 4788 5886
rect 4770 5886 4788 5904
rect 4770 5904 4788 5922
rect 4770 5922 4788 5940
rect 4770 5940 4788 5958
rect 4770 5958 4788 5976
rect 4770 5976 4788 5994
rect 4770 5994 4788 6012
rect 4770 6012 4788 6030
rect 4770 6030 4788 6048
rect 4770 6048 4788 6066
rect 4770 6066 4788 6084
rect 4770 6084 4788 6102
rect 4770 6102 4788 6120
rect 4770 6120 4788 6138
rect 4770 6138 4788 6156
rect 4770 6156 4788 6174
rect 4770 6174 4788 6192
rect 4770 6192 4788 6210
rect 4770 6210 4788 6228
rect 4770 6228 4788 6246
rect 4770 6246 4788 6264
rect 4770 6264 4788 6282
rect 4770 6282 4788 6300
rect 4770 6300 4788 6318
rect 4770 6318 4788 6336
rect 4770 6336 4788 6354
rect 4770 6354 4788 6372
rect 4770 6372 4788 6390
rect 4770 6390 4788 6408
rect 4770 6408 4788 6426
rect 4770 6426 4788 6444
rect 4770 6444 4788 6462
rect 4770 6462 4788 6480
rect 4770 6480 4788 6498
rect 4770 6498 4788 6516
rect 4770 6516 4788 6534
rect 4770 6534 4788 6552
rect 4770 6552 4788 6570
rect 4770 6570 4788 6588
rect 4770 6588 4788 6606
rect 4770 6606 4788 6624
rect 4770 6624 4788 6642
rect 4770 6642 4788 6660
rect 4770 6660 4788 6678
rect 4770 6678 4788 6696
rect 4770 6696 4788 6714
rect 4770 6714 4788 6732
rect 4770 6732 4788 6750
rect 4770 6750 4788 6768
rect 4770 6768 4788 6786
rect 4770 6786 4788 6804
rect 4770 6804 4788 6822
rect 4770 6822 4788 6840
rect 4770 6840 4788 6858
rect 4770 6858 4788 6876
rect 4770 6876 4788 6894
rect 4770 6894 4788 6912
rect 4770 6912 4788 6930
rect 4770 6930 4788 6948
rect 4770 6948 4788 6966
rect 4770 6966 4788 6984
rect 4770 6984 4788 7002
rect 4770 7002 4788 7020
rect 4770 7020 4788 7038
rect 4770 7038 4788 7056
rect 4770 7056 4788 7074
rect 4770 7074 4788 7092
rect 4770 7092 4788 7110
rect 4770 7110 4788 7128
rect 4770 7128 4788 7146
rect 4770 7146 4788 7164
rect 4770 7164 4788 7182
rect 4770 7182 4788 7200
rect 4770 7200 4788 7218
rect 4770 7218 4788 7236
rect 4770 7236 4788 7254
rect 4770 7254 4788 7272
rect 4770 7272 4788 7290
rect 4770 7290 4788 7308
rect 4770 7308 4788 7326
rect 4770 7326 4788 7344
rect 4770 7344 4788 7362
rect 4770 7362 4788 7380
rect 4770 7380 4788 7398
rect 4770 7398 4788 7416
rect 4770 7416 4788 7434
rect 4770 7434 4788 7452
rect 4770 7452 4788 7470
rect 4770 7470 4788 7488
rect 4788 180 4806 198
rect 4788 198 4806 216
rect 4788 216 4806 234
rect 4788 234 4806 252
rect 4788 252 4806 270
rect 4788 270 4806 288
rect 4788 288 4806 306
rect 4788 306 4806 324
rect 4788 324 4806 342
rect 4788 342 4806 360
rect 4788 360 4806 378
rect 4788 378 4806 396
rect 4788 396 4806 414
rect 4788 414 4806 432
rect 4788 432 4806 450
rect 4788 450 4806 468
rect 4788 468 4806 486
rect 4788 486 4806 504
rect 4788 504 4806 522
rect 4788 522 4806 540
rect 4788 540 4806 558
rect 4788 558 4806 576
rect 4788 576 4806 594
rect 4788 594 4806 612
rect 4788 612 4806 630
rect 4788 630 4806 648
rect 4788 648 4806 666
rect 4788 666 4806 684
rect 4788 684 4806 702
rect 4788 702 4806 720
rect 4788 720 4806 738
rect 4788 738 4806 756
rect 4788 864 4806 882
rect 4788 882 4806 900
rect 4788 900 4806 918
rect 4788 918 4806 936
rect 4788 936 4806 954
rect 4788 954 4806 972
rect 4788 972 4806 990
rect 4788 990 4806 1008
rect 4788 1008 4806 1026
rect 4788 1026 4806 1044
rect 4788 1044 4806 1062
rect 4788 1062 4806 1080
rect 4788 1080 4806 1098
rect 4788 1098 4806 1116
rect 4788 1116 4806 1134
rect 4788 1134 4806 1152
rect 4788 1152 4806 1170
rect 4788 1170 4806 1188
rect 4788 1188 4806 1206
rect 4788 1206 4806 1224
rect 4788 1224 4806 1242
rect 4788 1242 4806 1260
rect 4788 1260 4806 1278
rect 4788 1278 4806 1296
rect 4788 1296 4806 1314
rect 4788 1314 4806 1332
rect 4788 1332 4806 1350
rect 4788 1350 4806 1368
rect 4788 1368 4806 1386
rect 4788 1386 4806 1404
rect 4788 1404 4806 1422
rect 4788 1422 4806 1440
rect 4788 1440 4806 1458
rect 4788 1458 4806 1476
rect 4788 1476 4806 1494
rect 4788 1494 4806 1512
rect 4788 1512 4806 1530
rect 4788 1530 4806 1548
rect 4788 1548 4806 1566
rect 4788 1566 4806 1584
rect 4788 1584 4806 1602
rect 4788 1602 4806 1620
rect 4788 1620 4806 1638
rect 4788 1638 4806 1656
rect 4788 1656 4806 1674
rect 4788 1674 4806 1692
rect 4788 1692 4806 1710
rect 4788 1710 4806 1728
rect 4788 1728 4806 1746
rect 4788 1746 4806 1764
rect 4788 1764 4806 1782
rect 4788 1782 4806 1800
rect 4788 1800 4806 1818
rect 4788 1818 4806 1836
rect 4788 1836 4806 1854
rect 4788 1854 4806 1872
rect 4788 1872 4806 1890
rect 4788 1890 4806 1908
rect 4788 1908 4806 1926
rect 4788 1926 4806 1944
rect 4788 1944 4806 1962
rect 4788 1962 4806 1980
rect 4788 1980 4806 1998
rect 4788 1998 4806 2016
rect 4788 2016 4806 2034
rect 4788 2034 4806 2052
rect 4788 2052 4806 2070
rect 4788 2070 4806 2088
rect 4788 2322 4806 2340
rect 4788 2340 4806 2358
rect 4788 2358 4806 2376
rect 4788 2376 4806 2394
rect 4788 2394 4806 2412
rect 4788 2412 4806 2430
rect 4788 2430 4806 2448
rect 4788 2448 4806 2466
rect 4788 2466 4806 2484
rect 4788 2484 4806 2502
rect 4788 2502 4806 2520
rect 4788 2520 4806 2538
rect 4788 2538 4806 2556
rect 4788 2556 4806 2574
rect 4788 2574 4806 2592
rect 4788 2592 4806 2610
rect 4788 2610 4806 2628
rect 4788 2628 4806 2646
rect 4788 2646 4806 2664
rect 4788 2664 4806 2682
rect 4788 2682 4806 2700
rect 4788 2700 4806 2718
rect 4788 2718 4806 2736
rect 4788 2736 4806 2754
rect 4788 2754 4806 2772
rect 4788 2772 4806 2790
rect 4788 2790 4806 2808
rect 4788 2808 4806 2826
rect 4788 2826 4806 2844
rect 4788 2844 4806 2862
rect 4788 2862 4806 2880
rect 4788 2880 4806 2898
rect 4788 2898 4806 2916
rect 4788 2916 4806 2934
rect 4788 2934 4806 2952
rect 4788 2952 4806 2970
rect 4788 2970 4806 2988
rect 4788 2988 4806 3006
rect 4788 3006 4806 3024
rect 4788 3024 4806 3042
rect 4788 3042 4806 3060
rect 4788 3060 4806 3078
rect 4788 3078 4806 3096
rect 4788 3096 4806 3114
rect 4788 3114 4806 3132
rect 4788 3132 4806 3150
rect 4788 3150 4806 3168
rect 4788 3168 4806 3186
rect 4788 3186 4806 3204
rect 4788 3204 4806 3222
rect 4788 3222 4806 3240
rect 4788 3240 4806 3258
rect 4788 3258 4806 3276
rect 4788 3276 4806 3294
rect 4788 3294 4806 3312
rect 4788 3312 4806 3330
rect 4788 3330 4806 3348
rect 4788 3348 4806 3366
rect 4788 3366 4806 3384
rect 4788 3384 4806 3402
rect 4788 3402 4806 3420
rect 4788 3420 4806 3438
rect 4788 3438 4806 3456
rect 4788 3456 4806 3474
rect 4788 3474 4806 3492
rect 4788 3492 4806 3510
rect 4788 3510 4806 3528
rect 4788 3528 4806 3546
rect 4788 3546 4806 3564
rect 4788 3564 4806 3582
rect 4788 3582 4806 3600
rect 4788 3600 4806 3618
rect 4788 3618 4806 3636
rect 4788 3636 4806 3654
rect 4788 3654 4806 3672
rect 4788 3672 4806 3690
rect 4788 3690 4806 3708
rect 4788 3708 4806 3726
rect 4788 3726 4806 3744
rect 4788 3744 4806 3762
rect 4788 3762 4806 3780
rect 4788 3780 4806 3798
rect 4788 3798 4806 3816
rect 4788 3816 4806 3834
rect 4788 3834 4806 3852
rect 4788 3852 4806 3870
rect 4788 3870 4806 3888
rect 4788 3888 4806 3906
rect 4788 3906 4806 3924
rect 4788 3924 4806 3942
rect 4788 3942 4806 3960
rect 4788 3960 4806 3978
rect 4788 3978 4806 3996
rect 4788 3996 4806 4014
rect 4788 4014 4806 4032
rect 4788 4032 4806 4050
rect 4788 4050 4806 4068
rect 4788 4068 4806 4086
rect 4788 4086 4806 4104
rect 4788 4104 4806 4122
rect 4788 4122 4806 4140
rect 4788 4356 4806 4374
rect 4788 4374 4806 4392
rect 4788 4392 4806 4410
rect 4788 4410 4806 4428
rect 4788 4428 4806 4446
rect 4788 4446 4806 4464
rect 4788 4464 4806 4482
rect 4788 4482 4806 4500
rect 4788 4500 4806 4518
rect 4788 4518 4806 4536
rect 4788 4536 4806 4554
rect 4788 4554 4806 4572
rect 4788 4572 4806 4590
rect 4788 4590 4806 4608
rect 4788 4608 4806 4626
rect 4788 4626 4806 4644
rect 4788 4644 4806 4662
rect 4788 4662 4806 4680
rect 4788 4680 4806 4698
rect 4788 4698 4806 4716
rect 4788 4716 4806 4734
rect 4788 4734 4806 4752
rect 4788 4752 4806 4770
rect 4788 4770 4806 4788
rect 4788 4788 4806 4806
rect 4788 4806 4806 4824
rect 4788 4824 4806 4842
rect 4788 4842 4806 4860
rect 4788 4860 4806 4878
rect 4788 4878 4806 4896
rect 4788 4896 4806 4914
rect 4788 4914 4806 4932
rect 4788 4932 4806 4950
rect 4788 4950 4806 4968
rect 4788 4968 4806 4986
rect 4788 4986 4806 5004
rect 4788 5004 4806 5022
rect 4788 5022 4806 5040
rect 4788 5040 4806 5058
rect 4788 5058 4806 5076
rect 4788 5076 4806 5094
rect 4788 5094 4806 5112
rect 4788 5112 4806 5130
rect 4788 5130 4806 5148
rect 4788 5148 4806 5166
rect 4788 5166 4806 5184
rect 4788 5184 4806 5202
rect 4788 5202 4806 5220
rect 4788 5220 4806 5238
rect 4788 5238 4806 5256
rect 4788 5256 4806 5274
rect 4788 5274 4806 5292
rect 4788 5292 4806 5310
rect 4788 5310 4806 5328
rect 4788 5328 4806 5346
rect 4788 5346 4806 5364
rect 4788 5364 4806 5382
rect 4788 5382 4806 5400
rect 4788 5400 4806 5418
rect 4788 5418 4806 5436
rect 4788 5436 4806 5454
rect 4788 5454 4806 5472
rect 4788 5472 4806 5490
rect 4788 5490 4806 5508
rect 4788 5508 4806 5526
rect 4788 5526 4806 5544
rect 4788 5544 4806 5562
rect 4788 5562 4806 5580
rect 4788 5580 4806 5598
rect 4788 5598 4806 5616
rect 4788 5616 4806 5634
rect 4788 5634 4806 5652
rect 4788 5652 4806 5670
rect 4788 5670 4806 5688
rect 4788 5688 4806 5706
rect 4788 5706 4806 5724
rect 4788 5724 4806 5742
rect 4788 5742 4806 5760
rect 4788 5760 4806 5778
rect 4788 5778 4806 5796
rect 4788 5796 4806 5814
rect 4788 5814 4806 5832
rect 4788 5832 4806 5850
rect 4788 5850 4806 5868
rect 4788 5868 4806 5886
rect 4788 5886 4806 5904
rect 4788 5904 4806 5922
rect 4788 5922 4806 5940
rect 4788 5940 4806 5958
rect 4788 5958 4806 5976
rect 4788 5976 4806 5994
rect 4788 5994 4806 6012
rect 4788 6012 4806 6030
rect 4788 6030 4806 6048
rect 4788 6048 4806 6066
rect 4788 6066 4806 6084
rect 4788 6084 4806 6102
rect 4788 6102 4806 6120
rect 4788 6120 4806 6138
rect 4788 6138 4806 6156
rect 4788 6156 4806 6174
rect 4788 6174 4806 6192
rect 4788 6192 4806 6210
rect 4788 6210 4806 6228
rect 4788 6228 4806 6246
rect 4788 6246 4806 6264
rect 4788 6264 4806 6282
rect 4788 6282 4806 6300
rect 4788 6300 4806 6318
rect 4788 6318 4806 6336
rect 4788 6336 4806 6354
rect 4788 6354 4806 6372
rect 4788 6372 4806 6390
rect 4788 6390 4806 6408
rect 4788 6408 4806 6426
rect 4788 6426 4806 6444
rect 4788 6444 4806 6462
rect 4788 6462 4806 6480
rect 4788 6480 4806 6498
rect 4788 6498 4806 6516
rect 4788 6516 4806 6534
rect 4788 6534 4806 6552
rect 4788 6552 4806 6570
rect 4788 6570 4806 6588
rect 4788 6588 4806 6606
rect 4788 6606 4806 6624
rect 4788 6624 4806 6642
rect 4788 6642 4806 6660
rect 4788 6660 4806 6678
rect 4788 6678 4806 6696
rect 4788 6696 4806 6714
rect 4788 6714 4806 6732
rect 4788 6732 4806 6750
rect 4788 6750 4806 6768
rect 4788 6768 4806 6786
rect 4788 6786 4806 6804
rect 4788 6804 4806 6822
rect 4788 6822 4806 6840
rect 4788 6840 4806 6858
rect 4788 6858 4806 6876
rect 4788 6876 4806 6894
rect 4788 6894 4806 6912
rect 4788 6912 4806 6930
rect 4788 6930 4806 6948
rect 4788 6948 4806 6966
rect 4788 6966 4806 6984
rect 4788 6984 4806 7002
rect 4788 7002 4806 7020
rect 4788 7020 4806 7038
rect 4788 7038 4806 7056
rect 4788 7056 4806 7074
rect 4788 7074 4806 7092
rect 4788 7092 4806 7110
rect 4788 7110 4806 7128
rect 4788 7128 4806 7146
rect 4788 7146 4806 7164
rect 4788 7164 4806 7182
rect 4788 7182 4806 7200
rect 4788 7200 4806 7218
rect 4788 7218 4806 7236
rect 4788 7236 4806 7254
rect 4788 7254 4806 7272
rect 4788 7272 4806 7290
rect 4788 7290 4806 7308
rect 4788 7308 4806 7326
rect 4788 7326 4806 7344
rect 4788 7344 4806 7362
rect 4788 7362 4806 7380
rect 4788 7380 4806 7398
rect 4788 7398 4806 7416
rect 4788 7416 4806 7434
rect 4788 7434 4806 7452
rect 4788 7452 4806 7470
rect 4788 7470 4806 7488
rect 4788 7488 4806 7506
rect 4788 7506 4806 7524
rect 4806 198 4824 216
rect 4806 216 4824 234
rect 4806 234 4824 252
rect 4806 252 4824 270
rect 4806 270 4824 288
rect 4806 288 4824 306
rect 4806 306 4824 324
rect 4806 324 4824 342
rect 4806 342 4824 360
rect 4806 360 4824 378
rect 4806 378 4824 396
rect 4806 396 4824 414
rect 4806 414 4824 432
rect 4806 432 4824 450
rect 4806 450 4824 468
rect 4806 468 4824 486
rect 4806 486 4824 504
rect 4806 504 4824 522
rect 4806 522 4824 540
rect 4806 540 4824 558
rect 4806 558 4824 576
rect 4806 576 4824 594
rect 4806 594 4824 612
rect 4806 612 4824 630
rect 4806 630 4824 648
rect 4806 648 4824 666
rect 4806 666 4824 684
rect 4806 684 4824 702
rect 4806 702 4824 720
rect 4806 720 4824 738
rect 4806 738 4824 756
rect 4806 864 4824 882
rect 4806 882 4824 900
rect 4806 900 4824 918
rect 4806 918 4824 936
rect 4806 936 4824 954
rect 4806 954 4824 972
rect 4806 972 4824 990
rect 4806 990 4824 1008
rect 4806 1008 4824 1026
rect 4806 1026 4824 1044
rect 4806 1044 4824 1062
rect 4806 1062 4824 1080
rect 4806 1080 4824 1098
rect 4806 1098 4824 1116
rect 4806 1116 4824 1134
rect 4806 1134 4824 1152
rect 4806 1152 4824 1170
rect 4806 1170 4824 1188
rect 4806 1188 4824 1206
rect 4806 1206 4824 1224
rect 4806 1224 4824 1242
rect 4806 1242 4824 1260
rect 4806 1260 4824 1278
rect 4806 1278 4824 1296
rect 4806 1296 4824 1314
rect 4806 1314 4824 1332
rect 4806 1332 4824 1350
rect 4806 1350 4824 1368
rect 4806 1368 4824 1386
rect 4806 1386 4824 1404
rect 4806 1404 4824 1422
rect 4806 1422 4824 1440
rect 4806 1440 4824 1458
rect 4806 1458 4824 1476
rect 4806 1476 4824 1494
rect 4806 1494 4824 1512
rect 4806 1512 4824 1530
rect 4806 1530 4824 1548
rect 4806 1548 4824 1566
rect 4806 1566 4824 1584
rect 4806 1584 4824 1602
rect 4806 1602 4824 1620
rect 4806 1620 4824 1638
rect 4806 1638 4824 1656
rect 4806 1656 4824 1674
rect 4806 1674 4824 1692
rect 4806 1692 4824 1710
rect 4806 1710 4824 1728
rect 4806 1728 4824 1746
rect 4806 1746 4824 1764
rect 4806 1764 4824 1782
rect 4806 1782 4824 1800
rect 4806 1800 4824 1818
rect 4806 1818 4824 1836
rect 4806 1836 4824 1854
rect 4806 1854 4824 1872
rect 4806 1872 4824 1890
rect 4806 1890 4824 1908
rect 4806 1908 4824 1926
rect 4806 1926 4824 1944
rect 4806 1944 4824 1962
rect 4806 1962 4824 1980
rect 4806 1980 4824 1998
rect 4806 1998 4824 2016
rect 4806 2016 4824 2034
rect 4806 2034 4824 2052
rect 4806 2052 4824 2070
rect 4806 2070 4824 2088
rect 4806 2088 4824 2106
rect 4806 2322 4824 2340
rect 4806 2340 4824 2358
rect 4806 2358 4824 2376
rect 4806 2376 4824 2394
rect 4806 2394 4824 2412
rect 4806 2412 4824 2430
rect 4806 2430 4824 2448
rect 4806 2448 4824 2466
rect 4806 2466 4824 2484
rect 4806 2484 4824 2502
rect 4806 2502 4824 2520
rect 4806 2520 4824 2538
rect 4806 2538 4824 2556
rect 4806 2556 4824 2574
rect 4806 2574 4824 2592
rect 4806 2592 4824 2610
rect 4806 2610 4824 2628
rect 4806 2628 4824 2646
rect 4806 2646 4824 2664
rect 4806 2664 4824 2682
rect 4806 2682 4824 2700
rect 4806 2700 4824 2718
rect 4806 2718 4824 2736
rect 4806 2736 4824 2754
rect 4806 2754 4824 2772
rect 4806 2772 4824 2790
rect 4806 2790 4824 2808
rect 4806 2808 4824 2826
rect 4806 2826 4824 2844
rect 4806 2844 4824 2862
rect 4806 2862 4824 2880
rect 4806 2880 4824 2898
rect 4806 2898 4824 2916
rect 4806 2916 4824 2934
rect 4806 2934 4824 2952
rect 4806 2952 4824 2970
rect 4806 2970 4824 2988
rect 4806 2988 4824 3006
rect 4806 3006 4824 3024
rect 4806 3024 4824 3042
rect 4806 3042 4824 3060
rect 4806 3060 4824 3078
rect 4806 3078 4824 3096
rect 4806 3096 4824 3114
rect 4806 3114 4824 3132
rect 4806 3132 4824 3150
rect 4806 3150 4824 3168
rect 4806 3168 4824 3186
rect 4806 3186 4824 3204
rect 4806 3204 4824 3222
rect 4806 3222 4824 3240
rect 4806 3240 4824 3258
rect 4806 3258 4824 3276
rect 4806 3276 4824 3294
rect 4806 3294 4824 3312
rect 4806 3312 4824 3330
rect 4806 3330 4824 3348
rect 4806 3348 4824 3366
rect 4806 3366 4824 3384
rect 4806 3384 4824 3402
rect 4806 3402 4824 3420
rect 4806 3420 4824 3438
rect 4806 3438 4824 3456
rect 4806 3456 4824 3474
rect 4806 3474 4824 3492
rect 4806 3492 4824 3510
rect 4806 3510 4824 3528
rect 4806 3528 4824 3546
rect 4806 3546 4824 3564
rect 4806 3564 4824 3582
rect 4806 3582 4824 3600
rect 4806 3600 4824 3618
rect 4806 3618 4824 3636
rect 4806 3636 4824 3654
rect 4806 3654 4824 3672
rect 4806 3672 4824 3690
rect 4806 3690 4824 3708
rect 4806 3708 4824 3726
rect 4806 3726 4824 3744
rect 4806 3744 4824 3762
rect 4806 3762 4824 3780
rect 4806 3780 4824 3798
rect 4806 3798 4824 3816
rect 4806 3816 4824 3834
rect 4806 3834 4824 3852
rect 4806 3852 4824 3870
rect 4806 3870 4824 3888
rect 4806 3888 4824 3906
rect 4806 3906 4824 3924
rect 4806 3924 4824 3942
rect 4806 3942 4824 3960
rect 4806 3960 4824 3978
rect 4806 3978 4824 3996
rect 4806 3996 4824 4014
rect 4806 4014 4824 4032
rect 4806 4032 4824 4050
rect 4806 4050 4824 4068
rect 4806 4068 4824 4086
rect 4806 4086 4824 4104
rect 4806 4104 4824 4122
rect 4806 4122 4824 4140
rect 4806 4140 4824 4158
rect 4806 4158 4824 4176
rect 4806 4374 4824 4392
rect 4806 4392 4824 4410
rect 4806 4410 4824 4428
rect 4806 4428 4824 4446
rect 4806 4446 4824 4464
rect 4806 4464 4824 4482
rect 4806 4482 4824 4500
rect 4806 4500 4824 4518
rect 4806 4518 4824 4536
rect 4806 4536 4824 4554
rect 4806 4554 4824 4572
rect 4806 4572 4824 4590
rect 4806 4590 4824 4608
rect 4806 4608 4824 4626
rect 4806 4626 4824 4644
rect 4806 4644 4824 4662
rect 4806 4662 4824 4680
rect 4806 4680 4824 4698
rect 4806 4698 4824 4716
rect 4806 4716 4824 4734
rect 4806 4734 4824 4752
rect 4806 4752 4824 4770
rect 4806 4770 4824 4788
rect 4806 4788 4824 4806
rect 4806 4806 4824 4824
rect 4806 4824 4824 4842
rect 4806 4842 4824 4860
rect 4806 4860 4824 4878
rect 4806 4878 4824 4896
rect 4806 4896 4824 4914
rect 4806 4914 4824 4932
rect 4806 4932 4824 4950
rect 4806 4950 4824 4968
rect 4806 4968 4824 4986
rect 4806 4986 4824 5004
rect 4806 5004 4824 5022
rect 4806 5022 4824 5040
rect 4806 5040 4824 5058
rect 4806 5058 4824 5076
rect 4806 5076 4824 5094
rect 4806 5094 4824 5112
rect 4806 5112 4824 5130
rect 4806 5130 4824 5148
rect 4806 5148 4824 5166
rect 4806 5166 4824 5184
rect 4806 5184 4824 5202
rect 4806 5202 4824 5220
rect 4806 5220 4824 5238
rect 4806 5238 4824 5256
rect 4806 5256 4824 5274
rect 4806 5274 4824 5292
rect 4806 5292 4824 5310
rect 4806 5310 4824 5328
rect 4806 5328 4824 5346
rect 4806 5346 4824 5364
rect 4806 5364 4824 5382
rect 4806 5382 4824 5400
rect 4806 5400 4824 5418
rect 4806 5418 4824 5436
rect 4806 5436 4824 5454
rect 4806 5454 4824 5472
rect 4806 5472 4824 5490
rect 4806 5490 4824 5508
rect 4806 5508 4824 5526
rect 4806 5526 4824 5544
rect 4806 5544 4824 5562
rect 4806 5562 4824 5580
rect 4806 5580 4824 5598
rect 4806 5598 4824 5616
rect 4806 5616 4824 5634
rect 4806 5634 4824 5652
rect 4806 5652 4824 5670
rect 4806 5670 4824 5688
rect 4806 5688 4824 5706
rect 4806 5706 4824 5724
rect 4806 5724 4824 5742
rect 4806 5742 4824 5760
rect 4806 5760 4824 5778
rect 4806 5778 4824 5796
rect 4806 5796 4824 5814
rect 4806 5814 4824 5832
rect 4806 5832 4824 5850
rect 4806 5850 4824 5868
rect 4806 5868 4824 5886
rect 4806 5886 4824 5904
rect 4806 5904 4824 5922
rect 4806 5922 4824 5940
rect 4806 5940 4824 5958
rect 4806 5958 4824 5976
rect 4806 5976 4824 5994
rect 4806 5994 4824 6012
rect 4806 6012 4824 6030
rect 4806 6030 4824 6048
rect 4806 6048 4824 6066
rect 4806 6066 4824 6084
rect 4806 6084 4824 6102
rect 4806 6102 4824 6120
rect 4806 6120 4824 6138
rect 4806 6138 4824 6156
rect 4806 6156 4824 6174
rect 4806 6174 4824 6192
rect 4806 6192 4824 6210
rect 4806 6210 4824 6228
rect 4806 6228 4824 6246
rect 4806 6246 4824 6264
rect 4806 6264 4824 6282
rect 4806 6282 4824 6300
rect 4806 6300 4824 6318
rect 4806 6318 4824 6336
rect 4806 6336 4824 6354
rect 4806 6354 4824 6372
rect 4806 6372 4824 6390
rect 4806 6390 4824 6408
rect 4806 6408 4824 6426
rect 4806 6426 4824 6444
rect 4806 6444 4824 6462
rect 4806 6462 4824 6480
rect 4806 6480 4824 6498
rect 4806 6498 4824 6516
rect 4806 6516 4824 6534
rect 4806 6534 4824 6552
rect 4806 6552 4824 6570
rect 4806 6570 4824 6588
rect 4806 6588 4824 6606
rect 4806 6606 4824 6624
rect 4806 6624 4824 6642
rect 4806 6642 4824 6660
rect 4806 6660 4824 6678
rect 4806 6678 4824 6696
rect 4806 6696 4824 6714
rect 4806 6714 4824 6732
rect 4806 6732 4824 6750
rect 4806 6750 4824 6768
rect 4806 6768 4824 6786
rect 4806 6786 4824 6804
rect 4806 6804 4824 6822
rect 4806 6822 4824 6840
rect 4806 6840 4824 6858
rect 4806 6858 4824 6876
rect 4806 6876 4824 6894
rect 4806 6894 4824 6912
rect 4806 6912 4824 6930
rect 4806 6930 4824 6948
rect 4806 6948 4824 6966
rect 4806 6966 4824 6984
rect 4806 6984 4824 7002
rect 4806 7002 4824 7020
rect 4806 7020 4824 7038
rect 4806 7038 4824 7056
rect 4806 7056 4824 7074
rect 4806 7074 4824 7092
rect 4806 7092 4824 7110
rect 4806 7110 4824 7128
rect 4806 7128 4824 7146
rect 4806 7146 4824 7164
rect 4806 7164 4824 7182
rect 4806 7182 4824 7200
rect 4806 7200 4824 7218
rect 4806 7218 4824 7236
rect 4806 7236 4824 7254
rect 4806 7254 4824 7272
rect 4806 7272 4824 7290
rect 4806 7290 4824 7308
rect 4806 7308 4824 7326
rect 4806 7326 4824 7344
rect 4806 7344 4824 7362
rect 4806 7362 4824 7380
rect 4806 7380 4824 7398
rect 4806 7398 4824 7416
rect 4806 7416 4824 7434
rect 4806 7434 4824 7452
rect 4806 7452 4824 7470
rect 4806 7470 4824 7488
rect 4806 7488 4824 7506
rect 4806 7506 4824 7524
rect 4806 7524 4824 7542
rect 4824 198 4842 216
rect 4824 216 4842 234
rect 4824 234 4842 252
rect 4824 252 4842 270
rect 4824 270 4842 288
rect 4824 288 4842 306
rect 4824 306 4842 324
rect 4824 324 4842 342
rect 4824 342 4842 360
rect 4824 360 4842 378
rect 4824 378 4842 396
rect 4824 396 4842 414
rect 4824 414 4842 432
rect 4824 432 4842 450
rect 4824 450 4842 468
rect 4824 468 4842 486
rect 4824 486 4842 504
rect 4824 504 4842 522
rect 4824 522 4842 540
rect 4824 540 4842 558
rect 4824 558 4842 576
rect 4824 576 4842 594
rect 4824 594 4842 612
rect 4824 612 4842 630
rect 4824 630 4842 648
rect 4824 648 4842 666
rect 4824 666 4842 684
rect 4824 684 4842 702
rect 4824 702 4842 720
rect 4824 720 4842 738
rect 4824 738 4842 756
rect 4824 864 4842 882
rect 4824 882 4842 900
rect 4824 900 4842 918
rect 4824 918 4842 936
rect 4824 936 4842 954
rect 4824 954 4842 972
rect 4824 972 4842 990
rect 4824 990 4842 1008
rect 4824 1008 4842 1026
rect 4824 1026 4842 1044
rect 4824 1044 4842 1062
rect 4824 1062 4842 1080
rect 4824 1080 4842 1098
rect 4824 1098 4842 1116
rect 4824 1116 4842 1134
rect 4824 1134 4842 1152
rect 4824 1152 4842 1170
rect 4824 1170 4842 1188
rect 4824 1188 4842 1206
rect 4824 1206 4842 1224
rect 4824 1224 4842 1242
rect 4824 1242 4842 1260
rect 4824 1260 4842 1278
rect 4824 1278 4842 1296
rect 4824 1296 4842 1314
rect 4824 1314 4842 1332
rect 4824 1332 4842 1350
rect 4824 1350 4842 1368
rect 4824 1368 4842 1386
rect 4824 1386 4842 1404
rect 4824 1404 4842 1422
rect 4824 1422 4842 1440
rect 4824 1440 4842 1458
rect 4824 1458 4842 1476
rect 4824 1476 4842 1494
rect 4824 1494 4842 1512
rect 4824 1512 4842 1530
rect 4824 1530 4842 1548
rect 4824 1548 4842 1566
rect 4824 1566 4842 1584
rect 4824 1584 4842 1602
rect 4824 1602 4842 1620
rect 4824 1620 4842 1638
rect 4824 1638 4842 1656
rect 4824 1656 4842 1674
rect 4824 1674 4842 1692
rect 4824 1692 4842 1710
rect 4824 1710 4842 1728
rect 4824 1728 4842 1746
rect 4824 1746 4842 1764
rect 4824 1764 4842 1782
rect 4824 1782 4842 1800
rect 4824 1800 4842 1818
rect 4824 1818 4842 1836
rect 4824 1836 4842 1854
rect 4824 1854 4842 1872
rect 4824 1872 4842 1890
rect 4824 1890 4842 1908
rect 4824 1908 4842 1926
rect 4824 1926 4842 1944
rect 4824 1944 4842 1962
rect 4824 1962 4842 1980
rect 4824 1980 4842 1998
rect 4824 1998 4842 2016
rect 4824 2016 4842 2034
rect 4824 2034 4842 2052
rect 4824 2052 4842 2070
rect 4824 2070 4842 2088
rect 4824 2088 4842 2106
rect 4824 2106 4842 2124
rect 4824 2340 4842 2358
rect 4824 2358 4842 2376
rect 4824 2376 4842 2394
rect 4824 2394 4842 2412
rect 4824 2412 4842 2430
rect 4824 2430 4842 2448
rect 4824 2448 4842 2466
rect 4824 2466 4842 2484
rect 4824 2484 4842 2502
rect 4824 2502 4842 2520
rect 4824 2520 4842 2538
rect 4824 2538 4842 2556
rect 4824 2556 4842 2574
rect 4824 2574 4842 2592
rect 4824 2592 4842 2610
rect 4824 2610 4842 2628
rect 4824 2628 4842 2646
rect 4824 2646 4842 2664
rect 4824 2664 4842 2682
rect 4824 2682 4842 2700
rect 4824 2700 4842 2718
rect 4824 2718 4842 2736
rect 4824 2736 4842 2754
rect 4824 2754 4842 2772
rect 4824 2772 4842 2790
rect 4824 2790 4842 2808
rect 4824 2808 4842 2826
rect 4824 2826 4842 2844
rect 4824 2844 4842 2862
rect 4824 2862 4842 2880
rect 4824 2880 4842 2898
rect 4824 2898 4842 2916
rect 4824 2916 4842 2934
rect 4824 2934 4842 2952
rect 4824 2952 4842 2970
rect 4824 2970 4842 2988
rect 4824 2988 4842 3006
rect 4824 3006 4842 3024
rect 4824 3024 4842 3042
rect 4824 3042 4842 3060
rect 4824 3060 4842 3078
rect 4824 3078 4842 3096
rect 4824 3096 4842 3114
rect 4824 3114 4842 3132
rect 4824 3132 4842 3150
rect 4824 3150 4842 3168
rect 4824 3168 4842 3186
rect 4824 3186 4842 3204
rect 4824 3204 4842 3222
rect 4824 3222 4842 3240
rect 4824 3240 4842 3258
rect 4824 3258 4842 3276
rect 4824 3276 4842 3294
rect 4824 3294 4842 3312
rect 4824 3312 4842 3330
rect 4824 3330 4842 3348
rect 4824 3348 4842 3366
rect 4824 3366 4842 3384
rect 4824 3384 4842 3402
rect 4824 3402 4842 3420
rect 4824 3420 4842 3438
rect 4824 3438 4842 3456
rect 4824 3456 4842 3474
rect 4824 3474 4842 3492
rect 4824 3492 4842 3510
rect 4824 3510 4842 3528
rect 4824 3528 4842 3546
rect 4824 3546 4842 3564
rect 4824 3564 4842 3582
rect 4824 3582 4842 3600
rect 4824 3600 4842 3618
rect 4824 3618 4842 3636
rect 4824 3636 4842 3654
rect 4824 3654 4842 3672
rect 4824 3672 4842 3690
rect 4824 3690 4842 3708
rect 4824 3708 4842 3726
rect 4824 3726 4842 3744
rect 4824 3744 4842 3762
rect 4824 3762 4842 3780
rect 4824 3780 4842 3798
rect 4824 3798 4842 3816
rect 4824 3816 4842 3834
rect 4824 3834 4842 3852
rect 4824 3852 4842 3870
rect 4824 3870 4842 3888
rect 4824 3888 4842 3906
rect 4824 3906 4842 3924
rect 4824 3924 4842 3942
rect 4824 3942 4842 3960
rect 4824 3960 4842 3978
rect 4824 3978 4842 3996
rect 4824 3996 4842 4014
rect 4824 4014 4842 4032
rect 4824 4032 4842 4050
rect 4824 4050 4842 4068
rect 4824 4068 4842 4086
rect 4824 4086 4842 4104
rect 4824 4104 4842 4122
rect 4824 4122 4842 4140
rect 4824 4140 4842 4158
rect 4824 4158 4842 4176
rect 4824 4176 4842 4194
rect 4824 4392 4842 4410
rect 4824 4410 4842 4428
rect 4824 4428 4842 4446
rect 4824 4446 4842 4464
rect 4824 4464 4842 4482
rect 4824 4482 4842 4500
rect 4824 4500 4842 4518
rect 4824 4518 4842 4536
rect 4824 4536 4842 4554
rect 4824 4554 4842 4572
rect 4824 4572 4842 4590
rect 4824 4590 4842 4608
rect 4824 4608 4842 4626
rect 4824 4626 4842 4644
rect 4824 4644 4842 4662
rect 4824 4662 4842 4680
rect 4824 4680 4842 4698
rect 4824 4698 4842 4716
rect 4824 4716 4842 4734
rect 4824 4734 4842 4752
rect 4824 4752 4842 4770
rect 4824 4770 4842 4788
rect 4824 4788 4842 4806
rect 4824 4806 4842 4824
rect 4824 4824 4842 4842
rect 4824 4842 4842 4860
rect 4824 4860 4842 4878
rect 4824 4878 4842 4896
rect 4824 4896 4842 4914
rect 4824 4914 4842 4932
rect 4824 4932 4842 4950
rect 4824 4950 4842 4968
rect 4824 4968 4842 4986
rect 4824 4986 4842 5004
rect 4824 5004 4842 5022
rect 4824 5022 4842 5040
rect 4824 5040 4842 5058
rect 4824 5058 4842 5076
rect 4824 5076 4842 5094
rect 4824 5094 4842 5112
rect 4824 5112 4842 5130
rect 4824 5130 4842 5148
rect 4824 5148 4842 5166
rect 4824 5166 4842 5184
rect 4824 5184 4842 5202
rect 4824 5202 4842 5220
rect 4824 5220 4842 5238
rect 4824 5238 4842 5256
rect 4824 5256 4842 5274
rect 4824 5274 4842 5292
rect 4824 5292 4842 5310
rect 4824 5310 4842 5328
rect 4824 5328 4842 5346
rect 4824 5346 4842 5364
rect 4824 5364 4842 5382
rect 4824 5382 4842 5400
rect 4824 5400 4842 5418
rect 4824 5418 4842 5436
rect 4824 5436 4842 5454
rect 4824 5454 4842 5472
rect 4824 5472 4842 5490
rect 4824 5490 4842 5508
rect 4824 5508 4842 5526
rect 4824 5526 4842 5544
rect 4824 5544 4842 5562
rect 4824 5562 4842 5580
rect 4824 5580 4842 5598
rect 4824 5598 4842 5616
rect 4824 5616 4842 5634
rect 4824 5634 4842 5652
rect 4824 5652 4842 5670
rect 4824 5670 4842 5688
rect 4824 5688 4842 5706
rect 4824 5706 4842 5724
rect 4824 5724 4842 5742
rect 4824 5742 4842 5760
rect 4824 5760 4842 5778
rect 4824 5778 4842 5796
rect 4824 5796 4842 5814
rect 4824 5814 4842 5832
rect 4824 5832 4842 5850
rect 4824 5850 4842 5868
rect 4824 5868 4842 5886
rect 4824 5886 4842 5904
rect 4824 5904 4842 5922
rect 4824 5922 4842 5940
rect 4824 5940 4842 5958
rect 4824 5958 4842 5976
rect 4824 5976 4842 5994
rect 4824 5994 4842 6012
rect 4824 6012 4842 6030
rect 4824 6030 4842 6048
rect 4824 6048 4842 6066
rect 4824 6066 4842 6084
rect 4824 6084 4842 6102
rect 4824 6102 4842 6120
rect 4824 6120 4842 6138
rect 4824 6138 4842 6156
rect 4824 6156 4842 6174
rect 4824 6174 4842 6192
rect 4824 6192 4842 6210
rect 4824 6210 4842 6228
rect 4824 6228 4842 6246
rect 4824 6246 4842 6264
rect 4824 6264 4842 6282
rect 4824 6282 4842 6300
rect 4824 6300 4842 6318
rect 4824 6318 4842 6336
rect 4824 6336 4842 6354
rect 4824 6354 4842 6372
rect 4824 6372 4842 6390
rect 4824 6390 4842 6408
rect 4824 6408 4842 6426
rect 4824 6426 4842 6444
rect 4824 6444 4842 6462
rect 4824 6462 4842 6480
rect 4824 6480 4842 6498
rect 4824 6498 4842 6516
rect 4824 6516 4842 6534
rect 4824 6534 4842 6552
rect 4824 6552 4842 6570
rect 4824 6570 4842 6588
rect 4824 6588 4842 6606
rect 4824 6606 4842 6624
rect 4824 6624 4842 6642
rect 4824 6642 4842 6660
rect 4824 6660 4842 6678
rect 4824 6678 4842 6696
rect 4824 6696 4842 6714
rect 4824 6714 4842 6732
rect 4824 6732 4842 6750
rect 4824 6750 4842 6768
rect 4824 6768 4842 6786
rect 4824 6786 4842 6804
rect 4824 6804 4842 6822
rect 4824 6822 4842 6840
rect 4824 6840 4842 6858
rect 4824 6858 4842 6876
rect 4824 6876 4842 6894
rect 4824 6894 4842 6912
rect 4824 6912 4842 6930
rect 4824 6930 4842 6948
rect 4824 6948 4842 6966
rect 4824 6966 4842 6984
rect 4824 6984 4842 7002
rect 4824 7002 4842 7020
rect 4824 7020 4842 7038
rect 4824 7038 4842 7056
rect 4824 7056 4842 7074
rect 4824 7074 4842 7092
rect 4824 7092 4842 7110
rect 4824 7110 4842 7128
rect 4824 7128 4842 7146
rect 4824 7146 4842 7164
rect 4824 7164 4842 7182
rect 4824 7182 4842 7200
rect 4824 7200 4842 7218
rect 4824 7218 4842 7236
rect 4824 7236 4842 7254
rect 4824 7254 4842 7272
rect 4824 7272 4842 7290
rect 4824 7290 4842 7308
rect 4824 7308 4842 7326
rect 4824 7326 4842 7344
rect 4824 7344 4842 7362
rect 4824 7362 4842 7380
rect 4824 7380 4842 7398
rect 4824 7398 4842 7416
rect 4824 7416 4842 7434
rect 4824 7434 4842 7452
rect 4824 7452 4842 7470
rect 4824 7470 4842 7488
rect 4824 7488 4842 7506
rect 4824 7506 4842 7524
rect 4824 7524 4842 7542
rect 4824 7542 4842 7560
rect 4824 7560 4842 7578
rect 4842 198 4860 216
rect 4842 216 4860 234
rect 4842 234 4860 252
rect 4842 252 4860 270
rect 4842 270 4860 288
rect 4842 288 4860 306
rect 4842 306 4860 324
rect 4842 324 4860 342
rect 4842 342 4860 360
rect 4842 360 4860 378
rect 4842 378 4860 396
rect 4842 396 4860 414
rect 4842 414 4860 432
rect 4842 432 4860 450
rect 4842 450 4860 468
rect 4842 468 4860 486
rect 4842 486 4860 504
rect 4842 504 4860 522
rect 4842 522 4860 540
rect 4842 540 4860 558
rect 4842 558 4860 576
rect 4842 576 4860 594
rect 4842 594 4860 612
rect 4842 612 4860 630
rect 4842 630 4860 648
rect 4842 648 4860 666
rect 4842 666 4860 684
rect 4842 684 4860 702
rect 4842 702 4860 720
rect 4842 720 4860 738
rect 4842 738 4860 756
rect 4842 864 4860 882
rect 4842 882 4860 900
rect 4842 900 4860 918
rect 4842 918 4860 936
rect 4842 936 4860 954
rect 4842 954 4860 972
rect 4842 972 4860 990
rect 4842 990 4860 1008
rect 4842 1008 4860 1026
rect 4842 1026 4860 1044
rect 4842 1044 4860 1062
rect 4842 1062 4860 1080
rect 4842 1080 4860 1098
rect 4842 1098 4860 1116
rect 4842 1116 4860 1134
rect 4842 1134 4860 1152
rect 4842 1152 4860 1170
rect 4842 1170 4860 1188
rect 4842 1188 4860 1206
rect 4842 1206 4860 1224
rect 4842 1224 4860 1242
rect 4842 1242 4860 1260
rect 4842 1260 4860 1278
rect 4842 1278 4860 1296
rect 4842 1296 4860 1314
rect 4842 1314 4860 1332
rect 4842 1332 4860 1350
rect 4842 1350 4860 1368
rect 4842 1368 4860 1386
rect 4842 1386 4860 1404
rect 4842 1404 4860 1422
rect 4842 1422 4860 1440
rect 4842 1440 4860 1458
rect 4842 1458 4860 1476
rect 4842 1476 4860 1494
rect 4842 1494 4860 1512
rect 4842 1512 4860 1530
rect 4842 1530 4860 1548
rect 4842 1548 4860 1566
rect 4842 1566 4860 1584
rect 4842 1584 4860 1602
rect 4842 1602 4860 1620
rect 4842 1620 4860 1638
rect 4842 1638 4860 1656
rect 4842 1656 4860 1674
rect 4842 1674 4860 1692
rect 4842 1692 4860 1710
rect 4842 1710 4860 1728
rect 4842 1728 4860 1746
rect 4842 1746 4860 1764
rect 4842 1764 4860 1782
rect 4842 1782 4860 1800
rect 4842 1800 4860 1818
rect 4842 1818 4860 1836
rect 4842 1836 4860 1854
rect 4842 1854 4860 1872
rect 4842 1872 4860 1890
rect 4842 1890 4860 1908
rect 4842 1908 4860 1926
rect 4842 1926 4860 1944
rect 4842 1944 4860 1962
rect 4842 1962 4860 1980
rect 4842 1980 4860 1998
rect 4842 1998 4860 2016
rect 4842 2016 4860 2034
rect 4842 2034 4860 2052
rect 4842 2052 4860 2070
rect 4842 2070 4860 2088
rect 4842 2088 4860 2106
rect 4842 2106 4860 2124
rect 4842 2358 4860 2376
rect 4842 2376 4860 2394
rect 4842 2394 4860 2412
rect 4842 2412 4860 2430
rect 4842 2430 4860 2448
rect 4842 2448 4860 2466
rect 4842 2466 4860 2484
rect 4842 2484 4860 2502
rect 4842 2502 4860 2520
rect 4842 2520 4860 2538
rect 4842 2538 4860 2556
rect 4842 2556 4860 2574
rect 4842 2574 4860 2592
rect 4842 2592 4860 2610
rect 4842 2610 4860 2628
rect 4842 2628 4860 2646
rect 4842 2646 4860 2664
rect 4842 2664 4860 2682
rect 4842 2682 4860 2700
rect 4842 2700 4860 2718
rect 4842 2718 4860 2736
rect 4842 2736 4860 2754
rect 4842 2754 4860 2772
rect 4842 2772 4860 2790
rect 4842 2790 4860 2808
rect 4842 2808 4860 2826
rect 4842 2826 4860 2844
rect 4842 2844 4860 2862
rect 4842 2862 4860 2880
rect 4842 2880 4860 2898
rect 4842 2898 4860 2916
rect 4842 2916 4860 2934
rect 4842 2934 4860 2952
rect 4842 2952 4860 2970
rect 4842 2970 4860 2988
rect 4842 2988 4860 3006
rect 4842 3006 4860 3024
rect 4842 3024 4860 3042
rect 4842 3042 4860 3060
rect 4842 3060 4860 3078
rect 4842 3078 4860 3096
rect 4842 3096 4860 3114
rect 4842 3114 4860 3132
rect 4842 3132 4860 3150
rect 4842 3150 4860 3168
rect 4842 3168 4860 3186
rect 4842 3186 4860 3204
rect 4842 3204 4860 3222
rect 4842 3222 4860 3240
rect 4842 3240 4860 3258
rect 4842 3258 4860 3276
rect 4842 3276 4860 3294
rect 4842 3294 4860 3312
rect 4842 3312 4860 3330
rect 4842 3330 4860 3348
rect 4842 3348 4860 3366
rect 4842 3366 4860 3384
rect 4842 3384 4860 3402
rect 4842 3402 4860 3420
rect 4842 3420 4860 3438
rect 4842 3438 4860 3456
rect 4842 3456 4860 3474
rect 4842 3474 4860 3492
rect 4842 3492 4860 3510
rect 4842 3510 4860 3528
rect 4842 3528 4860 3546
rect 4842 3546 4860 3564
rect 4842 3564 4860 3582
rect 4842 3582 4860 3600
rect 4842 3600 4860 3618
rect 4842 3618 4860 3636
rect 4842 3636 4860 3654
rect 4842 3654 4860 3672
rect 4842 3672 4860 3690
rect 4842 3690 4860 3708
rect 4842 3708 4860 3726
rect 4842 3726 4860 3744
rect 4842 3744 4860 3762
rect 4842 3762 4860 3780
rect 4842 3780 4860 3798
rect 4842 3798 4860 3816
rect 4842 3816 4860 3834
rect 4842 3834 4860 3852
rect 4842 3852 4860 3870
rect 4842 3870 4860 3888
rect 4842 3888 4860 3906
rect 4842 3906 4860 3924
rect 4842 3924 4860 3942
rect 4842 3942 4860 3960
rect 4842 3960 4860 3978
rect 4842 3978 4860 3996
rect 4842 3996 4860 4014
rect 4842 4014 4860 4032
rect 4842 4032 4860 4050
rect 4842 4050 4860 4068
rect 4842 4068 4860 4086
rect 4842 4086 4860 4104
rect 4842 4104 4860 4122
rect 4842 4122 4860 4140
rect 4842 4140 4860 4158
rect 4842 4158 4860 4176
rect 4842 4176 4860 4194
rect 4842 4194 4860 4212
rect 4842 4410 4860 4428
rect 4842 4428 4860 4446
rect 4842 4446 4860 4464
rect 4842 4464 4860 4482
rect 4842 4482 4860 4500
rect 4842 4500 4860 4518
rect 4842 4518 4860 4536
rect 4842 4536 4860 4554
rect 4842 4554 4860 4572
rect 4842 4572 4860 4590
rect 4842 4590 4860 4608
rect 4842 4608 4860 4626
rect 4842 4626 4860 4644
rect 4842 4644 4860 4662
rect 4842 4662 4860 4680
rect 4842 4680 4860 4698
rect 4842 4698 4860 4716
rect 4842 4716 4860 4734
rect 4842 4734 4860 4752
rect 4842 4752 4860 4770
rect 4842 4770 4860 4788
rect 4842 4788 4860 4806
rect 4842 4806 4860 4824
rect 4842 4824 4860 4842
rect 4842 4842 4860 4860
rect 4842 4860 4860 4878
rect 4842 4878 4860 4896
rect 4842 4896 4860 4914
rect 4842 4914 4860 4932
rect 4842 4932 4860 4950
rect 4842 4950 4860 4968
rect 4842 4968 4860 4986
rect 4842 4986 4860 5004
rect 4842 5004 4860 5022
rect 4842 5022 4860 5040
rect 4842 5040 4860 5058
rect 4842 5058 4860 5076
rect 4842 5076 4860 5094
rect 4842 5094 4860 5112
rect 4842 5112 4860 5130
rect 4842 5130 4860 5148
rect 4842 5148 4860 5166
rect 4842 5166 4860 5184
rect 4842 5184 4860 5202
rect 4842 5202 4860 5220
rect 4842 5220 4860 5238
rect 4842 5238 4860 5256
rect 4842 5256 4860 5274
rect 4842 5274 4860 5292
rect 4842 5292 4860 5310
rect 4842 5310 4860 5328
rect 4842 5328 4860 5346
rect 4842 5346 4860 5364
rect 4842 5364 4860 5382
rect 4842 5382 4860 5400
rect 4842 5400 4860 5418
rect 4842 5418 4860 5436
rect 4842 5436 4860 5454
rect 4842 5454 4860 5472
rect 4842 5472 4860 5490
rect 4842 5490 4860 5508
rect 4842 5508 4860 5526
rect 4842 5526 4860 5544
rect 4842 5544 4860 5562
rect 4842 5562 4860 5580
rect 4842 5580 4860 5598
rect 4842 5598 4860 5616
rect 4842 5616 4860 5634
rect 4842 5634 4860 5652
rect 4842 5652 4860 5670
rect 4842 5670 4860 5688
rect 4842 5688 4860 5706
rect 4842 5706 4860 5724
rect 4842 5724 4860 5742
rect 4842 5742 4860 5760
rect 4842 5760 4860 5778
rect 4842 5778 4860 5796
rect 4842 5796 4860 5814
rect 4842 5814 4860 5832
rect 4842 5832 4860 5850
rect 4842 5850 4860 5868
rect 4842 5868 4860 5886
rect 4842 5886 4860 5904
rect 4842 5904 4860 5922
rect 4842 5922 4860 5940
rect 4842 5940 4860 5958
rect 4842 5958 4860 5976
rect 4842 5976 4860 5994
rect 4842 5994 4860 6012
rect 4842 6012 4860 6030
rect 4842 6030 4860 6048
rect 4842 6048 4860 6066
rect 4842 6066 4860 6084
rect 4842 6084 4860 6102
rect 4842 6102 4860 6120
rect 4842 6120 4860 6138
rect 4842 6138 4860 6156
rect 4842 6156 4860 6174
rect 4842 6174 4860 6192
rect 4842 6192 4860 6210
rect 4842 6210 4860 6228
rect 4842 6228 4860 6246
rect 4842 6246 4860 6264
rect 4842 6264 4860 6282
rect 4842 6282 4860 6300
rect 4842 6300 4860 6318
rect 4842 6318 4860 6336
rect 4842 6336 4860 6354
rect 4842 6354 4860 6372
rect 4842 6372 4860 6390
rect 4842 6390 4860 6408
rect 4842 6408 4860 6426
rect 4842 6426 4860 6444
rect 4842 6444 4860 6462
rect 4842 6462 4860 6480
rect 4842 6480 4860 6498
rect 4842 6498 4860 6516
rect 4842 6516 4860 6534
rect 4842 6534 4860 6552
rect 4842 6552 4860 6570
rect 4842 6570 4860 6588
rect 4842 6588 4860 6606
rect 4842 6606 4860 6624
rect 4842 6624 4860 6642
rect 4842 6642 4860 6660
rect 4842 6660 4860 6678
rect 4842 6678 4860 6696
rect 4842 6696 4860 6714
rect 4842 6714 4860 6732
rect 4842 6732 4860 6750
rect 4842 6750 4860 6768
rect 4842 6768 4860 6786
rect 4842 6786 4860 6804
rect 4842 6804 4860 6822
rect 4842 6822 4860 6840
rect 4842 6840 4860 6858
rect 4842 6858 4860 6876
rect 4842 6876 4860 6894
rect 4842 6894 4860 6912
rect 4842 6912 4860 6930
rect 4842 6930 4860 6948
rect 4842 6948 4860 6966
rect 4842 6966 4860 6984
rect 4842 6984 4860 7002
rect 4842 7002 4860 7020
rect 4842 7020 4860 7038
rect 4842 7038 4860 7056
rect 4842 7056 4860 7074
rect 4842 7074 4860 7092
rect 4842 7092 4860 7110
rect 4842 7110 4860 7128
rect 4842 7128 4860 7146
rect 4842 7146 4860 7164
rect 4842 7164 4860 7182
rect 4842 7182 4860 7200
rect 4842 7200 4860 7218
rect 4842 7218 4860 7236
rect 4842 7236 4860 7254
rect 4842 7254 4860 7272
rect 4842 7272 4860 7290
rect 4842 7290 4860 7308
rect 4842 7308 4860 7326
rect 4842 7326 4860 7344
rect 4842 7344 4860 7362
rect 4842 7362 4860 7380
rect 4842 7380 4860 7398
rect 4842 7398 4860 7416
rect 4842 7416 4860 7434
rect 4842 7434 4860 7452
rect 4842 7452 4860 7470
rect 4842 7470 4860 7488
rect 4842 7488 4860 7506
rect 4842 7506 4860 7524
rect 4842 7524 4860 7542
rect 4842 7542 4860 7560
rect 4842 7560 4860 7578
rect 4842 7578 4860 7596
rect 4860 216 4878 234
rect 4860 234 4878 252
rect 4860 252 4878 270
rect 4860 270 4878 288
rect 4860 288 4878 306
rect 4860 306 4878 324
rect 4860 324 4878 342
rect 4860 342 4878 360
rect 4860 360 4878 378
rect 4860 378 4878 396
rect 4860 396 4878 414
rect 4860 414 4878 432
rect 4860 432 4878 450
rect 4860 450 4878 468
rect 4860 468 4878 486
rect 4860 486 4878 504
rect 4860 504 4878 522
rect 4860 522 4878 540
rect 4860 540 4878 558
rect 4860 558 4878 576
rect 4860 576 4878 594
rect 4860 594 4878 612
rect 4860 612 4878 630
rect 4860 630 4878 648
rect 4860 648 4878 666
rect 4860 666 4878 684
rect 4860 684 4878 702
rect 4860 702 4878 720
rect 4860 720 4878 738
rect 4860 738 4878 756
rect 4860 864 4878 882
rect 4860 882 4878 900
rect 4860 900 4878 918
rect 4860 918 4878 936
rect 4860 936 4878 954
rect 4860 954 4878 972
rect 4860 972 4878 990
rect 4860 990 4878 1008
rect 4860 1008 4878 1026
rect 4860 1026 4878 1044
rect 4860 1044 4878 1062
rect 4860 1062 4878 1080
rect 4860 1080 4878 1098
rect 4860 1098 4878 1116
rect 4860 1116 4878 1134
rect 4860 1134 4878 1152
rect 4860 1152 4878 1170
rect 4860 1170 4878 1188
rect 4860 1188 4878 1206
rect 4860 1206 4878 1224
rect 4860 1224 4878 1242
rect 4860 1242 4878 1260
rect 4860 1260 4878 1278
rect 4860 1278 4878 1296
rect 4860 1296 4878 1314
rect 4860 1314 4878 1332
rect 4860 1332 4878 1350
rect 4860 1350 4878 1368
rect 4860 1368 4878 1386
rect 4860 1386 4878 1404
rect 4860 1404 4878 1422
rect 4860 1422 4878 1440
rect 4860 1440 4878 1458
rect 4860 1458 4878 1476
rect 4860 1476 4878 1494
rect 4860 1494 4878 1512
rect 4860 1512 4878 1530
rect 4860 1530 4878 1548
rect 4860 1548 4878 1566
rect 4860 1566 4878 1584
rect 4860 1584 4878 1602
rect 4860 1602 4878 1620
rect 4860 1620 4878 1638
rect 4860 1638 4878 1656
rect 4860 1656 4878 1674
rect 4860 1674 4878 1692
rect 4860 1692 4878 1710
rect 4860 1710 4878 1728
rect 4860 1728 4878 1746
rect 4860 1746 4878 1764
rect 4860 1764 4878 1782
rect 4860 1782 4878 1800
rect 4860 1800 4878 1818
rect 4860 1818 4878 1836
rect 4860 1836 4878 1854
rect 4860 1854 4878 1872
rect 4860 1872 4878 1890
rect 4860 1890 4878 1908
rect 4860 1908 4878 1926
rect 4860 1926 4878 1944
rect 4860 1944 4878 1962
rect 4860 1962 4878 1980
rect 4860 1980 4878 1998
rect 4860 1998 4878 2016
rect 4860 2016 4878 2034
rect 4860 2034 4878 2052
rect 4860 2052 4878 2070
rect 4860 2070 4878 2088
rect 4860 2088 4878 2106
rect 4860 2106 4878 2124
rect 4860 2124 4878 2142
rect 4860 2358 4878 2376
rect 4860 2376 4878 2394
rect 4860 2394 4878 2412
rect 4860 2412 4878 2430
rect 4860 2430 4878 2448
rect 4860 2448 4878 2466
rect 4860 2466 4878 2484
rect 4860 2484 4878 2502
rect 4860 2502 4878 2520
rect 4860 2520 4878 2538
rect 4860 2538 4878 2556
rect 4860 2556 4878 2574
rect 4860 2574 4878 2592
rect 4860 2592 4878 2610
rect 4860 2610 4878 2628
rect 4860 2628 4878 2646
rect 4860 2646 4878 2664
rect 4860 2664 4878 2682
rect 4860 2682 4878 2700
rect 4860 2700 4878 2718
rect 4860 2718 4878 2736
rect 4860 2736 4878 2754
rect 4860 2754 4878 2772
rect 4860 2772 4878 2790
rect 4860 2790 4878 2808
rect 4860 2808 4878 2826
rect 4860 2826 4878 2844
rect 4860 2844 4878 2862
rect 4860 2862 4878 2880
rect 4860 2880 4878 2898
rect 4860 2898 4878 2916
rect 4860 2916 4878 2934
rect 4860 2934 4878 2952
rect 4860 2952 4878 2970
rect 4860 2970 4878 2988
rect 4860 2988 4878 3006
rect 4860 3006 4878 3024
rect 4860 3024 4878 3042
rect 4860 3042 4878 3060
rect 4860 3060 4878 3078
rect 4860 3078 4878 3096
rect 4860 3096 4878 3114
rect 4860 3114 4878 3132
rect 4860 3132 4878 3150
rect 4860 3150 4878 3168
rect 4860 3168 4878 3186
rect 4860 3186 4878 3204
rect 4860 3204 4878 3222
rect 4860 3222 4878 3240
rect 4860 3240 4878 3258
rect 4860 3258 4878 3276
rect 4860 3276 4878 3294
rect 4860 3294 4878 3312
rect 4860 3312 4878 3330
rect 4860 3330 4878 3348
rect 4860 3348 4878 3366
rect 4860 3366 4878 3384
rect 4860 3384 4878 3402
rect 4860 3402 4878 3420
rect 4860 3420 4878 3438
rect 4860 3438 4878 3456
rect 4860 3456 4878 3474
rect 4860 3474 4878 3492
rect 4860 3492 4878 3510
rect 4860 3510 4878 3528
rect 4860 3528 4878 3546
rect 4860 3546 4878 3564
rect 4860 3564 4878 3582
rect 4860 3582 4878 3600
rect 4860 3600 4878 3618
rect 4860 3618 4878 3636
rect 4860 3636 4878 3654
rect 4860 3654 4878 3672
rect 4860 3672 4878 3690
rect 4860 3690 4878 3708
rect 4860 3708 4878 3726
rect 4860 3726 4878 3744
rect 4860 3744 4878 3762
rect 4860 3762 4878 3780
rect 4860 3780 4878 3798
rect 4860 3798 4878 3816
rect 4860 3816 4878 3834
rect 4860 3834 4878 3852
rect 4860 3852 4878 3870
rect 4860 3870 4878 3888
rect 4860 3888 4878 3906
rect 4860 3906 4878 3924
rect 4860 3924 4878 3942
rect 4860 3942 4878 3960
rect 4860 3960 4878 3978
rect 4860 3978 4878 3996
rect 4860 3996 4878 4014
rect 4860 4014 4878 4032
rect 4860 4032 4878 4050
rect 4860 4050 4878 4068
rect 4860 4068 4878 4086
rect 4860 4086 4878 4104
rect 4860 4104 4878 4122
rect 4860 4122 4878 4140
rect 4860 4140 4878 4158
rect 4860 4158 4878 4176
rect 4860 4176 4878 4194
rect 4860 4194 4878 4212
rect 4860 4212 4878 4230
rect 4860 4428 4878 4446
rect 4860 4446 4878 4464
rect 4860 4464 4878 4482
rect 4860 4482 4878 4500
rect 4860 4500 4878 4518
rect 4860 4518 4878 4536
rect 4860 4536 4878 4554
rect 4860 4554 4878 4572
rect 4860 4572 4878 4590
rect 4860 4590 4878 4608
rect 4860 4608 4878 4626
rect 4860 4626 4878 4644
rect 4860 4644 4878 4662
rect 4860 4662 4878 4680
rect 4860 4680 4878 4698
rect 4860 4698 4878 4716
rect 4860 4716 4878 4734
rect 4860 4734 4878 4752
rect 4860 4752 4878 4770
rect 4860 4770 4878 4788
rect 4860 4788 4878 4806
rect 4860 4806 4878 4824
rect 4860 4824 4878 4842
rect 4860 4842 4878 4860
rect 4860 4860 4878 4878
rect 4860 4878 4878 4896
rect 4860 4896 4878 4914
rect 4860 4914 4878 4932
rect 4860 4932 4878 4950
rect 4860 4950 4878 4968
rect 4860 4968 4878 4986
rect 4860 4986 4878 5004
rect 4860 5004 4878 5022
rect 4860 5022 4878 5040
rect 4860 5040 4878 5058
rect 4860 5058 4878 5076
rect 4860 5076 4878 5094
rect 4860 5094 4878 5112
rect 4860 5112 4878 5130
rect 4860 5130 4878 5148
rect 4860 5148 4878 5166
rect 4860 5166 4878 5184
rect 4860 5184 4878 5202
rect 4860 5202 4878 5220
rect 4860 5220 4878 5238
rect 4860 5238 4878 5256
rect 4860 5256 4878 5274
rect 4860 5274 4878 5292
rect 4860 5292 4878 5310
rect 4860 5310 4878 5328
rect 4860 5328 4878 5346
rect 4860 5346 4878 5364
rect 4860 5364 4878 5382
rect 4860 5382 4878 5400
rect 4860 5400 4878 5418
rect 4860 5418 4878 5436
rect 4860 5436 4878 5454
rect 4860 5454 4878 5472
rect 4860 5472 4878 5490
rect 4860 5490 4878 5508
rect 4860 5508 4878 5526
rect 4860 5526 4878 5544
rect 4860 5544 4878 5562
rect 4860 5562 4878 5580
rect 4860 5580 4878 5598
rect 4860 5598 4878 5616
rect 4860 5616 4878 5634
rect 4860 5634 4878 5652
rect 4860 5652 4878 5670
rect 4860 5670 4878 5688
rect 4860 5688 4878 5706
rect 4860 5706 4878 5724
rect 4860 5724 4878 5742
rect 4860 5742 4878 5760
rect 4860 5760 4878 5778
rect 4860 5778 4878 5796
rect 4860 5796 4878 5814
rect 4860 5814 4878 5832
rect 4860 5832 4878 5850
rect 4860 5850 4878 5868
rect 4860 5868 4878 5886
rect 4860 5886 4878 5904
rect 4860 5904 4878 5922
rect 4860 5922 4878 5940
rect 4860 5940 4878 5958
rect 4860 5958 4878 5976
rect 4860 5976 4878 5994
rect 4860 5994 4878 6012
rect 4860 6012 4878 6030
rect 4860 6030 4878 6048
rect 4860 6048 4878 6066
rect 4860 6066 4878 6084
rect 4860 6084 4878 6102
rect 4860 6102 4878 6120
rect 4860 6120 4878 6138
rect 4860 6138 4878 6156
rect 4860 6156 4878 6174
rect 4860 6174 4878 6192
rect 4860 6192 4878 6210
rect 4860 6210 4878 6228
rect 4860 6228 4878 6246
rect 4860 6246 4878 6264
rect 4860 6264 4878 6282
rect 4860 6282 4878 6300
rect 4860 6300 4878 6318
rect 4860 6318 4878 6336
rect 4860 6336 4878 6354
rect 4860 6354 4878 6372
rect 4860 6372 4878 6390
rect 4860 6390 4878 6408
rect 4860 6408 4878 6426
rect 4860 6426 4878 6444
rect 4860 6444 4878 6462
rect 4860 6462 4878 6480
rect 4860 6480 4878 6498
rect 4860 6498 4878 6516
rect 4860 6516 4878 6534
rect 4860 6534 4878 6552
rect 4860 6552 4878 6570
rect 4860 6570 4878 6588
rect 4860 6588 4878 6606
rect 4860 6606 4878 6624
rect 4860 6624 4878 6642
rect 4860 6642 4878 6660
rect 4860 6660 4878 6678
rect 4860 6678 4878 6696
rect 4860 6696 4878 6714
rect 4860 6714 4878 6732
rect 4860 6732 4878 6750
rect 4860 6750 4878 6768
rect 4860 6768 4878 6786
rect 4860 6786 4878 6804
rect 4860 6804 4878 6822
rect 4860 6822 4878 6840
rect 4860 6840 4878 6858
rect 4860 6858 4878 6876
rect 4860 6876 4878 6894
rect 4860 6894 4878 6912
rect 4860 6912 4878 6930
rect 4860 6930 4878 6948
rect 4860 6948 4878 6966
rect 4860 6966 4878 6984
rect 4860 6984 4878 7002
rect 4860 7002 4878 7020
rect 4860 7020 4878 7038
rect 4860 7038 4878 7056
rect 4860 7056 4878 7074
rect 4860 7074 4878 7092
rect 4860 7092 4878 7110
rect 4860 7110 4878 7128
rect 4860 7128 4878 7146
rect 4860 7146 4878 7164
rect 4860 7164 4878 7182
rect 4860 7182 4878 7200
rect 4860 7200 4878 7218
rect 4860 7218 4878 7236
rect 4860 7236 4878 7254
rect 4860 7254 4878 7272
rect 4860 7272 4878 7290
rect 4860 7290 4878 7308
rect 4860 7308 4878 7326
rect 4860 7326 4878 7344
rect 4860 7344 4878 7362
rect 4860 7362 4878 7380
rect 4860 7380 4878 7398
rect 4860 7398 4878 7416
rect 4860 7416 4878 7434
rect 4860 7434 4878 7452
rect 4860 7452 4878 7470
rect 4860 7470 4878 7488
rect 4860 7488 4878 7506
rect 4860 7506 4878 7524
rect 4860 7524 4878 7542
rect 4860 7542 4878 7560
rect 4860 7560 4878 7578
rect 4860 7578 4878 7596
rect 4860 7596 4878 7614
rect 4860 7614 4878 7632
rect 4878 216 4896 234
rect 4878 234 4896 252
rect 4878 252 4896 270
rect 4878 270 4896 288
rect 4878 288 4896 306
rect 4878 306 4896 324
rect 4878 324 4896 342
rect 4878 342 4896 360
rect 4878 360 4896 378
rect 4878 378 4896 396
rect 4878 396 4896 414
rect 4878 414 4896 432
rect 4878 432 4896 450
rect 4878 450 4896 468
rect 4878 468 4896 486
rect 4878 486 4896 504
rect 4878 504 4896 522
rect 4878 522 4896 540
rect 4878 540 4896 558
rect 4878 558 4896 576
rect 4878 576 4896 594
rect 4878 594 4896 612
rect 4878 612 4896 630
rect 4878 630 4896 648
rect 4878 648 4896 666
rect 4878 666 4896 684
rect 4878 684 4896 702
rect 4878 702 4896 720
rect 4878 720 4896 738
rect 4878 738 4896 756
rect 4878 864 4896 882
rect 4878 882 4896 900
rect 4878 900 4896 918
rect 4878 918 4896 936
rect 4878 936 4896 954
rect 4878 954 4896 972
rect 4878 972 4896 990
rect 4878 990 4896 1008
rect 4878 1008 4896 1026
rect 4878 1026 4896 1044
rect 4878 1044 4896 1062
rect 4878 1062 4896 1080
rect 4878 1080 4896 1098
rect 4878 1098 4896 1116
rect 4878 1116 4896 1134
rect 4878 1134 4896 1152
rect 4878 1152 4896 1170
rect 4878 1170 4896 1188
rect 4878 1188 4896 1206
rect 4878 1206 4896 1224
rect 4878 1224 4896 1242
rect 4878 1242 4896 1260
rect 4878 1260 4896 1278
rect 4878 1278 4896 1296
rect 4878 1296 4896 1314
rect 4878 1314 4896 1332
rect 4878 1332 4896 1350
rect 4878 1350 4896 1368
rect 4878 1368 4896 1386
rect 4878 1386 4896 1404
rect 4878 1404 4896 1422
rect 4878 1422 4896 1440
rect 4878 1440 4896 1458
rect 4878 1458 4896 1476
rect 4878 1476 4896 1494
rect 4878 1494 4896 1512
rect 4878 1512 4896 1530
rect 4878 1530 4896 1548
rect 4878 1548 4896 1566
rect 4878 1566 4896 1584
rect 4878 1584 4896 1602
rect 4878 1602 4896 1620
rect 4878 1620 4896 1638
rect 4878 1638 4896 1656
rect 4878 1656 4896 1674
rect 4878 1674 4896 1692
rect 4878 1692 4896 1710
rect 4878 1710 4896 1728
rect 4878 1728 4896 1746
rect 4878 1746 4896 1764
rect 4878 1764 4896 1782
rect 4878 1782 4896 1800
rect 4878 1800 4896 1818
rect 4878 1818 4896 1836
rect 4878 1836 4896 1854
rect 4878 1854 4896 1872
rect 4878 1872 4896 1890
rect 4878 1890 4896 1908
rect 4878 1908 4896 1926
rect 4878 1926 4896 1944
rect 4878 1944 4896 1962
rect 4878 1962 4896 1980
rect 4878 1980 4896 1998
rect 4878 1998 4896 2016
rect 4878 2016 4896 2034
rect 4878 2034 4896 2052
rect 4878 2052 4896 2070
rect 4878 2070 4896 2088
rect 4878 2088 4896 2106
rect 4878 2106 4896 2124
rect 4878 2124 4896 2142
rect 4878 2142 4896 2160
rect 4878 2376 4896 2394
rect 4878 2394 4896 2412
rect 4878 2412 4896 2430
rect 4878 2430 4896 2448
rect 4878 2448 4896 2466
rect 4878 2466 4896 2484
rect 4878 2484 4896 2502
rect 4878 2502 4896 2520
rect 4878 2520 4896 2538
rect 4878 2538 4896 2556
rect 4878 2556 4896 2574
rect 4878 2574 4896 2592
rect 4878 2592 4896 2610
rect 4878 2610 4896 2628
rect 4878 2628 4896 2646
rect 4878 2646 4896 2664
rect 4878 2664 4896 2682
rect 4878 2682 4896 2700
rect 4878 2700 4896 2718
rect 4878 2718 4896 2736
rect 4878 2736 4896 2754
rect 4878 2754 4896 2772
rect 4878 2772 4896 2790
rect 4878 2790 4896 2808
rect 4878 2808 4896 2826
rect 4878 2826 4896 2844
rect 4878 2844 4896 2862
rect 4878 2862 4896 2880
rect 4878 2880 4896 2898
rect 4878 2898 4896 2916
rect 4878 2916 4896 2934
rect 4878 2934 4896 2952
rect 4878 2952 4896 2970
rect 4878 2970 4896 2988
rect 4878 2988 4896 3006
rect 4878 3006 4896 3024
rect 4878 3024 4896 3042
rect 4878 3042 4896 3060
rect 4878 3060 4896 3078
rect 4878 3078 4896 3096
rect 4878 3096 4896 3114
rect 4878 3114 4896 3132
rect 4878 3132 4896 3150
rect 4878 3150 4896 3168
rect 4878 3168 4896 3186
rect 4878 3186 4896 3204
rect 4878 3204 4896 3222
rect 4878 3222 4896 3240
rect 4878 3240 4896 3258
rect 4878 3258 4896 3276
rect 4878 3276 4896 3294
rect 4878 3294 4896 3312
rect 4878 3312 4896 3330
rect 4878 3330 4896 3348
rect 4878 3348 4896 3366
rect 4878 3366 4896 3384
rect 4878 3384 4896 3402
rect 4878 3402 4896 3420
rect 4878 3420 4896 3438
rect 4878 3438 4896 3456
rect 4878 3456 4896 3474
rect 4878 3474 4896 3492
rect 4878 3492 4896 3510
rect 4878 3510 4896 3528
rect 4878 3528 4896 3546
rect 4878 3546 4896 3564
rect 4878 3564 4896 3582
rect 4878 3582 4896 3600
rect 4878 3600 4896 3618
rect 4878 3618 4896 3636
rect 4878 3636 4896 3654
rect 4878 3654 4896 3672
rect 4878 3672 4896 3690
rect 4878 3690 4896 3708
rect 4878 3708 4896 3726
rect 4878 3726 4896 3744
rect 4878 3744 4896 3762
rect 4878 3762 4896 3780
rect 4878 3780 4896 3798
rect 4878 3798 4896 3816
rect 4878 3816 4896 3834
rect 4878 3834 4896 3852
rect 4878 3852 4896 3870
rect 4878 3870 4896 3888
rect 4878 3888 4896 3906
rect 4878 3906 4896 3924
rect 4878 3924 4896 3942
rect 4878 3942 4896 3960
rect 4878 3960 4896 3978
rect 4878 3978 4896 3996
rect 4878 3996 4896 4014
rect 4878 4014 4896 4032
rect 4878 4032 4896 4050
rect 4878 4050 4896 4068
rect 4878 4068 4896 4086
rect 4878 4086 4896 4104
rect 4878 4104 4896 4122
rect 4878 4122 4896 4140
rect 4878 4140 4896 4158
rect 4878 4158 4896 4176
rect 4878 4176 4896 4194
rect 4878 4194 4896 4212
rect 4878 4212 4896 4230
rect 4878 4230 4896 4248
rect 4878 4446 4896 4464
rect 4878 4464 4896 4482
rect 4878 4482 4896 4500
rect 4878 4500 4896 4518
rect 4878 4518 4896 4536
rect 4878 4536 4896 4554
rect 4878 4554 4896 4572
rect 4878 4572 4896 4590
rect 4878 4590 4896 4608
rect 4878 4608 4896 4626
rect 4878 4626 4896 4644
rect 4878 4644 4896 4662
rect 4878 4662 4896 4680
rect 4878 4680 4896 4698
rect 4878 4698 4896 4716
rect 4878 4716 4896 4734
rect 4878 4734 4896 4752
rect 4878 4752 4896 4770
rect 4878 4770 4896 4788
rect 4878 4788 4896 4806
rect 4878 4806 4896 4824
rect 4878 4824 4896 4842
rect 4878 4842 4896 4860
rect 4878 4860 4896 4878
rect 4878 4878 4896 4896
rect 4878 4896 4896 4914
rect 4878 4914 4896 4932
rect 4878 4932 4896 4950
rect 4878 4950 4896 4968
rect 4878 4968 4896 4986
rect 4878 4986 4896 5004
rect 4878 5004 4896 5022
rect 4878 5022 4896 5040
rect 4878 5040 4896 5058
rect 4878 5058 4896 5076
rect 4878 5076 4896 5094
rect 4878 5094 4896 5112
rect 4878 5112 4896 5130
rect 4878 5130 4896 5148
rect 4878 5148 4896 5166
rect 4878 5166 4896 5184
rect 4878 5184 4896 5202
rect 4878 5202 4896 5220
rect 4878 5220 4896 5238
rect 4878 5238 4896 5256
rect 4878 5256 4896 5274
rect 4878 5274 4896 5292
rect 4878 5292 4896 5310
rect 4878 5310 4896 5328
rect 4878 5328 4896 5346
rect 4878 5346 4896 5364
rect 4878 5364 4896 5382
rect 4878 5382 4896 5400
rect 4878 5400 4896 5418
rect 4878 5418 4896 5436
rect 4878 5436 4896 5454
rect 4878 5454 4896 5472
rect 4878 5472 4896 5490
rect 4878 5490 4896 5508
rect 4878 5508 4896 5526
rect 4878 5526 4896 5544
rect 4878 5544 4896 5562
rect 4878 5562 4896 5580
rect 4878 5580 4896 5598
rect 4878 5598 4896 5616
rect 4878 5616 4896 5634
rect 4878 5634 4896 5652
rect 4878 5652 4896 5670
rect 4878 5670 4896 5688
rect 4878 5688 4896 5706
rect 4878 5706 4896 5724
rect 4878 5724 4896 5742
rect 4878 5742 4896 5760
rect 4878 5760 4896 5778
rect 4878 5778 4896 5796
rect 4878 5796 4896 5814
rect 4878 5814 4896 5832
rect 4878 5832 4896 5850
rect 4878 5850 4896 5868
rect 4878 5868 4896 5886
rect 4878 5886 4896 5904
rect 4878 5904 4896 5922
rect 4878 5922 4896 5940
rect 4878 5940 4896 5958
rect 4878 5958 4896 5976
rect 4878 5976 4896 5994
rect 4878 5994 4896 6012
rect 4878 6012 4896 6030
rect 4878 6030 4896 6048
rect 4878 6048 4896 6066
rect 4878 6066 4896 6084
rect 4878 6084 4896 6102
rect 4878 6102 4896 6120
rect 4878 6120 4896 6138
rect 4878 6138 4896 6156
rect 4878 6156 4896 6174
rect 4878 6174 4896 6192
rect 4878 6192 4896 6210
rect 4878 6210 4896 6228
rect 4878 6228 4896 6246
rect 4878 6246 4896 6264
rect 4878 6264 4896 6282
rect 4878 6282 4896 6300
rect 4878 6300 4896 6318
rect 4878 6318 4896 6336
rect 4878 6336 4896 6354
rect 4878 6354 4896 6372
rect 4878 6372 4896 6390
rect 4878 6390 4896 6408
rect 4878 6408 4896 6426
rect 4878 6426 4896 6444
rect 4878 6444 4896 6462
rect 4878 6462 4896 6480
rect 4878 6480 4896 6498
rect 4878 6498 4896 6516
rect 4878 6516 4896 6534
rect 4878 6534 4896 6552
rect 4878 6552 4896 6570
rect 4878 6570 4896 6588
rect 4878 6588 4896 6606
rect 4878 6606 4896 6624
rect 4878 6624 4896 6642
rect 4878 6642 4896 6660
rect 4878 6660 4896 6678
rect 4878 6678 4896 6696
rect 4878 6696 4896 6714
rect 4878 6714 4896 6732
rect 4878 6732 4896 6750
rect 4878 6750 4896 6768
rect 4878 6768 4896 6786
rect 4878 6786 4896 6804
rect 4878 6804 4896 6822
rect 4878 6822 4896 6840
rect 4878 6840 4896 6858
rect 4878 6858 4896 6876
rect 4878 6876 4896 6894
rect 4878 6894 4896 6912
rect 4878 6912 4896 6930
rect 4878 6930 4896 6948
rect 4878 6948 4896 6966
rect 4878 6966 4896 6984
rect 4878 6984 4896 7002
rect 4878 7002 4896 7020
rect 4878 7020 4896 7038
rect 4878 7038 4896 7056
rect 4878 7056 4896 7074
rect 4878 7074 4896 7092
rect 4878 7092 4896 7110
rect 4878 7110 4896 7128
rect 4878 7128 4896 7146
rect 4878 7146 4896 7164
rect 4878 7164 4896 7182
rect 4878 7182 4896 7200
rect 4878 7200 4896 7218
rect 4878 7218 4896 7236
rect 4878 7236 4896 7254
rect 4878 7254 4896 7272
rect 4878 7272 4896 7290
rect 4878 7290 4896 7308
rect 4878 7308 4896 7326
rect 4878 7326 4896 7344
rect 4878 7344 4896 7362
rect 4878 7362 4896 7380
rect 4878 7380 4896 7398
rect 4878 7398 4896 7416
rect 4878 7416 4896 7434
rect 4878 7434 4896 7452
rect 4878 7452 4896 7470
rect 4878 7470 4896 7488
rect 4878 7488 4896 7506
rect 4878 7506 4896 7524
rect 4878 7524 4896 7542
rect 4878 7542 4896 7560
rect 4878 7560 4896 7578
rect 4878 7578 4896 7596
rect 4878 7596 4896 7614
rect 4878 7614 4896 7632
rect 4878 7632 4896 7650
rect 4896 216 4914 234
rect 4896 234 4914 252
rect 4896 252 4914 270
rect 4896 270 4914 288
rect 4896 288 4914 306
rect 4896 306 4914 324
rect 4896 324 4914 342
rect 4896 342 4914 360
rect 4896 360 4914 378
rect 4896 378 4914 396
rect 4896 396 4914 414
rect 4896 414 4914 432
rect 4896 432 4914 450
rect 4896 450 4914 468
rect 4896 468 4914 486
rect 4896 486 4914 504
rect 4896 504 4914 522
rect 4896 522 4914 540
rect 4896 540 4914 558
rect 4896 558 4914 576
rect 4896 576 4914 594
rect 4896 594 4914 612
rect 4896 612 4914 630
rect 4896 630 4914 648
rect 4896 648 4914 666
rect 4896 666 4914 684
rect 4896 684 4914 702
rect 4896 702 4914 720
rect 4896 720 4914 738
rect 4896 738 4914 756
rect 4896 864 4914 882
rect 4896 882 4914 900
rect 4896 900 4914 918
rect 4896 918 4914 936
rect 4896 936 4914 954
rect 4896 954 4914 972
rect 4896 972 4914 990
rect 4896 990 4914 1008
rect 4896 1008 4914 1026
rect 4896 1026 4914 1044
rect 4896 1044 4914 1062
rect 4896 1062 4914 1080
rect 4896 1080 4914 1098
rect 4896 1098 4914 1116
rect 4896 1116 4914 1134
rect 4896 1134 4914 1152
rect 4896 1152 4914 1170
rect 4896 1170 4914 1188
rect 4896 1188 4914 1206
rect 4896 1206 4914 1224
rect 4896 1224 4914 1242
rect 4896 1242 4914 1260
rect 4896 1260 4914 1278
rect 4896 1278 4914 1296
rect 4896 1296 4914 1314
rect 4896 1314 4914 1332
rect 4896 1332 4914 1350
rect 4896 1350 4914 1368
rect 4896 1368 4914 1386
rect 4896 1386 4914 1404
rect 4896 1404 4914 1422
rect 4896 1422 4914 1440
rect 4896 1440 4914 1458
rect 4896 1458 4914 1476
rect 4896 1476 4914 1494
rect 4896 1494 4914 1512
rect 4896 1512 4914 1530
rect 4896 1530 4914 1548
rect 4896 1548 4914 1566
rect 4896 1566 4914 1584
rect 4896 1584 4914 1602
rect 4896 1602 4914 1620
rect 4896 1620 4914 1638
rect 4896 1638 4914 1656
rect 4896 1656 4914 1674
rect 4896 1674 4914 1692
rect 4896 1692 4914 1710
rect 4896 1710 4914 1728
rect 4896 1728 4914 1746
rect 4896 1746 4914 1764
rect 4896 1764 4914 1782
rect 4896 1782 4914 1800
rect 4896 1800 4914 1818
rect 4896 1818 4914 1836
rect 4896 1836 4914 1854
rect 4896 1854 4914 1872
rect 4896 1872 4914 1890
rect 4896 1890 4914 1908
rect 4896 1908 4914 1926
rect 4896 1926 4914 1944
rect 4896 1944 4914 1962
rect 4896 1962 4914 1980
rect 4896 1980 4914 1998
rect 4896 1998 4914 2016
rect 4896 2016 4914 2034
rect 4896 2034 4914 2052
rect 4896 2052 4914 2070
rect 4896 2070 4914 2088
rect 4896 2088 4914 2106
rect 4896 2106 4914 2124
rect 4896 2124 4914 2142
rect 4896 2142 4914 2160
rect 4896 2376 4914 2394
rect 4896 2394 4914 2412
rect 4896 2412 4914 2430
rect 4896 2430 4914 2448
rect 4896 2448 4914 2466
rect 4896 2466 4914 2484
rect 4896 2484 4914 2502
rect 4896 2502 4914 2520
rect 4896 2520 4914 2538
rect 4896 2538 4914 2556
rect 4896 2556 4914 2574
rect 4896 2574 4914 2592
rect 4896 2592 4914 2610
rect 4896 2610 4914 2628
rect 4896 2628 4914 2646
rect 4896 2646 4914 2664
rect 4896 2664 4914 2682
rect 4896 2682 4914 2700
rect 4896 2700 4914 2718
rect 4896 2718 4914 2736
rect 4896 2736 4914 2754
rect 4896 2754 4914 2772
rect 4896 2772 4914 2790
rect 4896 2790 4914 2808
rect 4896 2808 4914 2826
rect 4896 2826 4914 2844
rect 4896 2844 4914 2862
rect 4896 2862 4914 2880
rect 4896 2880 4914 2898
rect 4896 2898 4914 2916
rect 4896 2916 4914 2934
rect 4896 2934 4914 2952
rect 4896 2952 4914 2970
rect 4896 2970 4914 2988
rect 4896 2988 4914 3006
rect 4896 3006 4914 3024
rect 4896 3024 4914 3042
rect 4896 3042 4914 3060
rect 4896 3060 4914 3078
rect 4896 3078 4914 3096
rect 4896 3096 4914 3114
rect 4896 3114 4914 3132
rect 4896 3132 4914 3150
rect 4896 3150 4914 3168
rect 4896 3168 4914 3186
rect 4896 3186 4914 3204
rect 4896 3204 4914 3222
rect 4896 3222 4914 3240
rect 4896 3240 4914 3258
rect 4896 3258 4914 3276
rect 4896 3276 4914 3294
rect 4896 3294 4914 3312
rect 4896 3312 4914 3330
rect 4896 3330 4914 3348
rect 4896 3348 4914 3366
rect 4896 3366 4914 3384
rect 4896 3384 4914 3402
rect 4896 3402 4914 3420
rect 4896 3420 4914 3438
rect 4896 3438 4914 3456
rect 4896 3456 4914 3474
rect 4896 3474 4914 3492
rect 4896 3492 4914 3510
rect 4896 3510 4914 3528
rect 4896 3528 4914 3546
rect 4896 3546 4914 3564
rect 4896 3564 4914 3582
rect 4896 3582 4914 3600
rect 4896 3600 4914 3618
rect 4896 3618 4914 3636
rect 4896 3636 4914 3654
rect 4896 3654 4914 3672
rect 4896 3672 4914 3690
rect 4896 3690 4914 3708
rect 4896 3708 4914 3726
rect 4896 3726 4914 3744
rect 4896 3744 4914 3762
rect 4896 3762 4914 3780
rect 4896 3780 4914 3798
rect 4896 3798 4914 3816
rect 4896 3816 4914 3834
rect 4896 3834 4914 3852
rect 4896 3852 4914 3870
rect 4896 3870 4914 3888
rect 4896 3888 4914 3906
rect 4896 3906 4914 3924
rect 4896 3924 4914 3942
rect 4896 3942 4914 3960
rect 4896 3960 4914 3978
rect 4896 3978 4914 3996
rect 4896 3996 4914 4014
rect 4896 4014 4914 4032
rect 4896 4032 4914 4050
rect 4896 4050 4914 4068
rect 4896 4068 4914 4086
rect 4896 4086 4914 4104
rect 4896 4104 4914 4122
rect 4896 4122 4914 4140
rect 4896 4140 4914 4158
rect 4896 4158 4914 4176
rect 4896 4176 4914 4194
rect 4896 4194 4914 4212
rect 4896 4212 4914 4230
rect 4896 4230 4914 4248
rect 4896 4248 4914 4266
rect 4896 4482 4914 4500
rect 4896 4500 4914 4518
rect 4896 4518 4914 4536
rect 4896 4536 4914 4554
rect 4896 4554 4914 4572
rect 4896 4572 4914 4590
rect 4896 4590 4914 4608
rect 4896 4608 4914 4626
rect 4896 4626 4914 4644
rect 4896 4644 4914 4662
rect 4896 4662 4914 4680
rect 4896 4680 4914 4698
rect 4896 4698 4914 4716
rect 4896 4716 4914 4734
rect 4896 4734 4914 4752
rect 4896 4752 4914 4770
rect 4896 4770 4914 4788
rect 4896 4788 4914 4806
rect 4896 4806 4914 4824
rect 4896 4824 4914 4842
rect 4896 4842 4914 4860
rect 4896 4860 4914 4878
rect 4896 4878 4914 4896
rect 4896 4896 4914 4914
rect 4896 4914 4914 4932
rect 4896 4932 4914 4950
rect 4896 4950 4914 4968
rect 4896 4968 4914 4986
rect 4896 4986 4914 5004
rect 4896 5004 4914 5022
rect 4896 5022 4914 5040
rect 4896 5040 4914 5058
rect 4896 5058 4914 5076
rect 4896 5076 4914 5094
rect 4896 5094 4914 5112
rect 4896 5112 4914 5130
rect 4896 5130 4914 5148
rect 4896 5148 4914 5166
rect 4896 5166 4914 5184
rect 4896 5184 4914 5202
rect 4896 5202 4914 5220
rect 4896 5220 4914 5238
rect 4896 5238 4914 5256
rect 4896 5256 4914 5274
rect 4896 5274 4914 5292
rect 4896 5292 4914 5310
rect 4896 5310 4914 5328
rect 4896 5328 4914 5346
rect 4896 5346 4914 5364
rect 4896 5364 4914 5382
rect 4896 5382 4914 5400
rect 4896 5400 4914 5418
rect 4896 5418 4914 5436
rect 4896 5436 4914 5454
rect 4896 5454 4914 5472
rect 4896 5472 4914 5490
rect 4896 5490 4914 5508
rect 4896 5508 4914 5526
rect 4896 5526 4914 5544
rect 4896 5544 4914 5562
rect 4896 5562 4914 5580
rect 4896 5580 4914 5598
rect 4896 5598 4914 5616
rect 4896 5616 4914 5634
rect 4896 5634 4914 5652
rect 4896 5652 4914 5670
rect 4896 5670 4914 5688
rect 4896 5688 4914 5706
rect 4896 5706 4914 5724
rect 4896 5724 4914 5742
rect 4896 5742 4914 5760
rect 4896 5760 4914 5778
rect 4896 5778 4914 5796
rect 4896 5796 4914 5814
rect 4896 5814 4914 5832
rect 4896 5832 4914 5850
rect 4896 5850 4914 5868
rect 4896 5868 4914 5886
rect 4896 5886 4914 5904
rect 4896 5904 4914 5922
rect 4896 5922 4914 5940
rect 4896 5940 4914 5958
rect 4896 5958 4914 5976
rect 4896 5976 4914 5994
rect 4896 5994 4914 6012
rect 4896 6012 4914 6030
rect 4896 6030 4914 6048
rect 4896 6048 4914 6066
rect 4896 6066 4914 6084
rect 4896 6084 4914 6102
rect 4896 6102 4914 6120
rect 4896 6120 4914 6138
rect 4896 6138 4914 6156
rect 4896 6156 4914 6174
rect 4896 6174 4914 6192
rect 4896 6192 4914 6210
rect 4896 6210 4914 6228
rect 4896 6228 4914 6246
rect 4896 6246 4914 6264
rect 4896 6264 4914 6282
rect 4896 6282 4914 6300
rect 4896 6300 4914 6318
rect 4896 6318 4914 6336
rect 4896 6336 4914 6354
rect 4896 6354 4914 6372
rect 4896 6372 4914 6390
rect 4896 6390 4914 6408
rect 4896 6408 4914 6426
rect 4896 6426 4914 6444
rect 4896 6444 4914 6462
rect 4896 6462 4914 6480
rect 4896 6480 4914 6498
rect 4896 6498 4914 6516
rect 4896 6516 4914 6534
rect 4896 6534 4914 6552
rect 4896 6552 4914 6570
rect 4896 6570 4914 6588
rect 4896 6588 4914 6606
rect 4896 6606 4914 6624
rect 4896 6624 4914 6642
rect 4896 6642 4914 6660
rect 4896 6660 4914 6678
rect 4896 6678 4914 6696
rect 4896 6696 4914 6714
rect 4896 6714 4914 6732
rect 4896 6732 4914 6750
rect 4896 6750 4914 6768
rect 4896 6768 4914 6786
rect 4896 6786 4914 6804
rect 4896 6804 4914 6822
rect 4896 6822 4914 6840
rect 4896 6840 4914 6858
rect 4896 6858 4914 6876
rect 4896 6876 4914 6894
rect 4896 6894 4914 6912
rect 4896 6912 4914 6930
rect 4896 6930 4914 6948
rect 4896 6948 4914 6966
rect 4896 6966 4914 6984
rect 4896 6984 4914 7002
rect 4896 7002 4914 7020
rect 4896 7020 4914 7038
rect 4896 7038 4914 7056
rect 4896 7056 4914 7074
rect 4896 7074 4914 7092
rect 4896 7092 4914 7110
rect 4896 7110 4914 7128
rect 4896 7128 4914 7146
rect 4896 7146 4914 7164
rect 4896 7164 4914 7182
rect 4896 7182 4914 7200
rect 4896 7200 4914 7218
rect 4896 7218 4914 7236
rect 4896 7236 4914 7254
rect 4896 7254 4914 7272
rect 4896 7272 4914 7290
rect 4896 7290 4914 7308
rect 4896 7308 4914 7326
rect 4896 7326 4914 7344
rect 4896 7344 4914 7362
rect 4896 7362 4914 7380
rect 4896 7380 4914 7398
rect 4896 7398 4914 7416
rect 4896 7416 4914 7434
rect 4896 7434 4914 7452
rect 4896 7452 4914 7470
rect 4896 7470 4914 7488
rect 4896 7488 4914 7506
rect 4896 7506 4914 7524
rect 4896 7524 4914 7542
rect 4896 7542 4914 7560
rect 4896 7560 4914 7578
rect 4896 7578 4914 7596
rect 4896 7596 4914 7614
rect 4896 7614 4914 7632
rect 4896 7632 4914 7650
rect 4896 7650 4914 7668
rect 4896 7668 4914 7686
rect 4914 234 4932 252
rect 4914 252 4932 270
rect 4914 270 4932 288
rect 4914 288 4932 306
rect 4914 306 4932 324
rect 4914 324 4932 342
rect 4914 342 4932 360
rect 4914 360 4932 378
rect 4914 378 4932 396
rect 4914 396 4932 414
rect 4914 414 4932 432
rect 4914 432 4932 450
rect 4914 450 4932 468
rect 4914 468 4932 486
rect 4914 486 4932 504
rect 4914 504 4932 522
rect 4914 522 4932 540
rect 4914 540 4932 558
rect 4914 558 4932 576
rect 4914 576 4932 594
rect 4914 594 4932 612
rect 4914 612 4932 630
rect 4914 630 4932 648
rect 4914 648 4932 666
rect 4914 666 4932 684
rect 4914 684 4932 702
rect 4914 702 4932 720
rect 4914 720 4932 738
rect 4914 738 4932 756
rect 4914 864 4932 882
rect 4914 882 4932 900
rect 4914 900 4932 918
rect 4914 918 4932 936
rect 4914 936 4932 954
rect 4914 954 4932 972
rect 4914 972 4932 990
rect 4914 990 4932 1008
rect 4914 1008 4932 1026
rect 4914 1026 4932 1044
rect 4914 1044 4932 1062
rect 4914 1062 4932 1080
rect 4914 1080 4932 1098
rect 4914 1098 4932 1116
rect 4914 1116 4932 1134
rect 4914 1134 4932 1152
rect 4914 1152 4932 1170
rect 4914 1170 4932 1188
rect 4914 1188 4932 1206
rect 4914 1206 4932 1224
rect 4914 1224 4932 1242
rect 4914 1242 4932 1260
rect 4914 1260 4932 1278
rect 4914 1278 4932 1296
rect 4914 1296 4932 1314
rect 4914 1314 4932 1332
rect 4914 1332 4932 1350
rect 4914 1350 4932 1368
rect 4914 1368 4932 1386
rect 4914 1386 4932 1404
rect 4914 1404 4932 1422
rect 4914 1422 4932 1440
rect 4914 1440 4932 1458
rect 4914 1458 4932 1476
rect 4914 1476 4932 1494
rect 4914 1494 4932 1512
rect 4914 1512 4932 1530
rect 4914 1530 4932 1548
rect 4914 1548 4932 1566
rect 4914 1566 4932 1584
rect 4914 1584 4932 1602
rect 4914 1602 4932 1620
rect 4914 1620 4932 1638
rect 4914 1638 4932 1656
rect 4914 1656 4932 1674
rect 4914 1674 4932 1692
rect 4914 1692 4932 1710
rect 4914 1710 4932 1728
rect 4914 1728 4932 1746
rect 4914 1746 4932 1764
rect 4914 1764 4932 1782
rect 4914 1782 4932 1800
rect 4914 1800 4932 1818
rect 4914 1818 4932 1836
rect 4914 1836 4932 1854
rect 4914 1854 4932 1872
rect 4914 1872 4932 1890
rect 4914 1890 4932 1908
rect 4914 1908 4932 1926
rect 4914 1926 4932 1944
rect 4914 1944 4932 1962
rect 4914 1962 4932 1980
rect 4914 1980 4932 1998
rect 4914 1998 4932 2016
rect 4914 2016 4932 2034
rect 4914 2034 4932 2052
rect 4914 2052 4932 2070
rect 4914 2070 4932 2088
rect 4914 2088 4932 2106
rect 4914 2106 4932 2124
rect 4914 2124 4932 2142
rect 4914 2142 4932 2160
rect 4914 2160 4932 2178
rect 4914 2394 4932 2412
rect 4914 2412 4932 2430
rect 4914 2430 4932 2448
rect 4914 2448 4932 2466
rect 4914 2466 4932 2484
rect 4914 2484 4932 2502
rect 4914 2502 4932 2520
rect 4914 2520 4932 2538
rect 4914 2538 4932 2556
rect 4914 2556 4932 2574
rect 4914 2574 4932 2592
rect 4914 2592 4932 2610
rect 4914 2610 4932 2628
rect 4914 2628 4932 2646
rect 4914 2646 4932 2664
rect 4914 2664 4932 2682
rect 4914 2682 4932 2700
rect 4914 2700 4932 2718
rect 4914 2718 4932 2736
rect 4914 2736 4932 2754
rect 4914 2754 4932 2772
rect 4914 2772 4932 2790
rect 4914 2790 4932 2808
rect 4914 2808 4932 2826
rect 4914 2826 4932 2844
rect 4914 2844 4932 2862
rect 4914 2862 4932 2880
rect 4914 2880 4932 2898
rect 4914 2898 4932 2916
rect 4914 2916 4932 2934
rect 4914 2934 4932 2952
rect 4914 2952 4932 2970
rect 4914 2970 4932 2988
rect 4914 2988 4932 3006
rect 4914 3006 4932 3024
rect 4914 3024 4932 3042
rect 4914 3042 4932 3060
rect 4914 3060 4932 3078
rect 4914 3078 4932 3096
rect 4914 3096 4932 3114
rect 4914 3114 4932 3132
rect 4914 3132 4932 3150
rect 4914 3150 4932 3168
rect 4914 3168 4932 3186
rect 4914 3186 4932 3204
rect 4914 3204 4932 3222
rect 4914 3222 4932 3240
rect 4914 3240 4932 3258
rect 4914 3258 4932 3276
rect 4914 3276 4932 3294
rect 4914 3294 4932 3312
rect 4914 3312 4932 3330
rect 4914 3330 4932 3348
rect 4914 3348 4932 3366
rect 4914 3366 4932 3384
rect 4914 3384 4932 3402
rect 4914 3402 4932 3420
rect 4914 3420 4932 3438
rect 4914 3438 4932 3456
rect 4914 3456 4932 3474
rect 4914 3474 4932 3492
rect 4914 3492 4932 3510
rect 4914 3510 4932 3528
rect 4914 3528 4932 3546
rect 4914 3546 4932 3564
rect 4914 3564 4932 3582
rect 4914 3582 4932 3600
rect 4914 3600 4932 3618
rect 4914 3618 4932 3636
rect 4914 3636 4932 3654
rect 4914 3654 4932 3672
rect 4914 3672 4932 3690
rect 4914 3690 4932 3708
rect 4914 3708 4932 3726
rect 4914 3726 4932 3744
rect 4914 3744 4932 3762
rect 4914 3762 4932 3780
rect 4914 3780 4932 3798
rect 4914 3798 4932 3816
rect 4914 3816 4932 3834
rect 4914 3834 4932 3852
rect 4914 3852 4932 3870
rect 4914 3870 4932 3888
rect 4914 3888 4932 3906
rect 4914 3906 4932 3924
rect 4914 3924 4932 3942
rect 4914 3942 4932 3960
rect 4914 3960 4932 3978
rect 4914 3978 4932 3996
rect 4914 3996 4932 4014
rect 4914 4014 4932 4032
rect 4914 4032 4932 4050
rect 4914 4050 4932 4068
rect 4914 4068 4932 4086
rect 4914 4086 4932 4104
rect 4914 4104 4932 4122
rect 4914 4122 4932 4140
rect 4914 4140 4932 4158
rect 4914 4158 4932 4176
rect 4914 4176 4932 4194
rect 4914 4194 4932 4212
rect 4914 4212 4932 4230
rect 4914 4230 4932 4248
rect 4914 4248 4932 4266
rect 4914 4266 4932 4284
rect 4914 4500 4932 4518
rect 4914 4518 4932 4536
rect 4914 4536 4932 4554
rect 4914 4554 4932 4572
rect 4914 4572 4932 4590
rect 4914 4590 4932 4608
rect 4914 4608 4932 4626
rect 4914 4626 4932 4644
rect 4914 4644 4932 4662
rect 4914 4662 4932 4680
rect 4914 4680 4932 4698
rect 4914 4698 4932 4716
rect 4914 4716 4932 4734
rect 4914 4734 4932 4752
rect 4914 4752 4932 4770
rect 4914 4770 4932 4788
rect 4914 4788 4932 4806
rect 4914 4806 4932 4824
rect 4914 4824 4932 4842
rect 4914 4842 4932 4860
rect 4914 4860 4932 4878
rect 4914 4878 4932 4896
rect 4914 4896 4932 4914
rect 4914 4914 4932 4932
rect 4914 4932 4932 4950
rect 4914 4950 4932 4968
rect 4914 4968 4932 4986
rect 4914 4986 4932 5004
rect 4914 5004 4932 5022
rect 4914 5022 4932 5040
rect 4914 5040 4932 5058
rect 4914 5058 4932 5076
rect 4914 5076 4932 5094
rect 4914 5094 4932 5112
rect 4914 5112 4932 5130
rect 4914 5130 4932 5148
rect 4914 5148 4932 5166
rect 4914 5166 4932 5184
rect 4914 5184 4932 5202
rect 4914 5202 4932 5220
rect 4914 5220 4932 5238
rect 4914 5238 4932 5256
rect 4914 5256 4932 5274
rect 4914 5274 4932 5292
rect 4914 5292 4932 5310
rect 4914 5310 4932 5328
rect 4914 5328 4932 5346
rect 4914 5346 4932 5364
rect 4914 5364 4932 5382
rect 4914 5382 4932 5400
rect 4914 5400 4932 5418
rect 4914 5418 4932 5436
rect 4914 5436 4932 5454
rect 4914 5454 4932 5472
rect 4914 5472 4932 5490
rect 4914 5490 4932 5508
rect 4914 5508 4932 5526
rect 4914 5526 4932 5544
rect 4914 5544 4932 5562
rect 4914 5562 4932 5580
rect 4914 5580 4932 5598
rect 4914 5598 4932 5616
rect 4914 5616 4932 5634
rect 4914 5634 4932 5652
rect 4914 5652 4932 5670
rect 4914 5670 4932 5688
rect 4914 5688 4932 5706
rect 4914 5706 4932 5724
rect 4914 5724 4932 5742
rect 4914 5742 4932 5760
rect 4914 5760 4932 5778
rect 4914 5778 4932 5796
rect 4914 5796 4932 5814
rect 4914 5814 4932 5832
rect 4914 5832 4932 5850
rect 4914 5850 4932 5868
rect 4914 5868 4932 5886
rect 4914 5886 4932 5904
rect 4914 5904 4932 5922
rect 4914 5922 4932 5940
rect 4914 5940 4932 5958
rect 4914 5958 4932 5976
rect 4914 5976 4932 5994
rect 4914 5994 4932 6012
rect 4914 6012 4932 6030
rect 4914 6030 4932 6048
rect 4914 6048 4932 6066
rect 4914 6066 4932 6084
rect 4914 6084 4932 6102
rect 4914 6102 4932 6120
rect 4914 6120 4932 6138
rect 4914 6138 4932 6156
rect 4914 6156 4932 6174
rect 4914 6174 4932 6192
rect 4914 6192 4932 6210
rect 4914 6210 4932 6228
rect 4914 6228 4932 6246
rect 4914 6246 4932 6264
rect 4914 6264 4932 6282
rect 4914 6282 4932 6300
rect 4914 6300 4932 6318
rect 4914 6318 4932 6336
rect 4914 6336 4932 6354
rect 4914 6354 4932 6372
rect 4914 6372 4932 6390
rect 4914 6390 4932 6408
rect 4914 6408 4932 6426
rect 4914 6426 4932 6444
rect 4914 6444 4932 6462
rect 4914 6462 4932 6480
rect 4914 6480 4932 6498
rect 4914 6498 4932 6516
rect 4914 6516 4932 6534
rect 4914 6534 4932 6552
rect 4914 6552 4932 6570
rect 4914 6570 4932 6588
rect 4914 6588 4932 6606
rect 4914 6606 4932 6624
rect 4914 6624 4932 6642
rect 4914 6642 4932 6660
rect 4914 6660 4932 6678
rect 4914 6678 4932 6696
rect 4914 6696 4932 6714
rect 4914 6714 4932 6732
rect 4914 6732 4932 6750
rect 4914 6750 4932 6768
rect 4914 6768 4932 6786
rect 4914 6786 4932 6804
rect 4914 6804 4932 6822
rect 4914 6822 4932 6840
rect 4914 6840 4932 6858
rect 4914 6858 4932 6876
rect 4914 6876 4932 6894
rect 4914 6894 4932 6912
rect 4914 6912 4932 6930
rect 4914 6930 4932 6948
rect 4914 6948 4932 6966
rect 4914 6966 4932 6984
rect 4914 6984 4932 7002
rect 4914 7002 4932 7020
rect 4914 7020 4932 7038
rect 4914 7038 4932 7056
rect 4914 7056 4932 7074
rect 4914 7074 4932 7092
rect 4914 7092 4932 7110
rect 4914 7110 4932 7128
rect 4914 7128 4932 7146
rect 4914 7146 4932 7164
rect 4914 7164 4932 7182
rect 4914 7182 4932 7200
rect 4914 7200 4932 7218
rect 4914 7218 4932 7236
rect 4914 7236 4932 7254
rect 4914 7254 4932 7272
rect 4914 7272 4932 7290
rect 4914 7290 4932 7308
rect 4914 7308 4932 7326
rect 4914 7326 4932 7344
rect 4914 7344 4932 7362
rect 4914 7362 4932 7380
rect 4914 7380 4932 7398
rect 4914 7398 4932 7416
rect 4914 7416 4932 7434
rect 4914 7434 4932 7452
rect 4914 7452 4932 7470
rect 4914 7470 4932 7488
rect 4914 7488 4932 7506
rect 4914 7506 4932 7524
rect 4914 7524 4932 7542
rect 4914 7542 4932 7560
rect 4914 7560 4932 7578
rect 4914 7578 4932 7596
rect 4914 7596 4932 7614
rect 4914 7614 4932 7632
rect 4914 7632 4932 7650
rect 4914 7650 4932 7668
rect 4914 7668 4932 7686
rect 4914 7686 4932 7704
rect 4914 7704 4932 7722
rect 4932 234 4950 252
rect 4932 252 4950 270
rect 4932 270 4950 288
rect 4932 288 4950 306
rect 4932 306 4950 324
rect 4932 324 4950 342
rect 4932 342 4950 360
rect 4932 360 4950 378
rect 4932 378 4950 396
rect 4932 396 4950 414
rect 4932 414 4950 432
rect 4932 432 4950 450
rect 4932 450 4950 468
rect 4932 468 4950 486
rect 4932 486 4950 504
rect 4932 504 4950 522
rect 4932 522 4950 540
rect 4932 540 4950 558
rect 4932 558 4950 576
rect 4932 576 4950 594
rect 4932 594 4950 612
rect 4932 612 4950 630
rect 4932 630 4950 648
rect 4932 648 4950 666
rect 4932 666 4950 684
rect 4932 684 4950 702
rect 4932 702 4950 720
rect 4932 720 4950 738
rect 4932 738 4950 756
rect 4932 864 4950 882
rect 4932 882 4950 900
rect 4932 900 4950 918
rect 4932 918 4950 936
rect 4932 936 4950 954
rect 4932 954 4950 972
rect 4932 972 4950 990
rect 4932 990 4950 1008
rect 4932 1008 4950 1026
rect 4932 1026 4950 1044
rect 4932 1044 4950 1062
rect 4932 1062 4950 1080
rect 4932 1080 4950 1098
rect 4932 1098 4950 1116
rect 4932 1116 4950 1134
rect 4932 1134 4950 1152
rect 4932 1152 4950 1170
rect 4932 1170 4950 1188
rect 4932 1188 4950 1206
rect 4932 1206 4950 1224
rect 4932 1224 4950 1242
rect 4932 1242 4950 1260
rect 4932 1260 4950 1278
rect 4932 1278 4950 1296
rect 4932 1296 4950 1314
rect 4932 1314 4950 1332
rect 4932 1332 4950 1350
rect 4932 1350 4950 1368
rect 4932 1368 4950 1386
rect 4932 1386 4950 1404
rect 4932 1404 4950 1422
rect 4932 1422 4950 1440
rect 4932 1440 4950 1458
rect 4932 1458 4950 1476
rect 4932 1476 4950 1494
rect 4932 1494 4950 1512
rect 4932 1512 4950 1530
rect 4932 1530 4950 1548
rect 4932 1548 4950 1566
rect 4932 1566 4950 1584
rect 4932 1584 4950 1602
rect 4932 1602 4950 1620
rect 4932 1620 4950 1638
rect 4932 1638 4950 1656
rect 4932 1656 4950 1674
rect 4932 1674 4950 1692
rect 4932 1692 4950 1710
rect 4932 1710 4950 1728
rect 4932 1728 4950 1746
rect 4932 1746 4950 1764
rect 4932 1764 4950 1782
rect 4932 1782 4950 1800
rect 4932 1800 4950 1818
rect 4932 1818 4950 1836
rect 4932 1836 4950 1854
rect 4932 1854 4950 1872
rect 4932 1872 4950 1890
rect 4932 1890 4950 1908
rect 4932 1908 4950 1926
rect 4932 1926 4950 1944
rect 4932 1944 4950 1962
rect 4932 1962 4950 1980
rect 4932 1980 4950 1998
rect 4932 1998 4950 2016
rect 4932 2016 4950 2034
rect 4932 2034 4950 2052
rect 4932 2052 4950 2070
rect 4932 2070 4950 2088
rect 4932 2088 4950 2106
rect 4932 2106 4950 2124
rect 4932 2124 4950 2142
rect 4932 2142 4950 2160
rect 4932 2160 4950 2178
rect 4932 2412 4950 2430
rect 4932 2430 4950 2448
rect 4932 2448 4950 2466
rect 4932 2466 4950 2484
rect 4932 2484 4950 2502
rect 4932 2502 4950 2520
rect 4932 2520 4950 2538
rect 4932 2538 4950 2556
rect 4932 2556 4950 2574
rect 4932 2574 4950 2592
rect 4932 2592 4950 2610
rect 4932 2610 4950 2628
rect 4932 2628 4950 2646
rect 4932 2646 4950 2664
rect 4932 2664 4950 2682
rect 4932 2682 4950 2700
rect 4932 2700 4950 2718
rect 4932 2718 4950 2736
rect 4932 2736 4950 2754
rect 4932 2754 4950 2772
rect 4932 2772 4950 2790
rect 4932 2790 4950 2808
rect 4932 2808 4950 2826
rect 4932 2826 4950 2844
rect 4932 2844 4950 2862
rect 4932 2862 4950 2880
rect 4932 2880 4950 2898
rect 4932 2898 4950 2916
rect 4932 2916 4950 2934
rect 4932 2934 4950 2952
rect 4932 2952 4950 2970
rect 4932 2970 4950 2988
rect 4932 2988 4950 3006
rect 4932 3006 4950 3024
rect 4932 3024 4950 3042
rect 4932 3042 4950 3060
rect 4932 3060 4950 3078
rect 4932 3078 4950 3096
rect 4932 3096 4950 3114
rect 4932 3114 4950 3132
rect 4932 3132 4950 3150
rect 4932 3150 4950 3168
rect 4932 3168 4950 3186
rect 4932 3186 4950 3204
rect 4932 3204 4950 3222
rect 4932 3222 4950 3240
rect 4932 3240 4950 3258
rect 4932 3258 4950 3276
rect 4932 3276 4950 3294
rect 4932 3294 4950 3312
rect 4932 3312 4950 3330
rect 4932 3330 4950 3348
rect 4932 3348 4950 3366
rect 4932 3366 4950 3384
rect 4932 3384 4950 3402
rect 4932 3402 4950 3420
rect 4932 3420 4950 3438
rect 4932 3438 4950 3456
rect 4932 3456 4950 3474
rect 4932 3474 4950 3492
rect 4932 3492 4950 3510
rect 4932 3510 4950 3528
rect 4932 3528 4950 3546
rect 4932 3546 4950 3564
rect 4932 3564 4950 3582
rect 4932 3582 4950 3600
rect 4932 3600 4950 3618
rect 4932 3618 4950 3636
rect 4932 3636 4950 3654
rect 4932 3654 4950 3672
rect 4932 3672 4950 3690
rect 4932 3690 4950 3708
rect 4932 3708 4950 3726
rect 4932 3726 4950 3744
rect 4932 3744 4950 3762
rect 4932 3762 4950 3780
rect 4932 3780 4950 3798
rect 4932 3798 4950 3816
rect 4932 3816 4950 3834
rect 4932 3834 4950 3852
rect 4932 3852 4950 3870
rect 4932 3870 4950 3888
rect 4932 3888 4950 3906
rect 4932 3906 4950 3924
rect 4932 3924 4950 3942
rect 4932 3942 4950 3960
rect 4932 3960 4950 3978
rect 4932 3978 4950 3996
rect 4932 3996 4950 4014
rect 4932 4014 4950 4032
rect 4932 4032 4950 4050
rect 4932 4050 4950 4068
rect 4932 4068 4950 4086
rect 4932 4086 4950 4104
rect 4932 4104 4950 4122
rect 4932 4122 4950 4140
rect 4932 4140 4950 4158
rect 4932 4158 4950 4176
rect 4932 4176 4950 4194
rect 4932 4194 4950 4212
rect 4932 4212 4950 4230
rect 4932 4230 4950 4248
rect 4932 4248 4950 4266
rect 4932 4266 4950 4284
rect 4932 4284 4950 4302
rect 4932 4518 4950 4536
rect 4932 4536 4950 4554
rect 4932 4554 4950 4572
rect 4932 4572 4950 4590
rect 4932 4590 4950 4608
rect 4932 4608 4950 4626
rect 4932 4626 4950 4644
rect 4932 4644 4950 4662
rect 4932 4662 4950 4680
rect 4932 4680 4950 4698
rect 4932 4698 4950 4716
rect 4932 4716 4950 4734
rect 4932 4734 4950 4752
rect 4932 4752 4950 4770
rect 4932 4770 4950 4788
rect 4932 4788 4950 4806
rect 4932 4806 4950 4824
rect 4932 4824 4950 4842
rect 4932 4842 4950 4860
rect 4932 4860 4950 4878
rect 4932 4878 4950 4896
rect 4932 4896 4950 4914
rect 4932 4914 4950 4932
rect 4932 4932 4950 4950
rect 4932 4950 4950 4968
rect 4932 4968 4950 4986
rect 4932 4986 4950 5004
rect 4932 5004 4950 5022
rect 4932 5022 4950 5040
rect 4932 5040 4950 5058
rect 4932 5058 4950 5076
rect 4932 5076 4950 5094
rect 4932 5094 4950 5112
rect 4932 5112 4950 5130
rect 4932 5130 4950 5148
rect 4932 5148 4950 5166
rect 4932 5166 4950 5184
rect 4932 5184 4950 5202
rect 4932 5202 4950 5220
rect 4932 5220 4950 5238
rect 4932 5238 4950 5256
rect 4932 5256 4950 5274
rect 4932 5274 4950 5292
rect 4932 5292 4950 5310
rect 4932 5310 4950 5328
rect 4932 5328 4950 5346
rect 4932 5346 4950 5364
rect 4932 5364 4950 5382
rect 4932 5382 4950 5400
rect 4932 5400 4950 5418
rect 4932 5418 4950 5436
rect 4932 5436 4950 5454
rect 4932 5454 4950 5472
rect 4932 5472 4950 5490
rect 4932 5490 4950 5508
rect 4932 5508 4950 5526
rect 4932 5526 4950 5544
rect 4932 5544 4950 5562
rect 4932 5562 4950 5580
rect 4932 5580 4950 5598
rect 4932 5598 4950 5616
rect 4932 5616 4950 5634
rect 4932 5634 4950 5652
rect 4932 5652 4950 5670
rect 4932 5670 4950 5688
rect 4932 5688 4950 5706
rect 4932 5706 4950 5724
rect 4932 5724 4950 5742
rect 4932 5742 4950 5760
rect 4932 5760 4950 5778
rect 4932 5778 4950 5796
rect 4932 5796 4950 5814
rect 4932 5814 4950 5832
rect 4932 5832 4950 5850
rect 4932 5850 4950 5868
rect 4932 5868 4950 5886
rect 4932 5886 4950 5904
rect 4932 5904 4950 5922
rect 4932 5922 4950 5940
rect 4932 5940 4950 5958
rect 4932 5958 4950 5976
rect 4932 5976 4950 5994
rect 4932 5994 4950 6012
rect 4932 6012 4950 6030
rect 4932 6030 4950 6048
rect 4932 6048 4950 6066
rect 4932 6066 4950 6084
rect 4932 6084 4950 6102
rect 4932 6102 4950 6120
rect 4932 6120 4950 6138
rect 4932 6138 4950 6156
rect 4932 6156 4950 6174
rect 4932 6174 4950 6192
rect 4932 6192 4950 6210
rect 4932 6210 4950 6228
rect 4932 6228 4950 6246
rect 4932 6246 4950 6264
rect 4932 6264 4950 6282
rect 4932 6282 4950 6300
rect 4932 6300 4950 6318
rect 4932 6318 4950 6336
rect 4932 6336 4950 6354
rect 4932 6354 4950 6372
rect 4932 6372 4950 6390
rect 4932 6390 4950 6408
rect 4932 6408 4950 6426
rect 4932 6426 4950 6444
rect 4932 6444 4950 6462
rect 4932 6462 4950 6480
rect 4932 6480 4950 6498
rect 4932 6498 4950 6516
rect 4932 6516 4950 6534
rect 4932 6534 4950 6552
rect 4932 6552 4950 6570
rect 4932 6570 4950 6588
rect 4932 6588 4950 6606
rect 4932 6606 4950 6624
rect 4932 6624 4950 6642
rect 4932 6642 4950 6660
rect 4932 6660 4950 6678
rect 4932 6678 4950 6696
rect 4932 6696 4950 6714
rect 4932 6714 4950 6732
rect 4932 6732 4950 6750
rect 4932 6750 4950 6768
rect 4932 6768 4950 6786
rect 4932 6786 4950 6804
rect 4932 6804 4950 6822
rect 4932 6822 4950 6840
rect 4932 6840 4950 6858
rect 4932 6858 4950 6876
rect 4932 6876 4950 6894
rect 4932 6894 4950 6912
rect 4932 6912 4950 6930
rect 4932 6930 4950 6948
rect 4932 6948 4950 6966
rect 4932 6966 4950 6984
rect 4932 6984 4950 7002
rect 4932 7002 4950 7020
rect 4932 7020 4950 7038
rect 4932 7038 4950 7056
rect 4932 7056 4950 7074
rect 4932 7074 4950 7092
rect 4932 7092 4950 7110
rect 4932 7110 4950 7128
rect 4932 7128 4950 7146
rect 4932 7146 4950 7164
rect 4932 7164 4950 7182
rect 4932 7182 4950 7200
rect 4932 7200 4950 7218
rect 4932 7218 4950 7236
rect 4932 7236 4950 7254
rect 4932 7254 4950 7272
rect 4932 7272 4950 7290
rect 4932 7290 4950 7308
rect 4932 7308 4950 7326
rect 4932 7326 4950 7344
rect 4932 7344 4950 7362
rect 4932 7362 4950 7380
rect 4932 7380 4950 7398
rect 4932 7398 4950 7416
rect 4932 7416 4950 7434
rect 4932 7434 4950 7452
rect 4932 7452 4950 7470
rect 4932 7470 4950 7488
rect 4932 7488 4950 7506
rect 4932 7506 4950 7524
rect 4932 7524 4950 7542
rect 4932 7542 4950 7560
rect 4932 7560 4950 7578
rect 4932 7578 4950 7596
rect 4932 7596 4950 7614
rect 4932 7614 4950 7632
rect 4932 7632 4950 7650
rect 4932 7650 4950 7668
rect 4932 7668 4950 7686
rect 4932 7686 4950 7704
rect 4932 7704 4950 7722
rect 4932 7722 4950 7740
rect 4950 252 4968 270
rect 4950 270 4968 288
rect 4950 288 4968 306
rect 4950 306 4968 324
rect 4950 324 4968 342
rect 4950 342 4968 360
rect 4950 360 4968 378
rect 4950 378 4968 396
rect 4950 396 4968 414
rect 4950 414 4968 432
rect 4950 432 4968 450
rect 4950 450 4968 468
rect 4950 468 4968 486
rect 4950 486 4968 504
rect 4950 504 4968 522
rect 4950 522 4968 540
rect 4950 540 4968 558
rect 4950 558 4968 576
rect 4950 576 4968 594
rect 4950 594 4968 612
rect 4950 612 4968 630
rect 4950 630 4968 648
rect 4950 648 4968 666
rect 4950 666 4968 684
rect 4950 684 4968 702
rect 4950 702 4968 720
rect 4950 720 4968 738
rect 4950 738 4968 756
rect 4950 864 4968 882
rect 4950 882 4968 900
rect 4950 900 4968 918
rect 4950 918 4968 936
rect 4950 936 4968 954
rect 4950 954 4968 972
rect 4950 972 4968 990
rect 4950 990 4968 1008
rect 4950 1008 4968 1026
rect 4950 1026 4968 1044
rect 4950 1044 4968 1062
rect 4950 1062 4968 1080
rect 4950 1080 4968 1098
rect 4950 1098 4968 1116
rect 4950 1116 4968 1134
rect 4950 1134 4968 1152
rect 4950 1152 4968 1170
rect 4950 1170 4968 1188
rect 4950 1188 4968 1206
rect 4950 1206 4968 1224
rect 4950 1224 4968 1242
rect 4950 1242 4968 1260
rect 4950 1260 4968 1278
rect 4950 1278 4968 1296
rect 4950 1296 4968 1314
rect 4950 1314 4968 1332
rect 4950 1332 4968 1350
rect 4950 1350 4968 1368
rect 4950 1368 4968 1386
rect 4950 1386 4968 1404
rect 4950 1404 4968 1422
rect 4950 1422 4968 1440
rect 4950 1440 4968 1458
rect 4950 1458 4968 1476
rect 4950 1476 4968 1494
rect 4950 1494 4968 1512
rect 4950 1512 4968 1530
rect 4950 1530 4968 1548
rect 4950 1548 4968 1566
rect 4950 1566 4968 1584
rect 4950 1584 4968 1602
rect 4950 1602 4968 1620
rect 4950 1620 4968 1638
rect 4950 1638 4968 1656
rect 4950 1656 4968 1674
rect 4950 1674 4968 1692
rect 4950 1692 4968 1710
rect 4950 1710 4968 1728
rect 4950 1728 4968 1746
rect 4950 1746 4968 1764
rect 4950 1764 4968 1782
rect 4950 1782 4968 1800
rect 4950 1800 4968 1818
rect 4950 1818 4968 1836
rect 4950 1836 4968 1854
rect 4950 1854 4968 1872
rect 4950 1872 4968 1890
rect 4950 1890 4968 1908
rect 4950 1908 4968 1926
rect 4950 1926 4968 1944
rect 4950 1944 4968 1962
rect 4950 1962 4968 1980
rect 4950 1980 4968 1998
rect 4950 1998 4968 2016
rect 4950 2016 4968 2034
rect 4950 2034 4968 2052
rect 4950 2052 4968 2070
rect 4950 2070 4968 2088
rect 4950 2088 4968 2106
rect 4950 2106 4968 2124
rect 4950 2124 4968 2142
rect 4950 2142 4968 2160
rect 4950 2160 4968 2178
rect 4950 2178 4968 2196
rect 4950 2412 4968 2430
rect 4950 2430 4968 2448
rect 4950 2448 4968 2466
rect 4950 2466 4968 2484
rect 4950 2484 4968 2502
rect 4950 2502 4968 2520
rect 4950 2520 4968 2538
rect 4950 2538 4968 2556
rect 4950 2556 4968 2574
rect 4950 2574 4968 2592
rect 4950 2592 4968 2610
rect 4950 2610 4968 2628
rect 4950 2628 4968 2646
rect 4950 2646 4968 2664
rect 4950 2664 4968 2682
rect 4950 2682 4968 2700
rect 4950 2700 4968 2718
rect 4950 2718 4968 2736
rect 4950 2736 4968 2754
rect 4950 2754 4968 2772
rect 4950 2772 4968 2790
rect 4950 2790 4968 2808
rect 4950 2808 4968 2826
rect 4950 2826 4968 2844
rect 4950 2844 4968 2862
rect 4950 2862 4968 2880
rect 4950 2880 4968 2898
rect 4950 2898 4968 2916
rect 4950 2916 4968 2934
rect 4950 2934 4968 2952
rect 4950 2952 4968 2970
rect 4950 2970 4968 2988
rect 4950 2988 4968 3006
rect 4950 3006 4968 3024
rect 4950 3024 4968 3042
rect 4950 3042 4968 3060
rect 4950 3060 4968 3078
rect 4950 3078 4968 3096
rect 4950 3096 4968 3114
rect 4950 3114 4968 3132
rect 4950 3132 4968 3150
rect 4950 3150 4968 3168
rect 4950 3168 4968 3186
rect 4950 3186 4968 3204
rect 4950 3204 4968 3222
rect 4950 3222 4968 3240
rect 4950 3240 4968 3258
rect 4950 3258 4968 3276
rect 4950 3276 4968 3294
rect 4950 3294 4968 3312
rect 4950 3312 4968 3330
rect 4950 3330 4968 3348
rect 4950 3348 4968 3366
rect 4950 3366 4968 3384
rect 4950 3384 4968 3402
rect 4950 3402 4968 3420
rect 4950 3420 4968 3438
rect 4950 3438 4968 3456
rect 4950 3456 4968 3474
rect 4950 3474 4968 3492
rect 4950 3492 4968 3510
rect 4950 3510 4968 3528
rect 4950 3528 4968 3546
rect 4950 3546 4968 3564
rect 4950 3564 4968 3582
rect 4950 3582 4968 3600
rect 4950 3600 4968 3618
rect 4950 3618 4968 3636
rect 4950 3636 4968 3654
rect 4950 3654 4968 3672
rect 4950 3672 4968 3690
rect 4950 3690 4968 3708
rect 4950 3708 4968 3726
rect 4950 3726 4968 3744
rect 4950 3744 4968 3762
rect 4950 3762 4968 3780
rect 4950 3780 4968 3798
rect 4950 3798 4968 3816
rect 4950 3816 4968 3834
rect 4950 3834 4968 3852
rect 4950 3852 4968 3870
rect 4950 3870 4968 3888
rect 4950 3888 4968 3906
rect 4950 3906 4968 3924
rect 4950 3924 4968 3942
rect 4950 3942 4968 3960
rect 4950 3960 4968 3978
rect 4950 3978 4968 3996
rect 4950 3996 4968 4014
rect 4950 4014 4968 4032
rect 4950 4032 4968 4050
rect 4950 4050 4968 4068
rect 4950 4068 4968 4086
rect 4950 4086 4968 4104
rect 4950 4104 4968 4122
rect 4950 4122 4968 4140
rect 4950 4140 4968 4158
rect 4950 4158 4968 4176
rect 4950 4176 4968 4194
rect 4950 4194 4968 4212
rect 4950 4212 4968 4230
rect 4950 4230 4968 4248
rect 4950 4248 4968 4266
rect 4950 4266 4968 4284
rect 4950 4284 4968 4302
rect 4950 4302 4968 4320
rect 4950 4320 4968 4338
rect 4950 4536 4968 4554
rect 4950 4554 4968 4572
rect 4950 4572 4968 4590
rect 4950 4590 4968 4608
rect 4950 4608 4968 4626
rect 4950 4626 4968 4644
rect 4950 4644 4968 4662
rect 4950 4662 4968 4680
rect 4950 4680 4968 4698
rect 4950 4698 4968 4716
rect 4950 4716 4968 4734
rect 4950 4734 4968 4752
rect 4950 4752 4968 4770
rect 4950 4770 4968 4788
rect 4950 4788 4968 4806
rect 4950 4806 4968 4824
rect 4950 4824 4968 4842
rect 4950 4842 4968 4860
rect 4950 4860 4968 4878
rect 4950 4878 4968 4896
rect 4950 4896 4968 4914
rect 4950 4914 4968 4932
rect 4950 4932 4968 4950
rect 4950 4950 4968 4968
rect 4950 4968 4968 4986
rect 4950 4986 4968 5004
rect 4950 5004 4968 5022
rect 4950 5022 4968 5040
rect 4950 5040 4968 5058
rect 4950 5058 4968 5076
rect 4950 5076 4968 5094
rect 4950 5094 4968 5112
rect 4950 5112 4968 5130
rect 4950 5130 4968 5148
rect 4950 5148 4968 5166
rect 4950 5166 4968 5184
rect 4950 5184 4968 5202
rect 4950 5202 4968 5220
rect 4950 5220 4968 5238
rect 4950 5238 4968 5256
rect 4950 5256 4968 5274
rect 4950 5274 4968 5292
rect 4950 5292 4968 5310
rect 4950 5310 4968 5328
rect 4950 5328 4968 5346
rect 4950 5346 4968 5364
rect 4950 5364 4968 5382
rect 4950 5382 4968 5400
rect 4950 5400 4968 5418
rect 4950 5418 4968 5436
rect 4950 5436 4968 5454
rect 4950 5454 4968 5472
rect 4950 5472 4968 5490
rect 4950 5490 4968 5508
rect 4950 5508 4968 5526
rect 4950 5526 4968 5544
rect 4950 5544 4968 5562
rect 4950 5562 4968 5580
rect 4950 5580 4968 5598
rect 4950 5598 4968 5616
rect 4950 5616 4968 5634
rect 4950 5634 4968 5652
rect 4950 5652 4968 5670
rect 4950 5670 4968 5688
rect 4950 5688 4968 5706
rect 4950 5706 4968 5724
rect 4950 5724 4968 5742
rect 4950 5742 4968 5760
rect 4950 5760 4968 5778
rect 4950 5778 4968 5796
rect 4950 5796 4968 5814
rect 4950 5814 4968 5832
rect 4950 5832 4968 5850
rect 4950 5850 4968 5868
rect 4950 5868 4968 5886
rect 4950 5886 4968 5904
rect 4950 5904 4968 5922
rect 4950 5922 4968 5940
rect 4950 5940 4968 5958
rect 4950 5958 4968 5976
rect 4950 5976 4968 5994
rect 4950 5994 4968 6012
rect 4950 6012 4968 6030
rect 4950 6030 4968 6048
rect 4950 6048 4968 6066
rect 4950 6066 4968 6084
rect 4950 6084 4968 6102
rect 4950 6102 4968 6120
rect 4950 6120 4968 6138
rect 4950 6138 4968 6156
rect 4950 6156 4968 6174
rect 4950 6174 4968 6192
rect 4950 6192 4968 6210
rect 4950 6210 4968 6228
rect 4950 6228 4968 6246
rect 4950 6246 4968 6264
rect 4950 6264 4968 6282
rect 4950 6282 4968 6300
rect 4950 6300 4968 6318
rect 4950 6318 4968 6336
rect 4950 6336 4968 6354
rect 4950 6354 4968 6372
rect 4950 6372 4968 6390
rect 4950 6390 4968 6408
rect 4950 6408 4968 6426
rect 4950 6426 4968 6444
rect 4950 6444 4968 6462
rect 4950 6462 4968 6480
rect 4950 6480 4968 6498
rect 4950 6498 4968 6516
rect 4950 6516 4968 6534
rect 4950 6534 4968 6552
rect 4950 6552 4968 6570
rect 4950 6570 4968 6588
rect 4950 6588 4968 6606
rect 4950 6606 4968 6624
rect 4950 6624 4968 6642
rect 4950 6642 4968 6660
rect 4950 6660 4968 6678
rect 4950 6678 4968 6696
rect 4950 6696 4968 6714
rect 4950 6714 4968 6732
rect 4950 6732 4968 6750
rect 4950 6750 4968 6768
rect 4950 6768 4968 6786
rect 4950 6786 4968 6804
rect 4950 6804 4968 6822
rect 4950 6822 4968 6840
rect 4950 6840 4968 6858
rect 4950 6858 4968 6876
rect 4950 6876 4968 6894
rect 4950 6894 4968 6912
rect 4950 6912 4968 6930
rect 4950 6930 4968 6948
rect 4950 6948 4968 6966
rect 4950 6966 4968 6984
rect 4950 6984 4968 7002
rect 4950 7002 4968 7020
rect 4950 7020 4968 7038
rect 4950 7038 4968 7056
rect 4950 7056 4968 7074
rect 4950 7074 4968 7092
rect 4950 7092 4968 7110
rect 4950 7110 4968 7128
rect 4950 7128 4968 7146
rect 4950 7146 4968 7164
rect 4950 7164 4968 7182
rect 4950 7182 4968 7200
rect 4950 7200 4968 7218
rect 4950 7218 4968 7236
rect 4950 7236 4968 7254
rect 4950 7254 4968 7272
rect 4950 7272 4968 7290
rect 4950 7290 4968 7308
rect 4950 7308 4968 7326
rect 4950 7326 4968 7344
rect 4950 7344 4968 7362
rect 4950 7362 4968 7380
rect 4950 7380 4968 7398
rect 4950 7398 4968 7416
rect 4950 7416 4968 7434
rect 4950 7434 4968 7452
rect 4950 7452 4968 7470
rect 4950 7470 4968 7488
rect 4950 7488 4968 7506
rect 4950 7506 4968 7524
rect 4950 7524 4968 7542
rect 4950 7542 4968 7560
rect 4950 7560 4968 7578
rect 4950 7578 4968 7596
rect 4950 7596 4968 7614
rect 4950 7614 4968 7632
rect 4950 7632 4968 7650
rect 4950 7650 4968 7668
rect 4950 7668 4968 7686
rect 4950 7686 4968 7704
rect 4950 7704 4968 7722
rect 4950 7722 4968 7740
rect 4950 7740 4968 7758
rect 4950 7758 4968 7776
rect 4968 252 4986 270
rect 4968 270 4986 288
rect 4968 288 4986 306
rect 4968 306 4986 324
rect 4968 324 4986 342
rect 4968 342 4986 360
rect 4968 360 4986 378
rect 4968 378 4986 396
rect 4968 396 4986 414
rect 4968 414 4986 432
rect 4968 432 4986 450
rect 4968 450 4986 468
rect 4968 468 4986 486
rect 4968 486 4986 504
rect 4968 504 4986 522
rect 4968 522 4986 540
rect 4968 540 4986 558
rect 4968 558 4986 576
rect 4968 576 4986 594
rect 4968 594 4986 612
rect 4968 612 4986 630
rect 4968 630 4986 648
rect 4968 648 4986 666
rect 4968 666 4986 684
rect 4968 684 4986 702
rect 4968 702 4986 720
rect 4968 720 4986 738
rect 4968 738 4986 756
rect 4968 864 4986 882
rect 4968 882 4986 900
rect 4968 900 4986 918
rect 4968 918 4986 936
rect 4968 936 4986 954
rect 4968 954 4986 972
rect 4968 972 4986 990
rect 4968 990 4986 1008
rect 4968 1008 4986 1026
rect 4968 1026 4986 1044
rect 4968 1044 4986 1062
rect 4968 1062 4986 1080
rect 4968 1080 4986 1098
rect 4968 1098 4986 1116
rect 4968 1116 4986 1134
rect 4968 1134 4986 1152
rect 4968 1152 4986 1170
rect 4968 1170 4986 1188
rect 4968 1188 4986 1206
rect 4968 1206 4986 1224
rect 4968 1224 4986 1242
rect 4968 1242 4986 1260
rect 4968 1260 4986 1278
rect 4968 1278 4986 1296
rect 4968 1296 4986 1314
rect 4968 1314 4986 1332
rect 4968 1332 4986 1350
rect 4968 1350 4986 1368
rect 4968 1368 4986 1386
rect 4968 1386 4986 1404
rect 4968 1404 4986 1422
rect 4968 1422 4986 1440
rect 4968 1440 4986 1458
rect 4968 1458 4986 1476
rect 4968 1476 4986 1494
rect 4968 1494 4986 1512
rect 4968 1512 4986 1530
rect 4968 1530 4986 1548
rect 4968 1548 4986 1566
rect 4968 1566 4986 1584
rect 4968 1584 4986 1602
rect 4968 1602 4986 1620
rect 4968 1620 4986 1638
rect 4968 1638 4986 1656
rect 4968 1656 4986 1674
rect 4968 1674 4986 1692
rect 4968 1692 4986 1710
rect 4968 1710 4986 1728
rect 4968 1728 4986 1746
rect 4968 1746 4986 1764
rect 4968 1764 4986 1782
rect 4968 1782 4986 1800
rect 4968 1800 4986 1818
rect 4968 1818 4986 1836
rect 4968 1836 4986 1854
rect 4968 1854 4986 1872
rect 4968 1872 4986 1890
rect 4968 1890 4986 1908
rect 4968 1908 4986 1926
rect 4968 1926 4986 1944
rect 4968 1944 4986 1962
rect 4968 1962 4986 1980
rect 4968 1980 4986 1998
rect 4968 1998 4986 2016
rect 4968 2016 4986 2034
rect 4968 2034 4986 2052
rect 4968 2052 4986 2070
rect 4968 2070 4986 2088
rect 4968 2088 4986 2106
rect 4968 2106 4986 2124
rect 4968 2124 4986 2142
rect 4968 2142 4986 2160
rect 4968 2160 4986 2178
rect 4968 2178 4986 2196
rect 4968 2196 4986 2214
rect 4968 2430 4986 2448
rect 4968 2448 4986 2466
rect 4968 2466 4986 2484
rect 4968 2484 4986 2502
rect 4968 2502 4986 2520
rect 4968 2520 4986 2538
rect 4968 2538 4986 2556
rect 4968 2556 4986 2574
rect 4968 2574 4986 2592
rect 4968 2592 4986 2610
rect 4968 2610 4986 2628
rect 4968 2628 4986 2646
rect 4968 2646 4986 2664
rect 4968 2664 4986 2682
rect 4968 2682 4986 2700
rect 4968 2700 4986 2718
rect 4968 2718 4986 2736
rect 4968 2736 4986 2754
rect 4968 2754 4986 2772
rect 4968 2772 4986 2790
rect 4968 2790 4986 2808
rect 4968 2808 4986 2826
rect 4968 2826 4986 2844
rect 4968 2844 4986 2862
rect 4968 2862 4986 2880
rect 4968 2880 4986 2898
rect 4968 2898 4986 2916
rect 4968 2916 4986 2934
rect 4968 2934 4986 2952
rect 4968 2952 4986 2970
rect 4968 2970 4986 2988
rect 4968 2988 4986 3006
rect 4968 3006 4986 3024
rect 4968 3024 4986 3042
rect 4968 3042 4986 3060
rect 4968 3060 4986 3078
rect 4968 3078 4986 3096
rect 4968 3096 4986 3114
rect 4968 3114 4986 3132
rect 4968 3132 4986 3150
rect 4968 3150 4986 3168
rect 4968 3168 4986 3186
rect 4968 3186 4986 3204
rect 4968 3204 4986 3222
rect 4968 3222 4986 3240
rect 4968 3240 4986 3258
rect 4968 3258 4986 3276
rect 4968 3276 4986 3294
rect 4968 3294 4986 3312
rect 4968 3312 4986 3330
rect 4968 3330 4986 3348
rect 4968 3348 4986 3366
rect 4968 3366 4986 3384
rect 4968 3384 4986 3402
rect 4968 3402 4986 3420
rect 4968 3420 4986 3438
rect 4968 3438 4986 3456
rect 4968 3456 4986 3474
rect 4968 3474 4986 3492
rect 4968 3492 4986 3510
rect 4968 3510 4986 3528
rect 4968 3528 4986 3546
rect 4968 3546 4986 3564
rect 4968 3564 4986 3582
rect 4968 3582 4986 3600
rect 4968 3600 4986 3618
rect 4968 3618 4986 3636
rect 4968 3636 4986 3654
rect 4968 3654 4986 3672
rect 4968 3672 4986 3690
rect 4968 3690 4986 3708
rect 4968 3708 4986 3726
rect 4968 3726 4986 3744
rect 4968 3744 4986 3762
rect 4968 3762 4986 3780
rect 4968 3780 4986 3798
rect 4968 3798 4986 3816
rect 4968 3816 4986 3834
rect 4968 3834 4986 3852
rect 4968 3852 4986 3870
rect 4968 3870 4986 3888
rect 4968 3888 4986 3906
rect 4968 3906 4986 3924
rect 4968 3924 4986 3942
rect 4968 3942 4986 3960
rect 4968 3960 4986 3978
rect 4968 3978 4986 3996
rect 4968 3996 4986 4014
rect 4968 4014 4986 4032
rect 4968 4032 4986 4050
rect 4968 4050 4986 4068
rect 4968 4068 4986 4086
rect 4968 4086 4986 4104
rect 4968 4104 4986 4122
rect 4968 4122 4986 4140
rect 4968 4140 4986 4158
rect 4968 4158 4986 4176
rect 4968 4176 4986 4194
rect 4968 4194 4986 4212
rect 4968 4212 4986 4230
rect 4968 4230 4986 4248
rect 4968 4248 4986 4266
rect 4968 4266 4986 4284
rect 4968 4284 4986 4302
rect 4968 4302 4986 4320
rect 4968 4320 4986 4338
rect 4968 4338 4986 4356
rect 4968 4554 4986 4572
rect 4968 4572 4986 4590
rect 4968 4590 4986 4608
rect 4968 4608 4986 4626
rect 4968 4626 4986 4644
rect 4968 4644 4986 4662
rect 4968 4662 4986 4680
rect 4968 4680 4986 4698
rect 4968 4698 4986 4716
rect 4968 4716 4986 4734
rect 4968 4734 4986 4752
rect 4968 4752 4986 4770
rect 4968 4770 4986 4788
rect 4968 4788 4986 4806
rect 4968 4806 4986 4824
rect 4968 4824 4986 4842
rect 4968 4842 4986 4860
rect 4968 4860 4986 4878
rect 4968 4878 4986 4896
rect 4968 4896 4986 4914
rect 4968 4914 4986 4932
rect 4968 4932 4986 4950
rect 4968 4950 4986 4968
rect 4968 4968 4986 4986
rect 4968 4986 4986 5004
rect 4968 5004 4986 5022
rect 4968 5022 4986 5040
rect 4968 5040 4986 5058
rect 4968 5058 4986 5076
rect 4968 5076 4986 5094
rect 4968 5094 4986 5112
rect 4968 5112 4986 5130
rect 4968 5130 4986 5148
rect 4968 5148 4986 5166
rect 4968 5166 4986 5184
rect 4968 5184 4986 5202
rect 4968 5202 4986 5220
rect 4968 5220 4986 5238
rect 4968 5238 4986 5256
rect 4968 5256 4986 5274
rect 4968 5274 4986 5292
rect 4968 5292 4986 5310
rect 4968 5310 4986 5328
rect 4968 5328 4986 5346
rect 4968 5346 4986 5364
rect 4968 5364 4986 5382
rect 4968 5382 4986 5400
rect 4968 5400 4986 5418
rect 4968 5418 4986 5436
rect 4968 5436 4986 5454
rect 4968 5454 4986 5472
rect 4968 5472 4986 5490
rect 4968 5490 4986 5508
rect 4968 5508 4986 5526
rect 4968 5526 4986 5544
rect 4968 5544 4986 5562
rect 4968 5562 4986 5580
rect 4968 5580 4986 5598
rect 4968 5598 4986 5616
rect 4968 5616 4986 5634
rect 4968 5634 4986 5652
rect 4968 5652 4986 5670
rect 4968 5670 4986 5688
rect 4968 5688 4986 5706
rect 4968 5706 4986 5724
rect 4968 5724 4986 5742
rect 4968 5742 4986 5760
rect 4968 5760 4986 5778
rect 4968 5778 4986 5796
rect 4968 5796 4986 5814
rect 4968 5814 4986 5832
rect 4968 5832 4986 5850
rect 4968 5850 4986 5868
rect 4968 5868 4986 5886
rect 4968 5886 4986 5904
rect 4968 5904 4986 5922
rect 4968 5922 4986 5940
rect 4968 5940 4986 5958
rect 4968 5958 4986 5976
rect 4968 5976 4986 5994
rect 4968 5994 4986 6012
rect 4968 6012 4986 6030
rect 4968 6030 4986 6048
rect 4968 6048 4986 6066
rect 4968 6066 4986 6084
rect 4968 6084 4986 6102
rect 4968 6102 4986 6120
rect 4968 6120 4986 6138
rect 4968 6138 4986 6156
rect 4968 6156 4986 6174
rect 4968 6174 4986 6192
rect 4968 6192 4986 6210
rect 4968 6210 4986 6228
rect 4968 6228 4986 6246
rect 4968 6246 4986 6264
rect 4968 6264 4986 6282
rect 4968 6282 4986 6300
rect 4968 6300 4986 6318
rect 4968 6318 4986 6336
rect 4968 6336 4986 6354
rect 4968 6354 4986 6372
rect 4968 6372 4986 6390
rect 4968 6390 4986 6408
rect 4968 6408 4986 6426
rect 4968 6426 4986 6444
rect 4968 6444 4986 6462
rect 4968 6462 4986 6480
rect 4968 6480 4986 6498
rect 4968 6498 4986 6516
rect 4968 6516 4986 6534
rect 4968 6534 4986 6552
rect 4968 6552 4986 6570
rect 4968 6570 4986 6588
rect 4968 6588 4986 6606
rect 4968 6606 4986 6624
rect 4968 6624 4986 6642
rect 4968 6642 4986 6660
rect 4968 6660 4986 6678
rect 4968 6678 4986 6696
rect 4968 6696 4986 6714
rect 4968 6714 4986 6732
rect 4968 6732 4986 6750
rect 4968 6750 4986 6768
rect 4968 6768 4986 6786
rect 4968 6786 4986 6804
rect 4968 6804 4986 6822
rect 4968 6822 4986 6840
rect 4968 6840 4986 6858
rect 4968 6858 4986 6876
rect 4968 6876 4986 6894
rect 4968 6894 4986 6912
rect 4968 6912 4986 6930
rect 4968 6930 4986 6948
rect 4968 6948 4986 6966
rect 4968 6966 4986 6984
rect 4968 6984 4986 7002
rect 4968 7002 4986 7020
rect 4968 7020 4986 7038
rect 4968 7038 4986 7056
rect 4968 7056 4986 7074
rect 4968 7074 4986 7092
rect 4968 7092 4986 7110
rect 4968 7110 4986 7128
rect 4968 7128 4986 7146
rect 4968 7146 4986 7164
rect 4968 7164 4986 7182
rect 4968 7182 4986 7200
rect 4968 7200 4986 7218
rect 4968 7218 4986 7236
rect 4968 7236 4986 7254
rect 4968 7254 4986 7272
rect 4968 7272 4986 7290
rect 4968 7290 4986 7308
rect 4968 7308 4986 7326
rect 4968 7326 4986 7344
rect 4968 7344 4986 7362
rect 4968 7362 4986 7380
rect 4968 7380 4986 7398
rect 4968 7398 4986 7416
rect 4968 7416 4986 7434
rect 4968 7434 4986 7452
rect 4968 7452 4986 7470
rect 4968 7470 4986 7488
rect 4968 7488 4986 7506
rect 4968 7506 4986 7524
rect 4968 7524 4986 7542
rect 4968 7542 4986 7560
rect 4968 7560 4986 7578
rect 4968 7578 4986 7596
rect 4968 7596 4986 7614
rect 4968 7614 4986 7632
rect 4968 7632 4986 7650
rect 4968 7650 4986 7668
rect 4968 7668 4986 7686
rect 4968 7686 4986 7704
rect 4968 7704 4986 7722
rect 4968 7722 4986 7740
rect 4968 7740 4986 7758
rect 4968 7758 4986 7776
rect 4968 7776 4986 7794
rect 4986 252 5004 270
rect 4986 270 5004 288
rect 4986 288 5004 306
rect 4986 306 5004 324
rect 4986 324 5004 342
rect 4986 342 5004 360
rect 4986 360 5004 378
rect 4986 378 5004 396
rect 4986 396 5004 414
rect 4986 414 5004 432
rect 4986 432 5004 450
rect 4986 450 5004 468
rect 4986 468 5004 486
rect 4986 486 5004 504
rect 4986 504 5004 522
rect 4986 522 5004 540
rect 4986 540 5004 558
rect 4986 558 5004 576
rect 4986 576 5004 594
rect 4986 594 5004 612
rect 4986 612 5004 630
rect 4986 630 5004 648
rect 4986 648 5004 666
rect 4986 666 5004 684
rect 4986 684 5004 702
rect 4986 702 5004 720
rect 4986 720 5004 738
rect 4986 738 5004 756
rect 4986 864 5004 882
rect 4986 882 5004 900
rect 4986 900 5004 918
rect 4986 918 5004 936
rect 4986 936 5004 954
rect 4986 954 5004 972
rect 4986 972 5004 990
rect 4986 990 5004 1008
rect 4986 1008 5004 1026
rect 4986 1026 5004 1044
rect 4986 1044 5004 1062
rect 4986 1062 5004 1080
rect 4986 1080 5004 1098
rect 4986 1098 5004 1116
rect 4986 1116 5004 1134
rect 4986 1134 5004 1152
rect 4986 1152 5004 1170
rect 4986 1170 5004 1188
rect 4986 1188 5004 1206
rect 4986 1206 5004 1224
rect 4986 1224 5004 1242
rect 4986 1242 5004 1260
rect 4986 1260 5004 1278
rect 4986 1278 5004 1296
rect 4986 1296 5004 1314
rect 4986 1314 5004 1332
rect 4986 1332 5004 1350
rect 4986 1350 5004 1368
rect 4986 1368 5004 1386
rect 4986 1386 5004 1404
rect 4986 1404 5004 1422
rect 4986 1422 5004 1440
rect 4986 1440 5004 1458
rect 4986 1458 5004 1476
rect 4986 1476 5004 1494
rect 4986 1494 5004 1512
rect 4986 1512 5004 1530
rect 4986 1530 5004 1548
rect 4986 1548 5004 1566
rect 4986 1566 5004 1584
rect 4986 1584 5004 1602
rect 4986 1602 5004 1620
rect 4986 1620 5004 1638
rect 4986 1638 5004 1656
rect 4986 1656 5004 1674
rect 4986 1674 5004 1692
rect 4986 1692 5004 1710
rect 4986 1710 5004 1728
rect 4986 1728 5004 1746
rect 4986 1746 5004 1764
rect 4986 1764 5004 1782
rect 4986 1782 5004 1800
rect 4986 1800 5004 1818
rect 4986 1818 5004 1836
rect 4986 1836 5004 1854
rect 4986 1854 5004 1872
rect 4986 1872 5004 1890
rect 4986 1890 5004 1908
rect 4986 1908 5004 1926
rect 4986 1926 5004 1944
rect 4986 1944 5004 1962
rect 4986 1962 5004 1980
rect 4986 1980 5004 1998
rect 4986 1998 5004 2016
rect 4986 2016 5004 2034
rect 4986 2034 5004 2052
rect 4986 2052 5004 2070
rect 4986 2070 5004 2088
rect 4986 2088 5004 2106
rect 4986 2106 5004 2124
rect 4986 2124 5004 2142
rect 4986 2142 5004 2160
rect 4986 2160 5004 2178
rect 4986 2178 5004 2196
rect 4986 2196 5004 2214
rect 4986 2430 5004 2448
rect 4986 2448 5004 2466
rect 4986 2466 5004 2484
rect 4986 2484 5004 2502
rect 4986 2502 5004 2520
rect 4986 2520 5004 2538
rect 4986 2538 5004 2556
rect 4986 2556 5004 2574
rect 4986 2574 5004 2592
rect 4986 2592 5004 2610
rect 4986 2610 5004 2628
rect 4986 2628 5004 2646
rect 4986 2646 5004 2664
rect 4986 2664 5004 2682
rect 4986 2682 5004 2700
rect 4986 2700 5004 2718
rect 4986 2718 5004 2736
rect 4986 2736 5004 2754
rect 4986 2754 5004 2772
rect 4986 2772 5004 2790
rect 4986 2790 5004 2808
rect 4986 2808 5004 2826
rect 4986 2826 5004 2844
rect 4986 2844 5004 2862
rect 4986 2862 5004 2880
rect 4986 2880 5004 2898
rect 4986 2898 5004 2916
rect 4986 2916 5004 2934
rect 4986 2934 5004 2952
rect 4986 2952 5004 2970
rect 4986 2970 5004 2988
rect 4986 2988 5004 3006
rect 4986 3006 5004 3024
rect 4986 3024 5004 3042
rect 4986 3042 5004 3060
rect 4986 3060 5004 3078
rect 4986 3078 5004 3096
rect 4986 3096 5004 3114
rect 4986 3114 5004 3132
rect 4986 3132 5004 3150
rect 4986 3150 5004 3168
rect 4986 3168 5004 3186
rect 4986 3186 5004 3204
rect 4986 3204 5004 3222
rect 4986 3222 5004 3240
rect 4986 3240 5004 3258
rect 4986 3258 5004 3276
rect 4986 3276 5004 3294
rect 4986 3294 5004 3312
rect 4986 3312 5004 3330
rect 4986 3330 5004 3348
rect 4986 3348 5004 3366
rect 4986 3366 5004 3384
rect 4986 3384 5004 3402
rect 4986 3402 5004 3420
rect 4986 3420 5004 3438
rect 4986 3438 5004 3456
rect 4986 3456 5004 3474
rect 4986 3474 5004 3492
rect 4986 3492 5004 3510
rect 4986 3510 5004 3528
rect 4986 3528 5004 3546
rect 4986 3546 5004 3564
rect 4986 3564 5004 3582
rect 4986 3582 5004 3600
rect 4986 3600 5004 3618
rect 4986 3618 5004 3636
rect 4986 3636 5004 3654
rect 4986 3654 5004 3672
rect 4986 3672 5004 3690
rect 4986 3690 5004 3708
rect 4986 3708 5004 3726
rect 4986 3726 5004 3744
rect 4986 3744 5004 3762
rect 4986 3762 5004 3780
rect 4986 3780 5004 3798
rect 4986 3798 5004 3816
rect 4986 3816 5004 3834
rect 4986 3834 5004 3852
rect 4986 3852 5004 3870
rect 4986 3870 5004 3888
rect 4986 3888 5004 3906
rect 4986 3906 5004 3924
rect 4986 3924 5004 3942
rect 4986 3942 5004 3960
rect 4986 3960 5004 3978
rect 4986 3978 5004 3996
rect 4986 3996 5004 4014
rect 4986 4014 5004 4032
rect 4986 4032 5004 4050
rect 4986 4050 5004 4068
rect 4986 4068 5004 4086
rect 4986 4086 5004 4104
rect 4986 4104 5004 4122
rect 4986 4122 5004 4140
rect 4986 4140 5004 4158
rect 4986 4158 5004 4176
rect 4986 4176 5004 4194
rect 4986 4194 5004 4212
rect 4986 4212 5004 4230
rect 4986 4230 5004 4248
rect 4986 4248 5004 4266
rect 4986 4266 5004 4284
rect 4986 4284 5004 4302
rect 4986 4302 5004 4320
rect 4986 4320 5004 4338
rect 4986 4338 5004 4356
rect 4986 4356 5004 4374
rect 4986 4572 5004 4590
rect 4986 4590 5004 4608
rect 4986 4608 5004 4626
rect 4986 4626 5004 4644
rect 4986 4644 5004 4662
rect 4986 4662 5004 4680
rect 4986 4680 5004 4698
rect 4986 4698 5004 4716
rect 4986 4716 5004 4734
rect 4986 4734 5004 4752
rect 4986 4752 5004 4770
rect 4986 4770 5004 4788
rect 4986 4788 5004 4806
rect 4986 4806 5004 4824
rect 4986 4824 5004 4842
rect 4986 4842 5004 4860
rect 4986 4860 5004 4878
rect 4986 4878 5004 4896
rect 4986 4896 5004 4914
rect 4986 4914 5004 4932
rect 4986 4932 5004 4950
rect 4986 4950 5004 4968
rect 4986 4968 5004 4986
rect 4986 4986 5004 5004
rect 4986 5004 5004 5022
rect 4986 5022 5004 5040
rect 4986 5040 5004 5058
rect 4986 5058 5004 5076
rect 4986 5076 5004 5094
rect 4986 5094 5004 5112
rect 4986 5112 5004 5130
rect 4986 5130 5004 5148
rect 4986 5148 5004 5166
rect 4986 5166 5004 5184
rect 4986 5184 5004 5202
rect 4986 5202 5004 5220
rect 4986 5220 5004 5238
rect 4986 5238 5004 5256
rect 4986 5256 5004 5274
rect 4986 5274 5004 5292
rect 4986 5292 5004 5310
rect 4986 5310 5004 5328
rect 4986 5328 5004 5346
rect 4986 5346 5004 5364
rect 4986 5364 5004 5382
rect 4986 5382 5004 5400
rect 4986 5400 5004 5418
rect 4986 5418 5004 5436
rect 4986 5436 5004 5454
rect 4986 5454 5004 5472
rect 4986 5472 5004 5490
rect 4986 5490 5004 5508
rect 4986 5508 5004 5526
rect 4986 5526 5004 5544
rect 4986 5544 5004 5562
rect 4986 5562 5004 5580
rect 4986 5580 5004 5598
rect 4986 5598 5004 5616
rect 4986 5616 5004 5634
rect 4986 5634 5004 5652
rect 4986 5652 5004 5670
rect 4986 5670 5004 5688
rect 4986 5688 5004 5706
rect 4986 5706 5004 5724
rect 4986 5724 5004 5742
rect 4986 5742 5004 5760
rect 4986 5760 5004 5778
rect 4986 5778 5004 5796
rect 4986 5796 5004 5814
rect 4986 5814 5004 5832
rect 4986 5832 5004 5850
rect 4986 5850 5004 5868
rect 4986 5868 5004 5886
rect 4986 5886 5004 5904
rect 4986 5904 5004 5922
rect 4986 5922 5004 5940
rect 4986 5940 5004 5958
rect 4986 5958 5004 5976
rect 4986 5976 5004 5994
rect 4986 5994 5004 6012
rect 4986 6012 5004 6030
rect 4986 6030 5004 6048
rect 4986 6048 5004 6066
rect 4986 6066 5004 6084
rect 4986 6084 5004 6102
rect 4986 6102 5004 6120
rect 4986 6120 5004 6138
rect 4986 6138 5004 6156
rect 4986 6156 5004 6174
rect 4986 6174 5004 6192
rect 4986 6192 5004 6210
rect 4986 6210 5004 6228
rect 4986 6228 5004 6246
rect 4986 6246 5004 6264
rect 4986 6264 5004 6282
rect 4986 6282 5004 6300
rect 4986 6300 5004 6318
rect 4986 6318 5004 6336
rect 4986 6336 5004 6354
rect 4986 6354 5004 6372
rect 4986 6372 5004 6390
rect 4986 6390 5004 6408
rect 4986 6408 5004 6426
rect 4986 6426 5004 6444
rect 4986 6444 5004 6462
rect 4986 6462 5004 6480
rect 4986 6480 5004 6498
rect 4986 6498 5004 6516
rect 4986 6516 5004 6534
rect 4986 6534 5004 6552
rect 4986 6552 5004 6570
rect 4986 6570 5004 6588
rect 4986 6588 5004 6606
rect 4986 6606 5004 6624
rect 4986 6624 5004 6642
rect 4986 6642 5004 6660
rect 4986 6660 5004 6678
rect 4986 6678 5004 6696
rect 4986 6696 5004 6714
rect 4986 6714 5004 6732
rect 4986 6732 5004 6750
rect 4986 6750 5004 6768
rect 4986 6768 5004 6786
rect 4986 6786 5004 6804
rect 4986 6804 5004 6822
rect 4986 6822 5004 6840
rect 4986 6840 5004 6858
rect 4986 6858 5004 6876
rect 4986 6876 5004 6894
rect 4986 6894 5004 6912
rect 4986 6912 5004 6930
rect 4986 6930 5004 6948
rect 4986 6948 5004 6966
rect 4986 6966 5004 6984
rect 4986 6984 5004 7002
rect 4986 7002 5004 7020
rect 4986 7020 5004 7038
rect 4986 7038 5004 7056
rect 4986 7056 5004 7074
rect 4986 7074 5004 7092
rect 4986 7092 5004 7110
rect 4986 7110 5004 7128
rect 4986 7128 5004 7146
rect 4986 7146 5004 7164
rect 4986 7164 5004 7182
rect 4986 7182 5004 7200
rect 4986 7200 5004 7218
rect 4986 7218 5004 7236
rect 4986 7236 5004 7254
rect 4986 7254 5004 7272
rect 4986 7272 5004 7290
rect 4986 7290 5004 7308
rect 4986 7308 5004 7326
rect 4986 7326 5004 7344
rect 4986 7344 5004 7362
rect 4986 7362 5004 7380
rect 4986 7380 5004 7398
rect 4986 7398 5004 7416
rect 4986 7416 5004 7434
rect 4986 7434 5004 7452
rect 4986 7452 5004 7470
rect 4986 7470 5004 7488
rect 4986 7488 5004 7506
rect 4986 7506 5004 7524
rect 4986 7524 5004 7542
rect 4986 7542 5004 7560
rect 4986 7560 5004 7578
rect 4986 7578 5004 7596
rect 4986 7596 5004 7614
rect 4986 7614 5004 7632
rect 4986 7632 5004 7650
rect 4986 7650 5004 7668
rect 4986 7668 5004 7686
rect 4986 7686 5004 7704
rect 4986 7704 5004 7722
rect 4986 7722 5004 7740
rect 4986 7740 5004 7758
rect 4986 7758 5004 7776
rect 4986 7776 5004 7794
rect 4986 7794 5004 7812
rect 4986 7812 5004 7830
rect 5004 270 5022 288
rect 5004 288 5022 306
rect 5004 306 5022 324
rect 5004 324 5022 342
rect 5004 342 5022 360
rect 5004 360 5022 378
rect 5004 378 5022 396
rect 5004 396 5022 414
rect 5004 414 5022 432
rect 5004 432 5022 450
rect 5004 450 5022 468
rect 5004 468 5022 486
rect 5004 486 5022 504
rect 5004 504 5022 522
rect 5004 522 5022 540
rect 5004 540 5022 558
rect 5004 558 5022 576
rect 5004 576 5022 594
rect 5004 594 5022 612
rect 5004 612 5022 630
rect 5004 630 5022 648
rect 5004 648 5022 666
rect 5004 666 5022 684
rect 5004 684 5022 702
rect 5004 702 5022 720
rect 5004 720 5022 738
rect 5004 738 5022 756
rect 5004 864 5022 882
rect 5004 882 5022 900
rect 5004 900 5022 918
rect 5004 918 5022 936
rect 5004 936 5022 954
rect 5004 954 5022 972
rect 5004 972 5022 990
rect 5004 990 5022 1008
rect 5004 1008 5022 1026
rect 5004 1026 5022 1044
rect 5004 1044 5022 1062
rect 5004 1062 5022 1080
rect 5004 1080 5022 1098
rect 5004 1098 5022 1116
rect 5004 1116 5022 1134
rect 5004 1134 5022 1152
rect 5004 1152 5022 1170
rect 5004 1170 5022 1188
rect 5004 1188 5022 1206
rect 5004 1206 5022 1224
rect 5004 1224 5022 1242
rect 5004 1242 5022 1260
rect 5004 1260 5022 1278
rect 5004 1278 5022 1296
rect 5004 1296 5022 1314
rect 5004 1314 5022 1332
rect 5004 1332 5022 1350
rect 5004 1350 5022 1368
rect 5004 1368 5022 1386
rect 5004 1386 5022 1404
rect 5004 1404 5022 1422
rect 5004 1422 5022 1440
rect 5004 1440 5022 1458
rect 5004 1458 5022 1476
rect 5004 1476 5022 1494
rect 5004 1494 5022 1512
rect 5004 1512 5022 1530
rect 5004 1530 5022 1548
rect 5004 1548 5022 1566
rect 5004 1566 5022 1584
rect 5004 1584 5022 1602
rect 5004 1602 5022 1620
rect 5004 1620 5022 1638
rect 5004 1638 5022 1656
rect 5004 1656 5022 1674
rect 5004 1674 5022 1692
rect 5004 1692 5022 1710
rect 5004 1710 5022 1728
rect 5004 1728 5022 1746
rect 5004 1746 5022 1764
rect 5004 1764 5022 1782
rect 5004 1782 5022 1800
rect 5004 1800 5022 1818
rect 5004 1818 5022 1836
rect 5004 1836 5022 1854
rect 5004 1854 5022 1872
rect 5004 1872 5022 1890
rect 5004 1890 5022 1908
rect 5004 1908 5022 1926
rect 5004 1926 5022 1944
rect 5004 1944 5022 1962
rect 5004 1962 5022 1980
rect 5004 1980 5022 1998
rect 5004 1998 5022 2016
rect 5004 2016 5022 2034
rect 5004 2034 5022 2052
rect 5004 2052 5022 2070
rect 5004 2070 5022 2088
rect 5004 2088 5022 2106
rect 5004 2106 5022 2124
rect 5004 2124 5022 2142
rect 5004 2142 5022 2160
rect 5004 2160 5022 2178
rect 5004 2178 5022 2196
rect 5004 2196 5022 2214
rect 5004 2214 5022 2232
rect 5004 2448 5022 2466
rect 5004 2466 5022 2484
rect 5004 2484 5022 2502
rect 5004 2502 5022 2520
rect 5004 2520 5022 2538
rect 5004 2538 5022 2556
rect 5004 2556 5022 2574
rect 5004 2574 5022 2592
rect 5004 2592 5022 2610
rect 5004 2610 5022 2628
rect 5004 2628 5022 2646
rect 5004 2646 5022 2664
rect 5004 2664 5022 2682
rect 5004 2682 5022 2700
rect 5004 2700 5022 2718
rect 5004 2718 5022 2736
rect 5004 2736 5022 2754
rect 5004 2754 5022 2772
rect 5004 2772 5022 2790
rect 5004 2790 5022 2808
rect 5004 2808 5022 2826
rect 5004 2826 5022 2844
rect 5004 2844 5022 2862
rect 5004 2862 5022 2880
rect 5004 2880 5022 2898
rect 5004 2898 5022 2916
rect 5004 2916 5022 2934
rect 5004 2934 5022 2952
rect 5004 2952 5022 2970
rect 5004 2970 5022 2988
rect 5004 2988 5022 3006
rect 5004 3006 5022 3024
rect 5004 3024 5022 3042
rect 5004 3042 5022 3060
rect 5004 3060 5022 3078
rect 5004 3078 5022 3096
rect 5004 3096 5022 3114
rect 5004 3114 5022 3132
rect 5004 3132 5022 3150
rect 5004 3150 5022 3168
rect 5004 3168 5022 3186
rect 5004 3186 5022 3204
rect 5004 3204 5022 3222
rect 5004 3222 5022 3240
rect 5004 3240 5022 3258
rect 5004 3258 5022 3276
rect 5004 3276 5022 3294
rect 5004 3294 5022 3312
rect 5004 3312 5022 3330
rect 5004 3330 5022 3348
rect 5004 3348 5022 3366
rect 5004 3366 5022 3384
rect 5004 3384 5022 3402
rect 5004 3402 5022 3420
rect 5004 3420 5022 3438
rect 5004 3438 5022 3456
rect 5004 3456 5022 3474
rect 5004 3474 5022 3492
rect 5004 3492 5022 3510
rect 5004 3510 5022 3528
rect 5004 3528 5022 3546
rect 5004 3546 5022 3564
rect 5004 3564 5022 3582
rect 5004 3582 5022 3600
rect 5004 3600 5022 3618
rect 5004 3618 5022 3636
rect 5004 3636 5022 3654
rect 5004 3654 5022 3672
rect 5004 3672 5022 3690
rect 5004 3690 5022 3708
rect 5004 3708 5022 3726
rect 5004 3726 5022 3744
rect 5004 3744 5022 3762
rect 5004 3762 5022 3780
rect 5004 3780 5022 3798
rect 5004 3798 5022 3816
rect 5004 3816 5022 3834
rect 5004 3834 5022 3852
rect 5004 3852 5022 3870
rect 5004 3870 5022 3888
rect 5004 3888 5022 3906
rect 5004 3906 5022 3924
rect 5004 3924 5022 3942
rect 5004 3942 5022 3960
rect 5004 3960 5022 3978
rect 5004 3978 5022 3996
rect 5004 3996 5022 4014
rect 5004 4014 5022 4032
rect 5004 4032 5022 4050
rect 5004 4050 5022 4068
rect 5004 4068 5022 4086
rect 5004 4086 5022 4104
rect 5004 4104 5022 4122
rect 5004 4122 5022 4140
rect 5004 4140 5022 4158
rect 5004 4158 5022 4176
rect 5004 4176 5022 4194
rect 5004 4194 5022 4212
rect 5004 4212 5022 4230
rect 5004 4230 5022 4248
rect 5004 4248 5022 4266
rect 5004 4266 5022 4284
rect 5004 4284 5022 4302
rect 5004 4302 5022 4320
rect 5004 4320 5022 4338
rect 5004 4338 5022 4356
rect 5004 4356 5022 4374
rect 5004 4374 5022 4392
rect 5004 4590 5022 4608
rect 5004 4608 5022 4626
rect 5004 4626 5022 4644
rect 5004 4644 5022 4662
rect 5004 4662 5022 4680
rect 5004 4680 5022 4698
rect 5004 4698 5022 4716
rect 5004 4716 5022 4734
rect 5004 4734 5022 4752
rect 5004 4752 5022 4770
rect 5004 4770 5022 4788
rect 5004 4788 5022 4806
rect 5004 4806 5022 4824
rect 5004 4824 5022 4842
rect 5004 4842 5022 4860
rect 5004 4860 5022 4878
rect 5004 4878 5022 4896
rect 5004 4896 5022 4914
rect 5004 4914 5022 4932
rect 5004 4932 5022 4950
rect 5004 4950 5022 4968
rect 5004 4968 5022 4986
rect 5004 4986 5022 5004
rect 5004 5004 5022 5022
rect 5004 5022 5022 5040
rect 5004 5040 5022 5058
rect 5004 5058 5022 5076
rect 5004 5076 5022 5094
rect 5004 5094 5022 5112
rect 5004 5112 5022 5130
rect 5004 5130 5022 5148
rect 5004 5148 5022 5166
rect 5004 5166 5022 5184
rect 5004 5184 5022 5202
rect 5004 5202 5022 5220
rect 5004 5220 5022 5238
rect 5004 5238 5022 5256
rect 5004 5256 5022 5274
rect 5004 5274 5022 5292
rect 5004 5292 5022 5310
rect 5004 5310 5022 5328
rect 5004 5328 5022 5346
rect 5004 5346 5022 5364
rect 5004 5364 5022 5382
rect 5004 5382 5022 5400
rect 5004 5400 5022 5418
rect 5004 5418 5022 5436
rect 5004 5436 5022 5454
rect 5004 5454 5022 5472
rect 5004 5472 5022 5490
rect 5004 5490 5022 5508
rect 5004 5508 5022 5526
rect 5004 5526 5022 5544
rect 5004 5544 5022 5562
rect 5004 5562 5022 5580
rect 5004 5580 5022 5598
rect 5004 5598 5022 5616
rect 5004 5616 5022 5634
rect 5004 5634 5022 5652
rect 5004 5652 5022 5670
rect 5004 5670 5022 5688
rect 5004 5688 5022 5706
rect 5004 5706 5022 5724
rect 5004 5724 5022 5742
rect 5004 5742 5022 5760
rect 5004 5760 5022 5778
rect 5004 5778 5022 5796
rect 5004 5796 5022 5814
rect 5004 5814 5022 5832
rect 5004 5832 5022 5850
rect 5004 5850 5022 5868
rect 5004 5868 5022 5886
rect 5004 5886 5022 5904
rect 5004 5904 5022 5922
rect 5004 5922 5022 5940
rect 5004 5940 5022 5958
rect 5004 5958 5022 5976
rect 5004 5976 5022 5994
rect 5004 5994 5022 6012
rect 5004 6012 5022 6030
rect 5004 6030 5022 6048
rect 5004 6048 5022 6066
rect 5004 6066 5022 6084
rect 5004 6084 5022 6102
rect 5004 6102 5022 6120
rect 5004 6120 5022 6138
rect 5004 6138 5022 6156
rect 5004 6156 5022 6174
rect 5004 6174 5022 6192
rect 5004 6192 5022 6210
rect 5004 6210 5022 6228
rect 5004 6228 5022 6246
rect 5004 6246 5022 6264
rect 5004 6264 5022 6282
rect 5004 6282 5022 6300
rect 5004 6300 5022 6318
rect 5004 6318 5022 6336
rect 5004 6336 5022 6354
rect 5004 6354 5022 6372
rect 5004 6372 5022 6390
rect 5004 6390 5022 6408
rect 5004 6408 5022 6426
rect 5004 6426 5022 6444
rect 5004 6444 5022 6462
rect 5004 6462 5022 6480
rect 5004 6480 5022 6498
rect 5004 6498 5022 6516
rect 5004 6516 5022 6534
rect 5004 6534 5022 6552
rect 5004 6552 5022 6570
rect 5004 6570 5022 6588
rect 5004 6588 5022 6606
rect 5004 6606 5022 6624
rect 5004 6624 5022 6642
rect 5004 6642 5022 6660
rect 5004 6660 5022 6678
rect 5004 6678 5022 6696
rect 5004 6696 5022 6714
rect 5004 6714 5022 6732
rect 5004 6732 5022 6750
rect 5004 6750 5022 6768
rect 5004 6768 5022 6786
rect 5004 6786 5022 6804
rect 5004 6804 5022 6822
rect 5004 6822 5022 6840
rect 5004 6840 5022 6858
rect 5004 6858 5022 6876
rect 5004 6876 5022 6894
rect 5004 6894 5022 6912
rect 5004 6912 5022 6930
rect 5004 6930 5022 6948
rect 5004 6948 5022 6966
rect 5004 6966 5022 6984
rect 5004 6984 5022 7002
rect 5004 7002 5022 7020
rect 5004 7020 5022 7038
rect 5004 7038 5022 7056
rect 5004 7056 5022 7074
rect 5004 7074 5022 7092
rect 5004 7092 5022 7110
rect 5004 7110 5022 7128
rect 5004 7128 5022 7146
rect 5004 7146 5022 7164
rect 5004 7164 5022 7182
rect 5004 7182 5022 7200
rect 5004 7200 5022 7218
rect 5004 7218 5022 7236
rect 5004 7236 5022 7254
rect 5004 7254 5022 7272
rect 5004 7272 5022 7290
rect 5004 7290 5022 7308
rect 5004 7308 5022 7326
rect 5004 7326 5022 7344
rect 5004 7344 5022 7362
rect 5004 7362 5022 7380
rect 5004 7380 5022 7398
rect 5004 7398 5022 7416
rect 5004 7416 5022 7434
rect 5004 7434 5022 7452
rect 5004 7452 5022 7470
rect 5004 7470 5022 7488
rect 5004 7488 5022 7506
rect 5004 7506 5022 7524
rect 5004 7524 5022 7542
rect 5004 7542 5022 7560
rect 5004 7560 5022 7578
rect 5004 7578 5022 7596
rect 5004 7596 5022 7614
rect 5004 7614 5022 7632
rect 5004 7632 5022 7650
rect 5004 7650 5022 7668
rect 5004 7668 5022 7686
rect 5004 7686 5022 7704
rect 5004 7704 5022 7722
rect 5004 7722 5022 7740
rect 5004 7740 5022 7758
rect 5004 7758 5022 7776
rect 5004 7776 5022 7794
rect 5004 7794 5022 7812
rect 5004 7812 5022 7830
rect 5004 7830 5022 7848
rect 5022 270 5040 288
rect 5022 288 5040 306
rect 5022 306 5040 324
rect 5022 324 5040 342
rect 5022 342 5040 360
rect 5022 360 5040 378
rect 5022 378 5040 396
rect 5022 396 5040 414
rect 5022 414 5040 432
rect 5022 432 5040 450
rect 5022 450 5040 468
rect 5022 468 5040 486
rect 5022 486 5040 504
rect 5022 504 5040 522
rect 5022 522 5040 540
rect 5022 540 5040 558
rect 5022 558 5040 576
rect 5022 576 5040 594
rect 5022 594 5040 612
rect 5022 612 5040 630
rect 5022 630 5040 648
rect 5022 648 5040 666
rect 5022 666 5040 684
rect 5022 684 5040 702
rect 5022 702 5040 720
rect 5022 720 5040 738
rect 5022 738 5040 756
rect 5022 864 5040 882
rect 5022 882 5040 900
rect 5022 900 5040 918
rect 5022 918 5040 936
rect 5022 936 5040 954
rect 5022 954 5040 972
rect 5022 972 5040 990
rect 5022 990 5040 1008
rect 5022 1008 5040 1026
rect 5022 1026 5040 1044
rect 5022 1044 5040 1062
rect 5022 1062 5040 1080
rect 5022 1080 5040 1098
rect 5022 1098 5040 1116
rect 5022 1116 5040 1134
rect 5022 1134 5040 1152
rect 5022 1152 5040 1170
rect 5022 1170 5040 1188
rect 5022 1188 5040 1206
rect 5022 1206 5040 1224
rect 5022 1224 5040 1242
rect 5022 1242 5040 1260
rect 5022 1260 5040 1278
rect 5022 1278 5040 1296
rect 5022 1296 5040 1314
rect 5022 1314 5040 1332
rect 5022 1332 5040 1350
rect 5022 1350 5040 1368
rect 5022 1368 5040 1386
rect 5022 1386 5040 1404
rect 5022 1404 5040 1422
rect 5022 1422 5040 1440
rect 5022 1440 5040 1458
rect 5022 1458 5040 1476
rect 5022 1476 5040 1494
rect 5022 1494 5040 1512
rect 5022 1512 5040 1530
rect 5022 1530 5040 1548
rect 5022 1548 5040 1566
rect 5022 1566 5040 1584
rect 5022 1584 5040 1602
rect 5022 1602 5040 1620
rect 5022 1620 5040 1638
rect 5022 1638 5040 1656
rect 5022 1656 5040 1674
rect 5022 1674 5040 1692
rect 5022 1692 5040 1710
rect 5022 1710 5040 1728
rect 5022 1728 5040 1746
rect 5022 1746 5040 1764
rect 5022 1764 5040 1782
rect 5022 1782 5040 1800
rect 5022 1800 5040 1818
rect 5022 1818 5040 1836
rect 5022 1836 5040 1854
rect 5022 1854 5040 1872
rect 5022 1872 5040 1890
rect 5022 1890 5040 1908
rect 5022 1908 5040 1926
rect 5022 1926 5040 1944
rect 5022 1944 5040 1962
rect 5022 1962 5040 1980
rect 5022 1980 5040 1998
rect 5022 1998 5040 2016
rect 5022 2016 5040 2034
rect 5022 2034 5040 2052
rect 5022 2052 5040 2070
rect 5022 2070 5040 2088
rect 5022 2088 5040 2106
rect 5022 2106 5040 2124
rect 5022 2124 5040 2142
rect 5022 2142 5040 2160
rect 5022 2160 5040 2178
rect 5022 2178 5040 2196
rect 5022 2196 5040 2214
rect 5022 2214 5040 2232
rect 5022 2232 5040 2250
rect 5022 2466 5040 2484
rect 5022 2484 5040 2502
rect 5022 2502 5040 2520
rect 5022 2520 5040 2538
rect 5022 2538 5040 2556
rect 5022 2556 5040 2574
rect 5022 2574 5040 2592
rect 5022 2592 5040 2610
rect 5022 2610 5040 2628
rect 5022 2628 5040 2646
rect 5022 2646 5040 2664
rect 5022 2664 5040 2682
rect 5022 2682 5040 2700
rect 5022 2700 5040 2718
rect 5022 2718 5040 2736
rect 5022 2736 5040 2754
rect 5022 2754 5040 2772
rect 5022 2772 5040 2790
rect 5022 2790 5040 2808
rect 5022 2808 5040 2826
rect 5022 2826 5040 2844
rect 5022 2844 5040 2862
rect 5022 2862 5040 2880
rect 5022 2880 5040 2898
rect 5022 2898 5040 2916
rect 5022 2916 5040 2934
rect 5022 2934 5040 2952
rect 5022 2952 5040 2970
rect 5022 2970 5040 2988
rect 5022 2988 5040 3006
rect 5022 3006 5040 3024
rect 5022 3024 5040 3042
rect 5022 3042 5040 3060
rect 5022 3060 5040 3078
rect 5022 3078 5040 3096
rect 5022 3096 5040 3114
rect 5022 3114 5040 3132
rect 5022 3132 5040 3150
rect 5022 3150 5040 3168
rect 5022 3168 5040 3186
rect 5022 3186 5040 3204
rect 5022 3204 5040 3222
rect 5022 3222 5040 3240
rect 5022 3240 5040 3258
rect 5022 3258 5040 3276
rect 5022 3276 5040 3294
rect 5022 3294 5040 3312
rect 5022 3312 5040 3330
rect 5022 3330 5040 3348
rect 5022 3348 5040 3366
rect 5022 3366 5040 3384
rect 5022 3384 5040 3402
rect 5022 3402 5040 3420
rect 5022 3420 5040 3438
rect 5022 3438 5040 3456
rect 5022 3456 5040 3474
rect 5022 3474 5040 3492
rect 5022 3492 5040 3510
rect 5022 3510 5040 3528
rect 5022 3528 5040 3546
rect 5022 3546 5040 3564
rect 5022 3564 5040 3582
rect 5022 3582 5040 3600
rect 5022 3600 5040 3618
rect 5022 3618 5040 3636
rect 5022 3636 5040 3654
rect 5022 3654 5040 3672
rect 5022 3672 5040 3690
rect 5022 3690 5040 3708
rect 5022 3708 5040 3726
rect 5022 3726 5040 3744
rect 5022 3744 5040 3762
rect 5022 3762 5040 3780
rect 5022 3780 5040 3798
rect 5022 3798 5040 3816
rect 5022 3816 5040 3834
rect 5022 3834 5040 3852
rect 5022 3852 5040 3870
rect 5022 3870 5040 3888
rect 5022 3888 5040 3906
rect 5022 3906 5040 3924
rect 5022 3924 5040 3942
rect 5022 3942 5040 3960
rect 5022 3960 5040 3978
rect 5022 3978 5040 3996
rect 5022 3996 5040 4014
rect 5022 4014 5040 4032
rect 5022 4032 5040 4050
rect 5022 4050 5040 4068
rect 5022 4068 5040 4086
rect 5022 4086 5040 4104
rect 5022 4104 5040 4122
rect 5022 4122 5040 4140
rect 5022 4140 5040 4158
rect 5022 4158 5040 4176
rect 5022 4176 5040 4194
rect 5022 4194 5040 4212
rect 5022 4212 5040 4230
rect 5022 4230 5040 4248
rect 5022 4248 5040 4266
rect 5022 4266 5040 4284
rect 5022 4284 5040 4302
rect 5022 4302 5040 4320
rect 5022 4320 5040 4338
rect 5022 4338 5040 4356
rect 5022 4356 5040 4374
rect 5022 4374 5040 4392
rect 5022 4392 5040 4410
rect 5022 4626 5040 4644
rect 5022 4644 5040 4662
rect 5022 4662 5040 4680
rect 5022 4680 5040 4698
rect 5022 4698 5040 4716
rect 5022 4716 5040 4734
rect 5022 4734 5040 4752
rect 5022 4752 5040 4770
rect 5022 4770 5040 4788
rect 5022 4788 5040 4806
rect 5022 4806 5040 4824
rect 5022 4824 5040 4842
rect 5022 4842 5040 4860
rect 5022 4860 5040 4878
rect 5022 4878 5040 4896
rect 5022 4896 5040 4914
rect 5022 4914 5040 4932
rect 5022 4932 5040 4950
rect 5022 4950 5040 4968
rect 5022 4968 5040 4986
rect 5022 4986 5040 5004
rect 5022 5004 5040 5022
rect 5022 5022 5040 5040
rect 5022 5040 5040 5058
rect 5022 5058 5040 5076
rect 5022 5076 5040 5094
rect 5022 5094 5040 5112
rect 5022 5112 5040 5130
rect 5022 5130 5040 5148
rect 5022 5148 5040 5166
rect 5022 5166 5040 5184
rect 5022 5184 5040 5202
rect 5022 5202 5040 5220
rect 5022 5220 5040 5238
rect 5022 5238 5040 5256
rect 5022 5256 5040 5274
rect 5022 5274 5040 5292
rect 5022 5292 5040 5310
rect 5022 5310 5040 5328
rect 5022 5328 5040 5346
rect 5022 5346 5040 5364
rect 5022 5364 5040 5382
rect 5022 5382 5040 5400
rect 5022 5400 5040 5418
rect 5022 5418 5040 5436
rect 5022 5436 5040 5454
rect 5022 5454 5040 5472
rect 5022 5472 5040 5490
rect 5022 5490 5040 5508
rect 5022 5508 5040 5526
rect 5022 5526 5040 5544
rect 5022 5544 5040 5562
rect 5022 5562 5040 5580
rect 5022 5580 5040 5598
rect 5022 5598 5040 5616
rect 5022 5616 5040 5634
rect 5022 5634 5040 5652
rect 5022 5652 5040 5670
rect 5022 5670 5040 5688
rect 5022 5688 5040 5706
rect 5022 5706 5040 5724
rect 5022 5724 5040 5742
rect 5022 5742 5040 5760
rect 5022 5760 5040 5778
rect 5022 5778 5040 5796
rect 5022 5796 5040 5814
rect 5022 5814 5040 5832
rect 5022 5832 5040 5850
rect 5022 5850 5040 5868
rect 5022 5868 5040 5886
rect 5022 5886 5040 5904
rect 5022 5904 5040 5922
rect 5022 5922 5040 5940
rect 5022 5940 5040 5958
rect 5022 5958 5040 5976
rect 5022 5976 5040 5994
rect 5022 5994 5040 6012
rect 5022 6012 5040 6030
rect 5022 6030 5040 6048
rect 5022 6048 5040 6066
rect 5022 6066 5040 6084
rect 5022 6084 5040 6102
rect 5022 6102 5040 6120
rect 5022 6120 5040 6138
rect 5022 6138 5040 6156
rect 5022 6156 5040 6174
rect 5022 6174 5040 6192
rect 5022 6192 5040 6210
rect 5022 6210 5040 6228
rect 5022 6228 5040 6246
rect 5022 6246 5040 6264
rect 5022 6264 5040 6282
rect 5022 6282 5040 6300
rect 5022 6300 5040 6318
rect 5022 6318 5040 6336
rect 5022 6336 5040 6354
rect 5022 6354 5040 6372
rect 5022 6372 5040 6390
rect 5022 6390 5040 6408
rect 5022 6408 5040 6426
rect 5022 6426 5040 6444
rect 5022 6444 5040 6462
rect 5022 6462 5040 6480
rect 5022 6480 5040 6498
rect 5022 6498 5040 6516
rect 5022 6516 5040 6534
rect 5022 6534 5040 6552
rect 5022 6552 5040 6570
rect 5022 6570 5040 6588
rect 5022 6588 5040 6606
rect 5022 6606 5040 6624
rect 5022 6624 5040 6642
rect 5022 6642 5040 6660
rect 5022 6660 5040 6678
rect 5022 6678 5040 6696
rect 5022 6696 5040 6714
rect 5022 6714 5040 6732
rect 5022 6732 5040 6750
rect 5022 6750 5040 6768
rect 5022 6768 5040 6786
rect 5022 6786 5040 6804
rect 5022 6804 5040 6822
rect 5022 6822 5040 6840
rect 5022 6840 5040 6858
rect 5022 6858 5040 6876
rect 5022 6876 5040 6894
rect 5022 6894 5040 6912
rect 5022 6912 5040 6930
rect 5022 6930 5040 6948
rect 5022 6948 5040 6966
rect 5022 6966 5040 6984
rect 5022 6984 5040 7002
rect 5022 7002 5040 7020
rect 5022 7020 5040 7038
rect 5022 7038 5040 7056
rect 5022 7056 5040 7074
rect 5022 7074 5040 7092
rect 5022 7092 5040 7110
rect 5022 7110 5040 7128
rect 5022 7128 5040 7146
rect 5022 7146 5040 7164
rect 5022 7164 5040 7182
rect 5022 7182 5040 7200
rect 5022 7200 5040 7218
rect 5022 7218 5040 7236
rect 5022 7236 5040 7254
rect 5022 7254 5040 7272
rect 5022 7272 5040 7290
rect 5022 7290 5040 7308
rect 5022 7308 5040 7326
rect 5022 7326 5040 7344
rect 5022 7344 5040 7362
rect 5022 7362 5040 7380
rect 5022 7380 5040 7398
rect 5022 7398 5040 7416
rect 5022 7416 5040 7434
rect 5022 7434 5040 7452
rect 5022 7452 5040 7470
rect 5022 7470 5040 7488
rect 5022 7488 5040 7506
rect 5022 7506 5040 7524
rect 5022 7524 5040 7542
rect 5022 7542 5040 7560
rect 5022 7560 5040 7578
rect 5022 7578 5040 7596
rect 5022 7596 5040 7614
rect 5022 7614 5040 7632
rect 5022 7632 5040 7650
rect 5022 7650 5040 7668
rect 5022 7668 5040 7686
rect 5022 7686 5040 7704
rect 5022 7704 5040 7722
rect 5022 7722 5040 7740
rect 5022 7740 5040 7758
rect 5022 7758 5040 7776
rect 5022 7776 5040 7794
rect 5022 7794 5040 7812
rect 5022 7812 5040 7830
rect 5022 7830 5040 7848
rect 5022 7848 5040 7866
rect 5022 7866 5040 7884
rect 5040 288 5058 306
rect 5040 306 5058 324
rect 5040 324 5058 342
rect 5040 342 5058 360
rect 5040 360 5058 378
rect 5040 378 5058 396
rect 5040 396 5058 414
rect 5040 414 5058 432
rect 5040 432 5058 450
rect 5040 450 5058 468
rect 5040 468 5058 486
rect 5040 486 5058 504
rect 5040 504 5058 522
rect 5040 522 5058 540
rect 5040 540 5058 558
rect 5040 558 5058 576
rect 5040 576 5058 594
rect 5040 594 5058 612
rect 5040 612 5058 630
rect 5040 630 5058 648
rect 5040 648 5058 666
rect 5040 666 5058 684
rect 5040 684 5058 702
rect 5040 702 5058 720
rect 5040 720 5058 738
rect 5040 738 5058 756
rect 5040 882 5058 900
rect 5040 900 5058 918
rect 5040 918 5058 936
rect 5040 936 5058 954
rect 5040 954 5058 972
rect 5040 972 5058 990
rect 5040 990 5058 1008
rect 5040 1008 5058 1026
rect 5040 1026 5058 1044
rect 5040 1044 5058 1062
rect 5040 1062 5058 1080
rect 5040 1080 5058 1098
rect 5040 1098 5058 1116
rect 5040 1116 5058 1134
rect 5040 1134 5058 1152
rect 5040 1152 5058 1170
rect 5040 1170 5058 1188
rect 5040 1188 5058 1206
rect 5040 1206 5058 1224
rect 5040 1224 5058 1242
rect 5040 1242 5058 1260
rect 5040 1260 5058 1278
rect 5040 1278 5058 1296
rect 5040 1296 5058 1314
rect 5040 1314 5058 1332
rect 5040 1332 5058 1350
rect 5040 1350 5058 1368
rect 5040 1368 5058 1386
rect 5040 1386 5058 1404
rect 5040 1404 5058 1422
rect 5040 1422 5058 1440
rect 5040 1440 5058 1458
rect 5040 1458 5058 1476
rect 5040 1476 5058 1494
rect 5040 1494 5058 1512
rect 5040 1512 5058 1530
rect 5040 1530 5058 1548
rect 5040 1548 5058 1566
rect 5040 1566 5058 1584
rect 5040 1584 5058 1602
rect 5040 1602 5058 1620
rect 5040 1620 5058 1638
rect 5040 1638 5058 1656
rect 5040 1656 5058 1674
rect 5040 1674 5058 1692
rect 5040 1692 5058 1710
rect 5040 1710 5058 1728
rect 5040 1728 5058 1746
rect 5040 1746 5058 1764
rect 5040 1764 5058 1782
rect 5040 1782 5058 1800
rect 5040 1800 5058 1818
rect 5040 1818 5058 1836
rect 5040 1836 5058 1854
rect 5040 1854 5058 1872
rect 5040 1872 5058 1890
rect 5040 1890 5058 1908
rect 5040 1908 5058 1926
rect 5040 1926 5058 1944
rect 5040 1944 5058 1962
rect 5040 1962 5058 1980
rect 5040 1980 5058 1998
rect 5040 1998 5058 2016
rect 5040 2016 5058 2034
rect 5040 2034 5058 2052
rect 5040 2052 5058 2070
rect 5040 2070 5058 2088
rect 5040 2088 5058 2106
rect 5040 2106 5058 2124
rect 5040 2124 5058 2142
rect 5040 2142 5058 2160
rect 5040 2160 5058 2178
rect 5040 2178 5058 2196
rect 5040 2196 5058 2214
rect 5040 2214 5058 2232
rect 5040 2232 5058 2250
rect 5040 2466 5058 2484
rect 5040 2484 5058 2502
rect 5040 2502 5058 2520
rect 5040 2520 5058 2538
rect 5040 2538 5058 2556
rect 5040 2556 5058 2574
rect 5040 2574 5058 2592
rect 5040 2592 5058 2610
rect 5040 2610 5058 2628
rect 5040 2628 5058 2646
rect 5040 2646 5058 2664
rect 5040 2664 5058 2682
rect 5040 2682 5058 2700
rect 5040 2700 5058 2718
rect 5040 2718 5058 2736
rect 5040 2736 5058 2754
rect 5040 2754 5058 2772
rect 5040 2772 5058 2790
rect 5040 2790 5058 2808
rect 5040 2808 5058 2826
rect 5040 2826 5058 2844
rect 5040 2844 5058 2862
rect 5040 2862 5058 2880
rect 5040 2880 5058 2898
rect 5040 2898 5058 2916
rect 5040 2916 5058 2934
rect 5040 2934 5058 2952
rect 5040 2952 5058 2970
rect 5040 2970 5058 2988
rect 5040 2988 5058 3006
rect 5040 3006 5058 3024
rect 5040 3024 5058 3042
rect 5040 3042 5058 3060
rect 5040 3060 5058 3078
rect 5040 3078 5058 3096
rect 5040 3096 5058 3114
rect 5040 3114 5058 3132
rect 5040 3132 5058 3150
rect 5040 3150 5058 3168
rect 5040 3168 5058 3186
rect 5040 3186 5058 3204
rect 5040 3204 5058 3222
rect 5040 3222 5058 3240
rect 5040 3240 5058 3258
rect 5040 3258 5058 3276
rect 5040 3276 5058 3294
rect 5040 3294 5058 3312
rect 5040 3312 5058 3330
rect 5040 3330 5058 3348
rect 5040 3348 5058 3366
rect 5040 3366 5058 3384
rect 5040 3384 5058 3402
rect 5040 3402 5058 3420
rect 5040 3420 5058 3438
rect 5040 3438 5058 3456
rect 5040 3456 5058 3474
rect 5040 3474 5058 3492
rect 5040 3492 5058 3510
rect 5040 3510 5058 3528
rect 5040 3528 5058 3546
rect 5040 3546 5058 3564
rect 5040 3564 5058 3582
rect 5040 3582 5058 3600
rect 5040 3600 5058 3618
rect 5040 3618 5058 3636
rect 5040 3636 5058 3654
rect 5040 3654 5058 3672
rect 5040 3672 5058 3690
rect 5040 3690 5058 3708
rect 5040 3708 5058 3726
rect 5040 3726 5058 3744
rect 5040 3744 5058 3762
rect 5040 3762 5058 3780
rect 5040 3780 5058 3798
rect 5040 3798 5058 3816
rect 5040 3816 5058 3834
rect 5040 3834 5058 3852
rect 5040 3852 5058 3870
rect 5040 3870 5058 3888
rect 5040 3888 5058 3906
rect 5040 3906 5058 3924
rect 5040 3924 5058 3942
rect 5040 3942 5058 3960
rect 5040 3960 5058 3978
rect 5040 3978 5058 3996
rect 5040 3996 5058 4014
rect 5040 4014 5058 4032
rect 5040 4032 5058 4050
rect 5040 4050 5058 4068
rect 5040 4068 5058 4086
rect 5040 4086 5058 4104
rect 5040 4104 5058 4122
rect 5040 4122 5058 4140
rect 5040 4140 5058 4158
rect 5040 4158 5058 4176
rect 5040 4176 5058 4194
rect 5040 4194 5058 4212
rect 5040 4212 5058 4230
rect 5040 4230 5058 4248
rect 5040 4248 5058 4266
rect 5040 4266 5058 4284
rect 5040 4284 5058 4302
rect 5040 4302 5058 4320
rect 5040 4320 5058 4338
rect 5040 4338 5058 4356
rect 5040 4356 5058 4374
rect 5040 4374 5058 4392
rect 5040 4392 5058 4410
rect 5040 4410 5058 4428
rect 5040 4644 5058 4662
rect 5040 4662 5058 4680
rect 5040 4680 5058 4698
rect 5040 4698 5058 4716
rect 5040 4716 5058 4734
rect 5040 4734 5058 4752
rect 5040 4752 5058 4770
rect 5040 4770 5058 4788
rect 5040 4788 5058 4806
rect 5040 4806 5058 4824
rect 5040 4824 5058 4842
rect 5040 4842 5058 4860
rect 5040 4860 5058 4878
rect 5040 4878 5058 4896
rect 5040 4896 5058 4914
rect 5040 4914 5058 4932
rect 5040 4932 5058 4950
rect 5040 4950 5058 4968
rect 5040 4968 5058 4986
rect 5040 4986 5058 5004
rect 5040 5004 5058 5022
rect 5040 5022 5058 5040
rect 5040 5040 5058 5058
rect 5040 5058 5058 5076
rect 5040 5076 5058 5094
rect 5040 5094 5058 5112
rect 5040 5112 5058 5130
rect 5040 5130 5058 5148
rect 5040 5148 5058 5166
rect 5040 5166 5058 5184
rect 5040 5184 5058 5202
rect 5040 5202 5058 5220
rect 5040 5220 5058 5238
rect 5040 5238 5058 5256
rect 5040 5256 5058 5274
rect 5040 5274 5058 5292
rect 5040 5292 5058 5310
rect 5040 5310 5058 5328
rect 5040 5328 5058 5346
rect 5040 5346 5058 5364
rect 5040 5364 5058 5382
rect 5040 5382 5058 5400
rect 5040 5400 5058 5418
rect 5040 5418 5058 5436
rect 5040 5436 5058 5454
rect 5040 5454 5058 5472
rect 5040 5472 5058 5490
rect 5040 5490 5058 5508
rect 5040 5508 5058 5526
rect 5040 5526 5058 5544
rect 5040 5544 5058 5562
rect 5040 5562 5058 5580
rect 5040 5580 5058 5598
rect 5040 5598 5058 5616
rect 5040 5616 5058 5634
rect 5040 5634 5058 5652
rect 5040 5652 5058 5670
rect 5040 5670 5058 5688
rect 5040 5688 5058 5706
rect 5040 5706 5058 5724
rect 5040 5724 5058 5742
rect 5040 5742 5058 5760
rect 5040 5760 5058 5778
rect 5040 5778 5058 5796
rect 5040 5796 5058 5814
rect 5040 5814 5058 5832
rect 5040 5832 5058 5850
rect 5040 5850 5058 5868
rect 5040 5868 5058 5886
rect 5040 5886 5058 5904
rect 5040 5904 5058 5922
rect 5040 5922 5058 5940
rect 5040 5940 5058 5958
rect 5040 5958 5058 5976
rect 5040 5976 5058 5994
rect 5040 5994 5058 6012
rect 5040 6012 5058 6030
rect 5040 6030 5058 6048
rect 5040 6048 5058 6066
rect 5040 6066 5058 6084
rect 5040 6084 5058 6102
rect 5040 6102 5058 6120
rect 5040 6120 5058 6138
rect 5040 6138 5058 6156
rect 5040 6156 5058 6174
rect 5040 6174 5058 6192
rect 5040 6192 5058 6210
rect 5040 6210 5058 6228
rect 5040 6228 5058 6246
rect 5040 6246 5058 6264
rect 5040 6264 5058 6282
rect 5040 6282 5058 6300
rect 5040 6300 5058 6318
rect 5040 6318 5058 6336
rect 5040 6336 5058 6354
rect 5040 6354 5058 6372
rect 5040 6372 5058 6390
rect 5040 6390 5058 6408
rect 5040 6408 5058 6426
rect 5040 6426 5058 6444
rect 5040 6444 5058 6462
rect 5040 6462 5058 6480
rect 5040 6480 5058 6498
rect 5040 6498 5058 6516
rect 5040 6516 5058 6534
rect 5040 6534 5058 6552
rect 5040 6552 5058 6570
rect 5040 6570 5058 6588
rect 5040 6588 5058 6606
rect 5040 6606 5058 6624
rect 5040 6624 5058 6642
rect 5040 6642 5058 6660
rect 5040 6660 5058 6678
rect 5040 6678 5058 6696
rect 5040 6696 5058 6714
rect 5040 6714 5058 6732
rect 5040 6732 5058 6750
rect 5040 6750 5058 6768
rect 5040 6768 5058 6786
rect 5040 6786 5058 6804
rect 5040 6804 5058 6822
rect 5040 6822 5058 6840
rect 5040 6840 5058 6858
rect 5040 6858 5058 6876
rect 5040 6876 5058 6894
rect 5040 6894 5058 6912
rect 5040 6912 5058 6930
rect 5040 6930 5058 6948
rect 5040 6948 5058 6966
rect 5040 6966 5058 6984
rect 5040 6984 5058 7002
rect 5040 7002 5058 7020
rect 5040 7020 5058 7038
rect 5040 7038 5058 7056
rect 5040 7056 5058 7074
rect 5040 7074 5058 7092
rect 5040 7092 5058 7110
rect 5040 7110 5058 7128
rect 5040 7128 5058 7146
rect 5040 7146 5058 7164
rect 5040 7164 5058 7182
rect 5040 7182 5058 7200
rect 5040 7200 5058 7218
rect 5040 7218 5058 7236
rect 5040 7236 5058 7254
rect 5040 7254 5058 7272
rect 5040 7272 5058 7290
rect 5040 7290 5058 7308
rect 5040 7308 5058 7326
rect 5040 7326 5058 7344
rect 5040 7344 5058 7362
rect 5040 7362 5058 7380
rect 5040 7380 5058 7398
rect 5040 7398 5058 7416
rect 5040 7416 5058 7434
rect 5040 7434 5058 7452
rect 5040 7452 5058 7470
rect 5040 7470 5058 7488
rect 5040 7488 5058 7506
rect 5040 7506 5058 7524
rect 5040 7524 5058 7542
rect 5040 7542 5058 7560
rect 5040 7560 5058 7578
rect 5040 7578 5058 7596
rect 5040 7596 5058 7614
rect 5040 7614 5058 7632
rect 5040 7632 5058 7650
rect 5040 7650 5058 7668
rect 5040 7668 5058 7686
rect 5040 7686 5058 7704
rect 5040 7704 5058 7722
rect 5040 7722 5058 7740
rect 5040 7740 5058 7758
rect 5040 7758 5058 7776
rect 5040 7776 5058 7794
rect 5040 7794 5058 7812
rect 5040 7812 5058 7830
rect 5040 7830 5058 7848
rect 5040 7848 5058 7866
rect 5040 7866 5058 7884
rect 5040 7884 5058 7902
rect 5058 288 5076 306
rect 5058 306 5076 324
rect 5058 324 5076 342
rect 5058 342 5076 360
rect 5058 360 5076 378
rect 5058 378 5076 396
rect 5058 396 5076 414
rect 5058 414 5076 432
rect 5058 432 5076 450
rect 5058 450 5076 468
rect 5058 468 5076 486
rect 5058 486 5076 504
rect 5058 504 5076 522
rect 5058 522 5076 540
rect 5058 540 5076 558
rect 5058 558 5076 576
rect 5058 576 5076 594
rect 5058 594 5076 612
rect 5058 612 5076 630
rect 5058 630 5076 648
rect 5058 648 5076 666
rect 5058 666 5076 684
rect 5058 684 5076 702
rect 5058 702 5076 720
rect 5058 720 5076 738
rect 5058 738 5076 756
rect 5058 882 5076 900
rect 5058 900 5076 918
rect 5058 918 5076 936
rect 5058 936 5076 954
rect 5058 954 5076 972
rect 5058 972 5076 990
rect 5058 990 5076 1008
rect 5058 1008 5076 1026
rect 5058 1026 5076 1044
rect 5058 1044 5076 1062
rect 5058 1062 5076 1080
rect 5058 1080 5076 1098
rect 5058 1098 5076 1116
rect 5058 1116 5076 1134
rect 5058 1134 5076 1152
rect 5058 1152 5076 1170
rect 5058 1170 5076 1188
rect 5058 1188 5076 1206
rect 5058 1206 5076 1224
rect 5058 1224 5076 1242
rect 5058 1242 5076 1260
rect 5058 1260 5076 1278
rect 5058 1278 5076 1296
rect 5058 1296 5076 1314
rect 5058 1314 5076 1332
rect 5058 1332 5076 1350
rect 5058 1350 5076 1368
rect 5058 1368 5076 1386
rect 5058 1386 5076 1404
rect 5058 1404 5076 1422
rect 5058 1422 5076 1440
rect 5058 1440 5076 1458
rect 5058 1458 5076 1476
rect 5058 1476 5076 1494
rect 5058 1494 5076 1512
rect 5058 1512 5076 1530
rect 5058 1530 5076 1548
rect 5058 1548 5076 1566
rect 5058 1566 5076 1584
rect 5058 1584 5076 1602
rect 5058 1602 5076 1620
rect 5058 1620 5076 1638
rect 5058 1638 5076 1656
rect 5058 1656 5076 1674
rect 5058 1674 5076 1692
rect 5058 1692 5076 1710
rect 5058 1710 5076 1728
rect 5058 1728 5076 1746
rect 5058 1746 5076 1764
rect 5058 1764 5076 1782
rect 5058 1782 5076 1800
rect 5058 1800 5076 1818
rect 5058 1818 5076 1836
rect 5058 1836 5076 1854
rect 5058 1854 5076 1872
rect 5058 1872 5076 1890
rect 5058 1890 5076 1908
rect 5058 1908 5076 1926
rect 5058 1926 5076 1944
rect 5058 1944 5076 1962
rect 5058 1962 5076 1980
rect 5058 1980 5076 1998
rect 5058 1998 5076 2016
rect 5058 2016 5076 2034
rect 5058 2034 5076 2052
rect 5058 2052 5076 2070
rect 5058 2070 5076 2088
rect 5058 2088 5076 2106
rect 5058 2106 5076 2124
rect 5058 2124 5076 2142
rect 5058 2142 5076 2160
rect 5058 2160 5076 2178
rect 5058 2178 5076 2196
rect 5058 2196 5076 2214
rect 5058 2214 5076 2232
rect 5058 2232 5076 2250
rect 5058 2250 5076 2268
rect 5058 2484 5076 2502
rect 5058 2502 5076 2520
rect 5058 2520 5076 2538
rect 5058 2538 5076 2556
rect 5058 2556 5076 2574
rect 5058 2574 5076 2592
rect 5058 2592 5076 2610
rect 5058 2610 5076 2628
rect 5058 2628 5076 2646
rect 5058 2646 5076 2664
rect 5058 2664 5076 2682
rect 5058 2682 5076 2700
rect 5058 2700 5076 2718
rect 5058 2718 5076 2736
rect 5058 2736 5076 2754
rect 5058 2754 5076 2772
rect 5058 2772 5076 2790
rect 5058 2790 5076 2808
rect 5058 2808 5076 2826
rect 5058 2826 5076 2844
rect 5058 2844 5076 2862
rect 5058 2862 5076 2880
rect 5058 2880 5076 2898
rect 5058 2898 5076 2916
rect 5058 2916 5076 2934
rect 5058 2934 5076 2952
rect 5058 2952 5076 2970
rect 5058 2970 5076 2988
rect 5058 2988 5076 3006
rect 5058 3006 5076 3024
rect 5058 3024 5076 3042
rect 5058 3042 5076 3060
rect 5058 3060 5076 3078
rect 5058 3078 5076 3096
rect 5058 3096 5076 3114
rect 5058 3114 5076 3132
rect 5058 3132 5076 3150
rect 5058 3150 5076 3168
rect 5058 3168 5076 3186
rect 5058 3186 5076 3204
rect 5058 3204 5076 3222
rect 5058 3222 5076 3240
rect 5058 3240 5076 3258
rect 5058 3258 5076 3276
rect 5058 3276 5076 3294
rect 5058 3294 5076 3312
rect 5058 3312 5076 3330
rect 5058 3330 5076 3348
rect 5058 3348 5076 3366
rect 5058 3366 5076 3384
rect 5058 3384 5076 3402
rect 5058 3402 5076 3420
rect 5058 3420 5076 3438
rect 5058 3438 5076 3456
rect 5058 3456 5076 3474
rect 5058 3474 5076 3492
rect 5058 3492 5076 3510
rect 5058 3510 5076 3528
rect 5058 3528 5076 3546
rect 5058 3546 5076 3564
rect 5058 3564 5076 3582
rect 5058 3582 5076 3600
rect 5058 3600 5076 3618
rect 5058 3618 5076 3636
rect 5058 3636 5076 3654
rect 5058 3654 5076 3672
rect 5058 3672 5076 3690
rect 5058 3690 5076 3708
rect 5058 3708 5076 3726
rect 5058 3726 5076 3744
rect 5058 3744 5076 3762
rect 5058 3762 5076 3780
rect 5058 3780 5076 3798
rect 5058 3798 5076 3816
rect 5058 3816 5076 3834
rect 5058 3834 5076 3852
rect 5058 3852 5076 3870
rect 5058 3870 5076 3888
rect 5058 3888 5076 3906
rect 5058 3906 5076 3924
rect 5058 3924 5076 3942
rect 5058 3942 5076 3960
rect 5058 3960 5076 3978
rect 5058 3978 5076 3996
rect 5058 3996 5076 4014
rect 5058 4014 5076 4032
rect 5058 4032 5076 4050
rect 5058 4050 5076 4068
rect 5058 4068 5076 4086
rect 5058 4086 5076 4104
rect 5058 4104 5076 4122
rect 5058 4122 5076 4140
rect 5058 4140 5076 4158
rect 5058 4158 5076 4176
rect 5058 4176 5076 4194
rect 5058 4194 5076 4212
rect 5058 4212 5076 4230
rect 5058 4230 5076 4248
rect 5058 4248 5076 4266
rect 5058 4266 5076 4284
rect 5058 4284 5076 4302
rect 5058 4302 5076 4320
rect 5058 4320 5076 4338
rect 5058 4338 5076 4356
rect 5058 4356 5076 4374
rect 5058 4374 5076 4392
rect 5058 4392 5076 4410
rect 5058 4410 5076 4428
rect 5058 4428 5076 4446
rect 5058 4662 5076 4680
rect 5058 4680 5076 4698
rect 5058 4698 5076 4716
rect 5058 4716 5076 4734
rect 5058 4734 5076 4752
rect 5058 4752 5076 4770
rect 5058 4770 5076 4788
rect 5058 4788 5076 4806
rect 5058 4806 5076 4824
rect 5058 4824 5076 4842
rect 5058 4842 5076 4860
rect 5058 4860 5076 4878
rect 5058 4878 5076 4896
rect 5058 4896 5076 4914
rect 5058 4914 5076 4932
rect 5058 4932 5076 4950
rect 5058 4950 5076 4968
rect 5058 4968 5076 4986
rect 5058 4986 5076 5004
rect 5058 5004 5076 5022
rect 5058 5022 5076 5040
rect 5058 5040 5076 5058
rect 5058 5058 5076 5076
rect 5058 5076 5076 5094
rect 5058 5094 5076 5112
rect 5058 5112 5076 5130
rect 5058 5130 5076 5148
rect 5058 5148 5076 5166
rect 5058 5166 5076 5184
rect 5058 5184 5076 5202
rect 5058 5202 5076 5220
rect 5058 5220 5076 5238
rect 5058 5238 5076 5256
rect 5058 5256 5076 5274
rect 5058 5274 5076 5292
rect 5058 5292 5076 5310
rect 5058 5310 5076 5328
rect 5058 5328 5076 5346
rect 5058 5346 5076 5364
rect 5058 5364 5076 5382
rect 5058 5382 5076 5400
rect 5058 5400 5076 5418
rect 5058 5418 5076 5436
rect 5058 5436 5076 5454
rect 5058 5454 5076 5472
rect 5058 5472 5076 5490
rect 5058 5490 5076 5508
rect 5058 5508 5076 5526
rect 5058 5526 5076 5544
rect 5058 5544 5076 5562
rect 5058 5562 5076 5580
rect 5058 5580 5076 5598
rect 5058 5598 5076 5616
rect 5058 5616 5076 5634
rect 5058 5634 5076 5652
rect 5058 5652 5076 5670
rect 5058 5670 5076 5688
rect 5058 5688 5076 5706
rect 5058 5706 5076 5724
rect 5058 5724 5076 5742
rect 5058 5742 5076 5760
rect 5058 5760 5076 5778
rect 5058 5778 5076 5796
rect 5058 5796 5076 5814
rect 5058 5814 5076 5832
rect 5058 5832 5076 5850
rect 5058 5850 5076 5868
rect 5058 5868 5076 5886
rect 5058 5886 5076 5904
rect 5058 5904 5076 5922
rect 5058 5922 5076 5940
rect 5058 5940 5076 5958
rect 5058 5958 5076 5976
rect 5058 5976 5076 5994
rect 5058 5994 5076 6012
rect 5058 6012 5076 6030
rect 5058 6030 5076 6048
rect 5058 6048 5076 6066
rect 5058 6066 5076 6084
rect 5058 6084 5076 6102
rect 5058 6102 5076 6120
rect 5058 6120 5076 6138
rect 5058 6138 5076 6156
rect 5058 6156 5076 6174
rect 5058 6174 5076 6192
rect 5058 6192 5076 6210
rect 5058 6210 5076 6228
rect 5058 6228 5076 6246
rect 5058 6246 5076 6264
rect 5058 6264 5076 6282
rect 5058 6282 5076 6300
rect 5058 6300 5076 6318
rect 5058 6318 5076 6336
rect 5058 6336 5076 6354
rect 5058 6354 5076 6372
rect 5058 6372 5076 6390
rect 5058 6390 5076 6408
rect 5058 6408 5076 6426
rect 5058 6426 5076 6444
rect 5058 6444 5076 6462
rect 5058 6462 5076 6480
rect 5058 6480 5076 6498
rect 5058 6498 5076 6516
rect 5058 6516 5076 6534
rect 5058 6534 5076 6552
rect 5058 6552 5076 6570
rect 5058 6570 5076 6588
rect 5058 6588 5076 6606
rect 5058 6606 5076 6624
rect 5058 6624 5076 6642
rect 5058 6642 5076 6660
rect 5058 6660 5076 6678
rect 5058 6678 5076 6696
rect 5058 6696 5076 6714
rect 5058 6714 5076 6732
rect 5058 6732 5076 6750
rect 5058 6750 5076 6768
rect 5058 6768 5076 6786
rect 5058 6786 5076 6804
rect 5058 6804 5076 6822
rect 5058 6822 5076 6840
rect 5058 6840 5076 6858
rect 5058 6858 5076 6876
rect 5058 6876 5076 6894
rect 5058 6894 5076 6912
rect 5058 6912 5076 6930
rect 5058 6930 5076 6948
rect 5058 6948 5076 6966
rect 5058 6966 5076 6984
rect 5058 6984 5076 7002
rect 5058 7002 5076 7020
rect 5058 7020 5076 7038
rect 5058 7038 5076 7056
rect 5058 7056 5076 7074
rect 5058 7074 5076 7092
rect 5058 7092 5076 7110
rect 5058 7110 5076 7128
rect 5058 7128 5076 7146
rect 5058 7146 5076 7164
rect 5058 7164 5076 7182
rect 5058 7182 5076 7200
rect 5058 7200 5076 7218
rect 5058 7218 5076 7236
rect 5058 7236 5076 7254
rect 5058 7254 5076 7272
rect 5058 7272 5076 7290
rect 5058 7290 5076 7308
rect 5058 7308 5076 7326
rect 5058 7326 5076 7344
rect 5058 7344 5076 7362
rect 5058 7362 5076 7380
rect 5058 7380 5076 7398
rect 5058 7398 5076 7416
rect 5058 7416 5076 7434
rect 5058 7434 5076 7452
rect 5058 7452 5076 7470
rect 5058 7470 5076 7488
rect 5058 7488 5076 7506
rect 5058 7506 5076 7524
rect 5058 7524 5076 7542
rect 5058 7542 5076 7560
rect 5058 7560 5076 7578
rect 5058 7578 5076 7596
rect 5058 7596 5076 7614
rect 5058 7614 5076 7632
rect 5058 7632 5076 7650
rect 5058 7650 5076 7668
rect 5058 7668 5076 7686
rect 5058 7686 5076 7704
rect 5058 7704 5076 7722
rect 5058 7722 5076 7740
rect 5058 7740 5076 7758
rect 5058 7758 5076 7776
rect 5058 7776 5076 7794
rect 5058 7794 5076 7812
rect 5058 7812 5076 7830
rect 5058 7830 5076 7848
rect 5058 7848 5076 7866
rect 5058 7866 5076 7884
rect 5058 7884 5076 7902
rect 5058 7902 5076 7920
rect 5058 7920 5076 7938
rect 5076 288 5094 306
rect 5076 306 5094 324
rect 5076 324 5094 342
rect 5076 342 5094 360
rect 5076 360 5094 378
rect 5076 378 5094 396
rect 5076 396 5094 414
rect 5076 414 5094 432
rect 5076 432 5094 450
rect 5076 450 5094 468
rect 5076 468 5094 486
rect 5076 486 5094 504
rect 5076 504 5094 522
rect 5076 522 5094 540
rect 5076 540 5094 558
rect 5076 558 5094 576
rect 5076 576 5094 594
rect 5076 594 5094 612
rect 5076 612 5094 630
rect 5076 630 5094 648
rect 5076 648 5094 666
rect 5076 666 5094 684
rect 5076 684 5094 702
rect 5076 702 5094 720
rect 5076 720 5094 738
rect 5076 738 5094 756
rect 5076 882 5094 900
rect 5076 900 5094 918
rect 5076 918 5094 936
rect 5076 936 5094 954
rect 5076 954 5094 972
rect 5076 972 5094 990
rect 5076 990 5094 1008
rect 5076 1008 5094 1026
rect 5076 1026 5094 1044
rect 5076 1044 5094 1062
rect 5076 1062 5094 1080
rect 5076 1080 5094 1098
rect 5076 1098 5094 1116
rect 5076 1116 5094 1134
rect 5076 1134 5094 1152
rect 5076 1152 5094 1170
rect 5076 1170 5094 1188
rect 5076 1188 5094 1206
rect 5076 1206 5094 1224
rect 5076 1224 5094 1242
rect 5076 1242 5094 1260
rect 5076 1260 5094 1278
rect 5076 1278 5094 1296
rect 5076 1296 5094 1314
rect 5076 1314 5094 1332
rect 5076 1332 5094 1350
rect 5076 1350 5094 1368
rect 5076 1368 5094 1386
rect 5076 1386 5094 1404
rect 5076 1404 5094 1422
rect 5076 1422 5094 1440
rect 5076 1440 5094 1458
rect 5076 1458 5094 1476
rect 5076 1476 5094 1494
rect 5076 1494 5094 1512
rect 5076 1512 5094 1530
rect 5076 1530 5094 1548
rect 5076 1548 5094 1566
rect 5076 1566 5094 1584
rect 5076 1584 5094 1602
rect 5076 1602 5094 1620
rect 5076 1620 5094 1638
rect 5076 1638 5094 1656
rect 5076 1656 5094 1674
rect 5076 1674 5094 1692
rect 5076 1692 5094 1710
rect 5076 1710 5094 1728
rect 5076 1728 5094 1746
rect 5076 1746 5094 1764
rect 5076 1764 5094 1782
rect 5076 1782 5094 1800
rect 5076 1800 5094 1818
rect 5076 1818 5094 1836
rect 5076 1836 5094 1854
rect 5076 1854 5094 1872
rect 5076 1872 5094 1890
rect 5076 1890 5094 1908
rect 5076 1908 5094 1926
rect 5076 1926 5094 1944
rect 5076 1944 5094 1962
rect 5076 1962 5094 1980
rect 5076 1980 5094 1998
rect 5076 1998 5094 2016
rect 5076 2016 5094 2034
rect 5076 2034 5094 2052
rect 5076 2052 5094 2070
rect 5076 2070 5094 2088
rect 5076 2088 5094 2106
rect 5076 2106 5094 2124
rect 5076 2124 5094 2142
rect 5076 2142 5094 2160
rect 5076 2160 5094 2178
rect 5076 2178 5094 2196
rect 5076 2196 5094 2214
rect 5076 2214 5094 2232
rect 5076 2232 5094 2250
rect 5076 2250 5094 2268
rect 5076 2484 5094 2502
rect 5076 2502 5094 2520
rect 5076 2520 5094 2538
rect 5076 2538 5094 2556
rect 5076 2556 5094 2574
rect 5076 2574 5094 2592
rect 5076 2592 5094 2610
rect 5076 2610 5094 2628
rect 5076 2628 5094 2646
rect 5076 2646 5094 2664
rect 5076 2664 5094 2682
rect 5076 2682 5094 2700
rect 5076 2700 5094 2718
rect 5076 2718 5094 2736
rect 5076 2736 5094 2754
rect 5076 2754 5094 2772
rect 5076 2772 5094 2790
rect 5076 2790 5094 2808
rect 5076 2808 5094 2826
rect 5076 2826 5094 2844
rect 5076 2844 5094 2862
rect 5076 2862 5094 2880
rect 5076 2880 5094 2898
rect 5076 2898 5094 2916
rect 5076 2916 5094 2934
rect 5076 2934 5094 2952
rect 5076 2952 5094 2970
rect 5076 2970 5094 2988
rect 5076 2988 5094 3006
rect 5076 3006 5094 3024
rect 5076 3024 5094 3042
rect 5076 3042 5094 3060
rect 5076 3060 5094 3078
rect 5076 3078 5094 3096
rect 5076 3096 5094 3114
rect 5076 3114 5094 3132
rect 5076 3132 5094 3150
rect 5076 3150 5094 3168
rect 5076 3168 5094 3186
rect 5076 3186 5094 3204
rect 5076 3204 5094 3222
rect 5076 3222 5094 3240
rect 5076 3240 5094 3258
rect 5076 3258 5094 3276
rect 5076 3276 5094 3294
rect 5076 3294 5094 3312
rect 5076 3312 5094 3330
rect 5076 3330 5094 3348
rect 5076 3348 5094 3366
rect 5076 3366 5094 3384
rect 5076 3384 5094 3402
rect 5076 3402 5094 3420
rect 5076 3420 5094 3438
rect 5076 3438 5094 3456
rect 5076 3456 5094 3474
rect 5076 3474 5094 3492
rect 5076 3492 5094 3510
rect 5076 3510 5094 3528
rect 5076 3528 5094 3546
rect 5076 3546 5094 3564
rect 5076 3564 5094 3582
rect 5076 3582 5094 3600
rect 5076 3600 5094 3618
rect 5076 3618 5094 3636
rect 5076 3636 5094 3654
rect 5076 3654 5094 3672
rect 5076 3672 5094 3690
rect 5076 3690 5094 3708
rect 5076 3708 5094 3726
rect 5076 3726 5094 3744
rect 5076 3744 5094 3762
rect 5076 3762 5094 3780
rect 5076 3780 5094 3798
rect 5076 3798 5094 3816
rect 5076 3816 5094 3834
rect 5076 3834 5094 3852
rect 5076 3852 5094 3870
rect 5076 3870 5094 3888
rect 5076 3888 5094 3906
rect 5076 3906 5094 3924
rect 5076 3924 5094 3942
rect 5076 3942 5094 3960
rect 5076 3960 5094 3978
rect 5076 3978 5094 3996
rect 5076 3996 5094 4014
rect 5076 4014 5094 4032
rect 5076 4032 5094 4050
rect 5076 4050 5094 4068
rect 5076 4068 5094 4086
rect 5076 4086 5094 4104
rect 5076 4104 5094 4122
rect 5076 4122 5094 4140
rect 5076 4140 5094 4158
rect 5076 4158 5094 4176
rect 5076 4176 5094 4194
rect 5076 4194 5094 4212
rect 5076 4212 5094 4230
rect 5076 4230 5094 4248
rect 5076 4248 5094 4266
rect 5076 4266 5094 4284
rect 5076 4284 5094 4302
rect 5076 4302 5094 4320
rect 5076 4320 5094 4338
rect 5076 4338 5094 4356
rect 5076 4356 5094 4374
rect 5076 4374 5094 4392
rect 5076 4392 5094 4410
rect 5076 4410 5094 4428
rect 5076 4428 5094 4446
rect 5076 4446 5094 4464
rect 5076 4680 5094 4698
rect 5076 4698 5094 4716
rect 5076 4716 5094 4734
rect 5076 4734 5094 4752
rect 5076 4752 5094 4770
rect 5076 4770 5094 4788
rect 5076 4788 5094 4806
rect 5076 4806 5094 4824
rect 5076 4824 5094 4842
rect 5076 4842 5094 4860
rect 5076 4860 5094 4878
rect 5076 4878 5094 4896
rect 5076 4896 5094 4914
rect 5076 4914 5094 4932
rect 5076 4932 5094 4950
rect 5076 4950 5094 4968
rect 5076 4968 5094 4986
rect 5076 4986 5094 5004
rect 5076 5004 5094 5022
rect 5076 5022 5094 5040
rect 5076 5040 5094 5058
rect 5076 5058 5094 5076
rect 5076 5076 5094 5094
rect 5076 5094 5094 5112
rect 5076 5112 5094 5130
rect 5076 5130 5094 5148
rect 5076 5148 5094 5166
rect 5076 5166 5094 5184
rect 5076 5184 5094 5202
rect 5076 5202 5094 5220
rect 5076 5220 5094 5238
rect 5076 5238 5094 5256
rect 5076 5256 5094 5274
rect 5076 5274 5094 5292
rect 5076 5292 5094 5310
rect 5076 5310 5094 5328
rect 5076 5328 5094 5346
rect 5076 5346 5094 5364
rect 5076 5364 5094 5382
rect 5076 5382 5094 5400
rect 5076 5400 5094 5418
rect 5076 5418 5094 5436
rect 5076 5436 5094 5454
rect 5076 5454 5094 5472
rect 5076 5472 5094 5490
rect 5076 5490 5094 5508
rect 5076 5508 5094 5526
rect 5076 5526 5094 5544
rect 5076 5544 5094 5562
rect 5076 5562 5094 5580
rect 5076 5580 5094 5598
rect 5076 5598 5094 5616
rect 5076 5616 5094 5634
rect 5076 5634 5094 5652
rect 5076 5652 5094 5670
rect 5076 5670 5094 5688
rect 5076 5688 5094 5706
rect 5076 5706 5094 5724
rect 5076 5724 5094 5742
rect 5076 5742 5094 5760
rect 5076 5760 5094 5778
rect 5076 5778 5094 5796
rect 5076 5796 5094 5814
rect 5076 5814 5094 5832
rect 5076 5832 5094 5850
rect 5076 5850 5094 5868
rect 5076 5868 5094 5886
rect 5076 5886 5094 5904
rect 5076 5904 5094 5922
rect 5076 5922 5094 5940
rect 5076 5940 5094 5958
rect 5076 5958 5094 5976
rect 5076 5976 5094 5994
rect 5076 5994 5094 6012
rect 5076 6012 5094 6030
rect 5076 6030 5094 6048
rect 5076 6048 5094 6066
rect 5076 6066 5094 6084
rect 5076 6084 5094 6102
rect 5076 6102 5094 6120
rect 5076 6120 5094 6138
rect 5076 6138 5094 6156
rect 5076 6156 5094 6174
rect 5076 6174 5094 6192
rect 5076 6192 5094 6210
rect 5076 6210 5094 6228
rect 5076 6228 5094 6246
rect 5076 6246 5094 6264
rect 5076 6264 5094 6282
rect 5076 6282 5094 6300
rect 5076 6300 5094 6318
rect 5076 6318 5094 6336
rect 5076 6336 5094 6354
rect 5076 6354 5094 6372
rect 5076 6372 5094 6390
rect 5076 6390 5094 6408
rect 5076 6408 5094 6426
rect 5076 6426 5094 6444
rect 5076 6444 5094 6462
rect 5076 6462 5094 6480
rect 5076 6480 5094 6498
rect 5076 6498 5094 6516
rect 5076 6516 5094 6534
rect 5076 6534 5094 6552
rect 5076 6552 5094 6570
rect 5076 6570 5094 6588
rect 5076 6588 5094 6606
rect 5076 6606 5094 6624
rect 5076 6624 5094 6642
rect 5076 6642 5094 6660
rect 5076 6660 5094 6678
rect 5076 6678 5094 6696
rect 5076 6696 5094 6714
rect 5076 6714 5094 6732
rect 5076 6732 5094 6750
rect 5076 6750 5094 6768
rect 5076 6768 5094 6786
rect 5076 6786 5094 6804
rect 5076 6804 5094 6822
rect 5076 6822 5094 6840
rect 5076 6840 5094 6858
rect 5076 6858 5094 6876
rect 5076 6876 5094 6894
rect 5076 6894 5094 6912
rect 5076 6912 5094 6930
rect 5076 6930 5094 6948
rect 5076 6948 5094 6966
rect 5076 6966 5094 6984
rect 5076 6984 5094 7002
rect 5076 7002 5094 7020
rect 5076 7020 5094 7038
rect 5076 7038 5094 7056
rect 5076 7056 5094 7074
rect 5076 7074 5094 7092
rect 5076 7092 5094 7110
rect 5076 7110 5094 7128
rect 5076 7128 5094 7146
rect 5076 7146 5094 7164
rect 5076 7164 5094 7182
rect 5076 7182 5094 7200
rect 5076 7200 5094 7218
rect 5076 7218 5094 7236
rect 5076 7236 5094 7254
rect 5076 7254 5094 7272
rect 5076 7272 5094 7290
rect 5076 7290 5094 7308
rect 5076 7308 5094 7326
rect 5076 7326 5094 7344
rect 5076 7344 5094 7362
rect 5076 7362 5094 7380
rect 5076 7380 5094 7398
rect 5076 7398 5094 7416
rect 5076 7416 5094 7434
rect 5076 7434 5094 7452
rect 5076 7452 5094 7470
rect 5076 7470 5094 7488
rect 5076 7488 5094 7506
rect 5076 7506 5094 7524
rect 5076 7524 5094 7542
rect 5076 7542 5094 7560
rect 5076 7560 5094 7578
rect 5076 7578 5094 7596
rect 5076 7596 5094 7614
rect 5076 7614 5094 7632
rect 5076 7632 5094 7650
rect 5076 7650 5094 7668
rect 5076 7668 5094 7686
rect 5076 7686 5094 7704
rect 5076 7704 5094 7722
rect 5076 7722 5094 7740
rect 5076 7740 5094 7758
rect 5076 7758 5094 7776
rect 5076 7776 5094 7794
rect 5076 7794 5094 7812
rect 5076 7812 5094 7830
rect 5076 7830 5094 7848
rect 5076 7848 5094 7866
rect 5076 7866 5094 7884
rect 5076 7884 5094 7902
rect 5076 7902 5094 7920
rect 5076 7920 5094 7938
rect 5076 7938 5094 7956
rect 5094 306 5112 324
rect 5094 324 5112 342
rect 5094 342 5112 360
rect 5094 360 5112 378
rect 5094 378 5112 396
rect 5094 396 5112 414
rect 5094 414 5112 432
rect 5094 432 5112 450
rect 5094 450 5112 468
rect 5094 468 5112 486
rect 5094 486 5112 504
rect 5094 504 5112 522
rect 5094 522 5112 540
rect 5094 540 5112 558
rect 5094 558 5112 576
rect 5094 576 5112 594
rect 5094 594 5112 612
rect 5094 612 5112 630
rect 5094 630 5112 648
rect 5094 648 5112 666
rect 5094 666 5112 684
rect 5094 684 5112 702
rect 5094 702 5112 720
rect 5094 720 5112 738
rect 5094 738 5112 756
rect 5094 756 5112 774
rect 5094 900 5112 918
rect 5094 918 5112 936
rect 5094 936 5112 954
rect 5094 954 5112 972
rect 5094 972 5112 990
rect 5094 990 5112 1008
rect 5094 1008 5112 1026
rect 5094 1026 5112 1044
rect 5094 1044 5112 1062
rect 5094 1062 5112 1080
rect 5094 1080 5112 1098
rect 5094 1098 5112 1116
rect 5094 1116 5112 1134
rect 5094 1134 5112 1152
rect 5094 1152 5112 1170
rect 5094 1170 5112 1188
rect 5094 1188 5112 1206
rect 5094 1206 5112 1224
rect 5094 1224 5112 1242
rect 5094 1242 5112 1260
rect 5094 1260 5112 1278
rect 5094 1278 5112 1296
rect 5094 1296 5112 1314
rect 5094 1314 5112 1332
rect 5094 1332 5112 1350
rect 5094 1350 5112 1368
rect 5094 1368 5112 1386
rect 5094 1386 5112 1404
rect 5094 1404 5112 1422
rect 5094 1422 5112 1440
rect 5094 1440 5112 1458
rect 5094 1458 5112 1476
rect 5094 1476 5112 1494
rect 5094 1494 5112 1512
rect 5094 1512 5112 1530
rect 5094 1530 5112 1548
rect 5094 1548 5112 1566
rect 5094 1566 5112 1584
rect 5094 1584 5112 1602
rect 5094 1602 5112 1620
rect 5094 1620 5112 1638
rect 5094 1638 5112 1656
rect 5094 1656 5112 1674
rect 5094 1674 5112 1692
rect 5094 1692 5112 1710
rect 5094 1710 5112 1728
rect 5094 1728 5112 1746
rect 5094 1746 5112 1764
rect 5094 1764 5112 1782
rect 5094 1782 5112 1800
rect 5094 1800 5112 1818
rect 5094 1818 5112 1836
rect 5094 1836 5112 1854
rect 5094 1854 5112 1872
rect 5094 1872 5112 1890
rect 5094 1890 5112 1908
rect 5094 1908 5112 1926
rect 5094 1926 5112 1944
rect 5094 1944 5112 1962
rect 5094 1962 5112 1980
rect 5094 1980 5112 1998
rect 5094 1998 5112 2016
rect 5094 2016 5112 2034
rect 5094 2034 5112 2052
rect 5094 2052 5112 2070
rect 5094 2070 5112 2088
rect 5094 2088 5112 2106
rect 5094 2106 5112 2124
rect 5094 2124 5112 2142
rect 5094 2142 5112 2160
rect 5094 2160 5112 2178
rect 5094 2178 5112 2196
rect 5094 2196 5112 2214
rect 5094 2214 5112 2232
rect 5094 2232 5112 2250
rect 5094 2250 5112 2268
rect 5094 2268 5112 2286
rect 5094 2502 5112 2520
rect 5094 2520 5112 2538
rect 5094 2538 5112 2556
rect 5094 2556 5112 2574
rect 5094 2574 5112 2592
rect 5094 2592 5112 2610
rect 5094 2610 5112 2628
rect 5094 2628 5112 2646
rect 5094 2646 5112 2664
rect 5094 2664 5112 2682
rect 5094 2682 5112 2700
rect 5094 2700 5112 2718
rect 5094 2718 5112 2736
rect 5094 2736 5112 2754
rect 5094 2754 5112 2772
rect 5094 2772 5112 2790
rect 5094 2790 5112 2808
rect 5094 2808 5112 2826
rect 5094 2826 5112 2844
rect 5094 2844 5112 2862
rect 5094 2862 5112 2880
rect 5094 2880 5112 2898
rect 5094 2898 5112 2916
rect 5094 2916 5112 2934
rect 5094 2934 5112 2952
rect 5094 2952 5112 2970
rect 5094 2970 5112 2988
rect 5094 2988 5112 3006
rect 5094 3006 5112 3024
rect 5094 3024 5112 3042
rect 5094 3042 5112 3060
rect 5094 3060 5112 3078
rect 5094 3078 5112 3096
rect 5094 3096 5112 3114
rect 5094 3114 5112 3132
rect 5094 3132 5112 3150
rect 5094 3150 5112 3168
rect 5094 3168 5112 3186
rect 5094 3186 5112 3204
rect 5094 3204 5112 3222
rect 5094 3222 5112 3240
rect 5094 3240 5112 3258
rect 5094 3258 5112 3276
rect 5094 3276 5112 3294
rect 5094 3294 5112 3312
rect 5094 3312 5112 3330
rect 5094 3330 5112 3348
rect 5094 3348 5112 3366
rect 5094 3366 5112 3384
rect 5094 3384 5112 3402
rect 5094 3402 5112 3420
rect 5094 3420 5112 3438
rect 5094 3438 5112 3456
rect 5094 3456 5112 3474
rect 5094 3474 5112 3492
rect 5094 3492 5112 3510
rect 5094 3510 5112 3528
rect 5094 3528 5112 3546
rect 5094 3546 5112 3564
rect 5094 3564 5112 3582
rect 5094 3582 5112 3600
rect 5094 3600 5112 3618
rect 5094 3618 5112 3636
rect 5094 3636 5112 3654
rect 5094 3654 5112 3672
rect 5094 3672 5112 3690
rect 5094 3690 5112 3708
rect 5094 3708 5112 3726
rect 5094 3726 5112 3744
rect 5094 3744 5112 3762
rect 5094 3762 5112 3780
rect 5094 3780 5112 3798
rect 5094 3798 5112 3816
rect 5094 3816 5112 3834
rect 5094 3834 5112 3852
rect 5094 3852 5112 3870
rect 5094 3870 5112 3888
rect 5094 3888 5112 3906
rect 5094 3906 5112 3924
rect 5094 3924 5112 3942
rect 5094 3942 5112 3960
rect 5094 3960 5112 3978
rect 5094 3978 5112 3996
rect 5094 3996 5112 4014
rect 5094 4014 5112 4032
rect 5094 4032 5112 4050
rect 5094 4050 5112 4068
rect 5094 4068 5112 4086
rect 5094 4086 5112 4104
rect 5094 4104 5112 4122
rect 5094 4122 5112 4140
rect 5094 4140 5112 4158
rect 5094 4158 5112 4176
rect 5094 4176 5112 4194
rect 5094 4194 5112 4212
rect 5094 4212 5112 4230
rect 5094 4230 5112 4248
rect 5094 4248 5112 4266
rect 5094 4266 5112 4284
rect 5094 4284 5112 4302
rect 5094 4302 5112 4320
rect 5094 4320 5112 4338
rect 5094 4338 5112 4356
rect 5094 4356 5112 4374
rect 5094 4374 5112 4392
rect 5094 4392 5112 4410
rect 5094 4410 5112 4428
rect 5094 4428 5112 4446
rect 5094 4446 5112 4464
rect 5094 4464 5112 4482
rect 5094 4698 5112 4716
rect 5094 4716 5112 4734
rect 5094 4734 5112 4752
rect 5094 4752 5112 4770
rect 5094 4770 5112 4788
rect 5094 4788 5112 4806
rect 5094 4806 5112 4824
rect 5094 4824 5112 4842
rect 5094 4842 5112 4860
rect 5094 4860 5112 4878
rect 5094 4878 5112 4896
rect 5094 4896 5112 4914
rect 5094 4914 5112 4932
rect 5094 4932 5112 4950
rect 5094 4950 5112 4968
rect 5094 4968 5112 4986
rect 5094 4986 5112 5004
rect 5094 5004 5112 5022
rect 5094 5022 5112 5040
rect 5094 5040 5112 5058
rect 5094 5058 5112 5076
rect 5094 5076 5112 5094
rect 5094 5094 5112 5112
rect 5094 5112 5112 5130
rect 5094 5130 5112 5148
rect 5094 5148 5112 5166
rect 5094 5166 5112 5184
rect 5094 5184 5112 5202
rect 5094 5202 5112 5220
rect 5094 5220 5112 5238
rect 5094 5238 5112 5256
rect 5094 5256 5112 5274
rect 5094 5274 5112 5292
rect 5094 5292 5112 5310
rect 5094 5310 5112 5328
rect 5094 5328 5112 5346
rect 5094 5346 5112 5364
rect 5094 5364 5112 5382
rect 5094 5382 5112 5400
rect 5094 5400 5112 5418
rect 5094 5418 5112 5436
rect 5094 5436 5112 5454
rect 5094 5454 5112 5472
rect 5094 5472 5112 5490
rect 5094 5490 5112 5508
rect 5094 5508 5112 5526
rect 5094 5526 5112 5544
rect 5094 5544 5112 5562
rect 5094 5562 5112 5580
rect 5094 5580 5112 5598
rect 5094 5598 5112 5616
rect 5094 5616 5112 5634
rect 5094 5634 5112 5652
rect 5094 5652 5112 5670
rect 5094 5670 5112 5688
rect 5094 5688 5112 5706
rect 5094 5706 5112 5724
rect 5094 5724 5112 5742
rect 5094 5742 5112 5760
rect 5094 5760 5112 5778
rect 5094 5778 5112 5796
rect 5094 5796 5112 5814
rect 5094 5814 5112 5832
rect 5094 5832 5112 5850
rect 5094 5850 5112 5868
rect 5094 5868 5112 5886
rect 5094 5886 5112 5904
rect 5094 5904 5112 5922
rect 5094 5922 5112 5940
rect 5094 5940 5112 5958
rect 5094 5958 5112 5976
rect 5094 5976 5112 5994
rect 5094 5994 5112 6012
rect 5094 6012 5112 6030
rect 5094 6030 5112 6048
rect 5094 6048 5112 6066
rect 5094 6066 5112 6084
rect 5094 6084 5112 6102
rect 5094 6102 5112 6120
rect 5094 6120 5112 6138
rect 5094 6138 5112 6156
rect 5094 6156 5112 6174
rect 5094 6174 5112 6192
rect 5094 6192 5112 6210
rect 5094 6210 5112 6228
rect 5094 6228 5112 6246
rect 5094 6246 5112 6264
rect 5094 6264 5112 6282
rect 5094 6282 5112 6300
rect 5094 6300 5112 6318
rect 5094 6318 5112 6336
rect 5094 6336 5112 6354
rect 5094 6354 5112 6372
rect 5094 6372 5112 6390
rect 5094 6390 5112 6408
rect 5094 6408 5112 6426
rect 5094 6426 5112 6444
rect 5094 6444 5112 6462
rect 5094 6462 5112 6480
rect 5094 6480 5112 6498
rect 5094 6498 5112 6516
rect 5094 6516 5112 6534
rect 5094 6534 5112 6552
rect 5094 6552 5112 6570
rect 5094 6570 5112 6588
rect 5094 6588 5112 6606
rect 5094 6606 5112 6624
rect 5094 6624 5112 6642
rect 5094 6642 5112 6660
rect 5094 6660 5112 6678
rect 5094 6678 5112 6696
rect 5094 6696 5112 6714
rect 5094 6714 5112 6732
rect 5094 6732 5112 6750
rect 5094 6750 5112 6768
rect 5094 6768 5112 6786
rect 5094 6786 5112 6804
rect 5094 6804 5112 6822
rect 5094 6822 5112 6840
rect 5094 6840 5112 6858
rect 5094 6858 5112 6876
rect 5094 6876 5112 6894
rect 5094 6894 5112 6912
rect 5094 6912 5112 6930
rect 5094 6930 5112 6948
rect 5094 6948 5112 6966
rect 5094 6966 5112 6984
rect 5094 6984 5112 7002
rect 5094 7002 5112 7020
rect 5094 7020 5112 7038
rect 5094 7038 5112 7056
rect 5094 7056 5112 7074
rect 5094 7074 5112 7092
rect 5094 7092 5112 7110
rect 5094 7110 5112 7128
rect 5094 7128 5112 7146
rect 5094 7146 5112 7164
rect 5094 7164 5112 7182
rect 5094 7182 5112 7200
rect 5094 7200 5112 7218
rect 5094 7218 5112 7236
rect 5094 7236 5112 7254
rect 5094 7254 5112 7272
rect 5094 7272 5112 7290
rect 5094 7290 5112 7308
rect 5094 7308 5112 7326
rect 5094 7326 5112 7344
rect 5094 7344 5112 7362
rect 5094 7362 5112 7380
rect 5094 7380 5112 7398
rect 5094 7398 5112 7416
rect 5094 7416 5112 7434
rect 5094 7434 5112 7452
rect 5094 7452 5112 7470
rect 5094 7470 5112 7488
rect 5094 7488 5112 7506
rect 5094 7506 5112 7524
rect 5094 7524 5112 7542
rect 5094 7542 5112 7560
rect 5094 7560 5112 7578
rect 5094 7578 5112 7596
rect 5094 7596 5112 7614
rect 5094 7614 5112 7632
rect 5094 7632 5112 7650
rect 5094 7650 5112 7668
rect 5094 7668 5112 7686
rect 5094 7686 5112 7704
rect 5094 7704 5112 7722
rect 5094 7722 5112 7740
rect 5094 7740 5112 7758
rect 5094 7758 5112 7776
rect 5094 7776 5112 7794
rect 5094 7794 5112 7812
rect 5094 7812 5112 7830
rect 5094 7830 5112 7848
rect 5094 7848 5112 7866
rect 5094 7866 5112 7884
rect 5094 7884 5112 7902
rect 5094 7902 5112 7920
rect 5094 7920 5112 7938
rect 5094 7938 5112 7956
rect 5094 7956 5112 7974
rect 5094 7974 5112 7992
rect 5112 306 5130 324
rect 5112 324 5130 342
rect 5112 342 5130 360
rect 5112 360 5130 378
rect 5112 378 5130 396
rect 5112 396 5130 414
rect 5112 414 5130 432
rect 5112 432 5130 450
rect 5112 450 5130 468
rect 5112 468 5130 486
rect 5112 486 5130 504
rect 5112 504 5130 522
rect 5112 522 5130 540
rect 5112 540 5130 558
rect 5112 558 5130 576
rect 5112 576 5130 594
rect 5112 594 5130 612
rect 5112 612 5130 630
rect 5112 630 5130 648
rect 5112 648 5130 666
rect 5112 666 5130 684
rect 5112 684 5130 702
rect 5112 702 5130 720
rect 5112 720 5130 738
rect 5112 738 5130 756
rect 5112 756 5130 774
rect 5112 900 5130 918
rect 5112 918 5130 936
rect 5112 936 5130 954
rect 5112 954 5130 972
rect 5112 972 5130 990
rect 5112 990 5130 1008
rect 5112 1008 5130 1026
rect 5112 1026 5130 1044
rect 5112 1044 5130 1062
rect 5112 1062 5130 1080
rect 5112 1080 5130 1098
rect 5112 1098 5130 1116
rect 5112 1116 5130 1134
rect 5112 1134 5130 1152
rect 5112 1152 5130 1170
rect 5112 1170 5130 1188
rect 5112 1188 5130 1206
rect 5112 1206 5130 1224
rect 5112 1224 5130 1242
rect 5112 1242 5130 1260
rect 5112 1260 5130 1278
rect 5112 1278 5130 1296
rect 5112 1296 5130 1314
rect 5112 1314 5130 1332
rect 5112 1332 5130 1350
rect 5112 1350 5130 1368
rect 5112 1368 5130 1386
rect 5112 1386 5130 1404
rect 5112 1404 5130 1422
rect 5112 1422 5130 1440
rect 5112 1440 5130 1458
rect 5112 1458 5130 1476
rect 5112 1476 5130 1494
rect 5112 1494 5130 1512
rect 5112 1512 5130 1530
rect 5112 1530 5130 1548
rect 5112 1548 5130 1566
rect 5112 1566 5130 1584
rect 5112 1584 5130 1602
rect 5112 1602 5130 1620
rect 5112 1620 5130 1638
rect 5112 1638 5130 1656
rect 5112 1656 5130 1674
rect 5112 1674 5130 1692
rect 5112 1692 5130 1710
rect 5112 1710 5130 1728
rect 5112 1728 5130 1746
rect 5112 1746 5130 1764
rect 5112 1764 5130 1782
rect 5112 1782 5130 1800
rect 5112 1800 5130 1818
rect 5112 1818 5130 1836
rect 5112 1836 5130 1854
rect 5112 1854 5130 1872
rect 5112 1872 5130 1890
rect 5112 1890 5130 1908
rect 5112 1908 5130 1926
rect 5112 1926 5130 1944
rect 5112 1944 5130 1962
rect 5112 1962 5130 1980
rect 5112 1980 5130 1998
rect 5112 1998 5130 2016
rect 5112 2016 5130 2034
rect 5112 2034 5130 2052
rect 5112 2052 5130 2070
rect 5112 2070 5130 2088
rect 5112 2088 5130 2106
rect 5112 2106 5130 2124
rect 5112 2124 5130 2142
rect 5112 2142 5130 2160
rect 5112 2160 5130 2178
rect 5112 2178 5130 2196
rect 5112 2196 5130 2214
rect 5112 2214 5130 2232
rect 5112 2232 5130 2250
rect 5112 2250 5130 2268
rect 5112 2268 5130 2286
rect 5112 2286 5130 2304
rect 5112 2502 5130 2520
rect 5112 2520 5130 2538
rect 5112 2538 5130 2556
rect 5112 2556 5130 2574
rect 5112 2574 5130 2592
rect 5112 2592 5130 2610
rect 5112 2610 5130 2628
rect 5112 2628 5130 2646
rect 5112 2646 5130 2664
rect 5112 2664 5130 2682
rect 5112 2682 5130 2700
rect 5112 2700 5130 2718
rect 5112 2718 5130 2736
rect 5112 2736 5130 2754
rect 5112 2754 5130 2772
rect 5112 2772 5130 2790
rect 5112 2790 5130 2808
rect 5112 2808 5130 2826
rect 5112 2826 5130 2844
rect 5112 2844 5130 2862
rect 5112 2862 5130 2880
rect 5112 2880 5130 2898
rect 5112 2898 5130 2916
rect 5112 2916 5130 2934
rect 5112 2934 5130 2952
rect 5112 2952 5130 2970
rect 5112 2970 5130 2988
rect 5112 2988 5130 3006
rect 5112 3006 5130 3024
rect 5112 3024 5130 3042
rect 5112 3042 5130 3060
rect 5112 3060 5130 3078
rect 5112 3078 5130 3096
rect 5112 3096 5130 3114
rect 5112 3114 5130 3132
rect 5112 3132 5130 3150
rect 5112 3150 5130 3168
rect 5112 3168 5130 3186
rect 5112 3186 5130 3204
rect 5112 3204 5130 3222
rect 5112 3222 5130 3240
rect 5112 3240 5130 3258
rect 5112 3258 5130 3276
rect 5112 3276 5130 3294
rect 5112 3294 5130 3312
rect 5112 3312 5130 3330
rect 5112 3330 5130 3348
rect 5112 3348 5130 3366
rect 5112 3366 5130 3384
rect 5112 3384 5130 3402
rect 5112 3402 5130 3420
rect 5112 3420 5130 3438
rect 5112 3438 5130 3456
rect 5112 3456 5130 3474
rect 5112 3474 5130 3492
rect 5112 3492 5130 3510
rect 5112 3510 5130 3528
rect 5112 3528 5130 3546
rect 5112 3546 5130 3564
rect 5112 3564 5130 3582
rect 5112 3582 5130 3600
rect 5112 3600 5130 3618
rect 5112 3618 5130 3636
rect 5112 3636 5130 3654
rect 5112 3654 5130 3672
rect 5112 3672 5130 3690
rect 5112 3690 5130 3708
rect 5112 3708 5130 3726
rect 5112 3726 5130 3744
rect 5112 3744 5130 3762
rect 5112 3762 5130 3780
rect 5112 3780 5130 3798
rect 5112 3798 5130 3816
rect 5112 3816 5130 3834
rect 5112 3834 5130 3852
rect 5112 3852 5130 3870
rect 5112 3870 5130 3888
rect 5112 3888 5130 3906
rect 5112 3906 5130 3924
rect 5112 3924 5130 3942
rect 5112 3942 5130 3960
rect 5112 3960 5130 3978
rect 5112 3978 5130 3996
rect 5112 3996 5130 4014
rect 5112 4014 5130 4032
rect 5112 4032 5130 4050
rect 5112 4050 5130 4068
rect 5112 4068 5130 4086
rect 5112 4086 5130 4104
rect 5112 4104 5130 4122
rect 5112 4122 5130 4140
rect 5112 4140 5130 4158
rect 5112 4158 5130 4176
rect 5112 4176 5130 4194
rect 5112 4194 5130 4212
rect 5112 4212 5130 4230
rect 5112 4230 5130 4248
rect 5112 4248 5130 4266
rect 5112 4266 5130 4284
rect 5112 4284 5130 4302
rect 5112 4302 5130 4320
rect 5112 4320 5130 4338
rect 5112 4338 5130 4356
rect 5112 4356 5130 4374
rect 5112 4374 5130 4392
rect 5112 4392 5130 4410
rect 5112 4410 5130 4428
rect 5112 4428 5130 4446
rect 5112 4446 5130 4464
rect 5112 4464 5130 4482
rect 5112 4482 5130 4500
rect 5112 4716 5130 4734
rect 5112 4734 5130 4752
rect 5112 4752 5130 4770
rect 5112 4770 5130 4788
rect 5112 4788 5130 4806
rect 5112 4806 5130 4824
rect 5112 4824 5130 4842
rect 5112 4842 5130 4860
rect 5112 4860 5130 4878
rect 5112 4878 5130 4896
rect 5112 4896 5130 4914
rect 5112 4914 5130 4932
rect 5112 4932 5130 4950
rect 5112 4950 5130 4968
rect 5112 4968 5130 4986
rect 5112 4986 5130 5004
rect 5112 5004 5130 5022
rect 5112 5022 5130 5040
rect 5112 5040 5130 5058
rect 5112 5058 5130 5076
rect 5112 5076 5130 5094
rect 5112 5094 5130 5112
rect 5112 5112 5130 5130
rect 5112 5130 5130 5148
rect 5112 5148 5130 5166
rect 5112 5166 5130 5184
rect 5112 5184 5130 5202
rect 5112 5202 5130 5220
rect 5112 5220 5130 5238
rect 5112 5238 5130 5256
rect 5112 5256 5130 5274
rect 5112 5274 5130 5292
rect 5112 5292 5130 5310
rect 5112 5310 5130 5328
rect 5112 5328 5130 5346
rect 5112 5346 5130 5364
rect 5112 5364 5130 5382
rect 5112 5382 5130 5400
rect 5112 5400 5130 5418
rect 5112 5418 5130 5436
rect 5112 5436 5130 5454
rect 5112 5454 5130 5472
rect 5112 5472 5130 5490
rect 5112 5490 5130 5508
rect 5112 5508 5130 5526
rect 5112 5526 5130 5544
rect 5112 5544 5130 5562
rect 5112 5562 5130 5580
rect 5112 5580 5130 5598
rect 5112 5598 5130 5616
rect 5112 5616 5130 5634
rect 5112 5634 5130 5652
rect 5112 5652 5130 5670
rect 5112 5670 5130 5688
rect 5112 5688 5130 5706
rect 5112 5706 5130 5724
rect 5112 5724 5130 5742
rect 5112 5742 5130 5760
rect 5112 5760 5130 5778
rect 5112 5778 5130 5796
rect 5112 5796 5130 5814
rect 5112 5814 5130 5832
rect 5112 5832 5130 5850
rect 5112 5850 5130 5868
rect 5112 5868 5130 5886
rect 5112 5886 5130 5904
rect 5112 5904 5130 5922
rect 5112 5922 5130 5940
rect 5112 5940 5130 5958
rect 5112 5958 5130 5976
rect 5112 5976 5130 5994
rect 5112 5994 5130 6012
rect 5112 6012 5130 6030
rect 5112 6030 5130 6048
rect 5112 6048 5130 6066
rect 5112 6066 5130 6084
rect 5112 6084 5130 6102
rect 5112 6102 5130 6120
rect 5112 6120 5130 6138
rect 5112 6138 5130 6156
rect 5112 6156 5130 6174
rect 5112 6174 5130 6192
rect 5112 6192 5130 6210
rect 5112 6210 5130 6228
rect 5112 6228 5130 6246
rect 5112 6246 5130 6264
rect 5112 6264 5130 6282
rect 5112 6282 5130 6300
rect 5112 6300 5130 6318
rect 5112 6318 5130 6336
rect 5112 6336 5130 6354
rect 5112 6354 5130 6372
rect 5112 6372 5130 6390
rect 5112 6390 5130 6408
rect 5112 6408 5130 6426
rect 5112 6426 5130 6444
rect 5112 6444 5130 6462
rect 5112 6462 5130 6480
rect 5112 6480 5130 6498
rect 5112 6498 5130 6516
rect 5112 6516 5130 6534
rect 5112 6534 5130 6552
rect 5112 6552 5130 6570
rect 5112 6570 5130 6588
rect 5112 6588 5130 6606
rect 5112 6606 5130 6624
rect 5112 6624 5130 6642
rect 5112 6642 5130 6660
rect 5112 6660 5130 6678
rect 5112 6678 5130 6696
rect 5112 6696 5130 6714
rect 5112 6714 5130 6732
rect 5112 6732 5130 6750
rect 5112 6750 5130 6768
rect 5112 6768 5130 6786
rect 5112 6786 5130 6804
rect 5112 6804 5130 6822
rect 5112 6822 5130 6840
rect 5112 6840 5130 6858
rect 5112 6858 5130 6876
rect 5112 6876 5130 6894
rect 5112 6894 5130 6912
rect 5112 6912 5130 6930
rect 5112 6930 5130 6948
rect 5112 6948 5130 6966
rect 5112 6966 5130 6984
rect 5112 6984 5130 7002
rect 5112 7002 5130 7020
rect 5112 7020 5130 7038
rect 5112 7038 5130 7056
rect 5112 7056 5130 7074
rect 5112 7074 5130 7092
rect 5112 7092 5130 7110
rect 5112 7110 5130 7128
rect 5112 7128 5130 7146
rect 5112 7146 5130 7164
rect 5112 7164 5130 7182
rect 5112 7182 5130 7200
rect 5112 7200 5130 7218
rect 5112 7218 5130 7236
rect 5112 7236 5130 7254
rect 5112 7254 5130 7272
rect 5112 7272 5130 7290
rect 5112 7290 5130 7308
rect 5112 7308 5130 7326
rect 5112 7326 5130 7344
rect 5112 7344 5130 7362
rect 5112 7362 5130 7380
rect 5112 7380 5130 7398
rect 5112 7398 5130 7416
rect 5112 7416 5130 7434
rect 5112 7434 5130 7452
rect 5112 7452 5130 7470
rect 5112 7470 5130 7488
rect 5112 7488 5130 7506
rect 5112 7506 5130 7524
rect 5112 7524 5130 7542
rect 5112 7542 5130 7560
rect 5112 7560 5130 7578
rect 5112 7578 5130 7596
rect 5112 7596 5130 7614
rect 5112 7614 5130 7632
rect 5112 7632 5130 7650
rect 5112 7650 5130 7668
rect 5112 7668 5130 7686
rect 5112 7686 5130 7704
rect 5112 7704 5130 7722
rect 5112 7722 5130 7740
rect 5112 7740 5130 7758
rect 5112 7758 5130 7776
rect 5112 7776 5130 7794
rect 5112 7794 5130 7812
rect 5112 7812 5130 7830
rect 5112 7830 5130 7848
rect 5112 7848 5130 7866
rect 5112 7866 5130 7884
rect 5112 7884 5130 7902
rect 5112 7902 5130 7920
rect 5112 7920 5130 7938
rect 5112 7938 5130 7956
rect 5112 7956 5130 7974
rect 5112 7974 5130 7992
rect 5112 7992 5130 8010
rect 5130 324 5148 342
rect 5130 342 5148 360
rect 5130 360 5148 378
rect 5130 378 5148 396
rect 5130 396 5148 414
rect 5130 414 5148 432
rect 5130 432 5148 450
rect 5130 450 5148 468
rect 5130 468 5148 486
rect 5130 486 5148 504
rect 5130 504 5148 522
rect 5130 522 5148 540
rect 5130 540 5148 558
rect 5130 558 5148 576
rect 5130 576 5148 594
rect 5130 594 5148 612
rect 5130 612 5148 630
rect 5130 630 5148 648
rect 5130 648 5148 666
rect 5130 666 5148 684
rect 5130 684 5148 702
rect 5130 702 5148 720
rect 5130 720 5148 738
rect 5130 738 5148 756
rect 5130 756 5148 774
rect 5130 918 5148 936
rect 5130 936 5148 954
rect 5130 954 5148 972
rect 5130 972 5148 990
rect 5130 990 5148 1008
rect 5130 1008 5148 1026
rect 5130 1026 5148 1044
rect 5130 1044 5148 1062
rect 5130 1062 5148 1080
rect 5130 1080 5148 1098
rect 5130 1098 5148 1116
rect 5130 1116 5148 1134
rect 5130 1134 5148 1152
rect 5130 1152 5148 1170
rect 5130 1170 5148 1188
rect 5130 1188 5148 1206
rect 5130 1206 5148 1224
rect 5130 1224 5148 1242
rect 5130 1242 5148 1260
rect 5130 1260 5148 1278
rect 5130 1278 5148 1296
rect 5130 1296 5148 1314
rect 5130 1314 5148 1332
rect 5130 1332 5148 1350
rect 5130 1350 5148 1368
rect 5130 1368 5148 1386
rect 5130 1386 5148 1404
rect 5130 1404 5148 1422
rect 5130 1422 5148 1440
rect 5130 1440 5148 1458
rect 5130 1458 5148 1476
rect 5130 1476 5148 1494
rect 5130 1494 5148 1512
rect 5130 1512 5148 1530
rect 5130 1530 5148 1548
rect 5130 1548 5148 1566
rect 5130 1566 5148 1584
rect 5130 1584 5148 1602
rect 5130 1602 5148 1620
rect 5130 1620 5148 1638
rect 5130 1638 5148 1656
rect 5130 1656 5148 1674
rect 5130 1674 5148 1692
rect 5130 1692 5148 1710
rect 5130 1710 5148 1728
rect 5130 1728 5148 1746
rect 5130 1746 5148 1764
rect 5130 1764 5148 1782
rect 5130 1782 5148 1800
rect 5130 1800 5148 1818
rect 5130 1818 5148 1836
rect 5130 1836 5148 1854
rect 5130 1854 5148 1872
rect 5130 1872 5148 1890
rect 5130 1890 5148 1908
rect 5130 1908 5148 1926
rect 5130 1926 5148 1944
rect 5130 1944 5148 1962
rect 5130 1962 5148 1980
rect 5130 1980 5148 1998
rect 5130 1998 5148 2016
rect 5130 2016 5148 2034
rect 5130 2034 5148 2052
rect 5130 2052 5148 2070
rect 5130 2070 5148 2088
rect 5130 2088 5148 2106
rect 5130 2106 5148 2124
rect 5130 2124 5148 2142
rect 5130 2142 5148 2160
rect 5130 2160 5148 2178
rect 5130 2178 5148 2196
rect 5130 2196 5148 2214
rect 5130 2214 5148 2232
rect 5130 2232 5148 2250
rect 5130 2250 5148 2268
rect 5130 2268 5148 2286
rect 5130 2286 5148 2304
rect 5130 2520 5148 2538
rect 5130 2538 5148 2556
rect 5130 2556 5148 2574
rect 5130 2574 5148 2592
rect 5130 2592 5148 2610
rect 5130 2610 5148 2628
rect 5130 2628 5148 2646
rect 5130 2646 5148 2664
rect 5130 2664 5148 2682
rect 5130 2682 5148 2700
rect 5130 2700 5148 2718
rect 5130 2718 5148 2736
rect 5130 2736 5148 2754
rect 5130 2754 5148 2772
rect 5130 2772 5148 2790
rect 5130 2790 5148 2808
rect 5130 2808 5148 2826
rect 5130 2826 5148 2844
rect 5130 2844 5148 2862
rect 5130 2862 5148 2880
rect 5130 2880 5148 2898
rect 5130 2898 5148 2916
rect 5130 2916 5148 2934
rect 5130 2934 5148 2952
rect 5130 2952 5148 2970
rect 5130 2970 5148 2988
rect 5130 2988 5148 3006
rect 5130 3006 5148 3024
rect 5130 3024 5148 3042
rect 5130 3042 5148 3060
rect 5130 3060 5148 3078
rect 5130 3078 5148 3096
rect 5130 3096 5148 3114
rect 5130 3114 5148 3132
rect 5130 3132 5148 3150
rect 5130 3150 5148 3168
rect 5130 3168 5148 3186
rect 5130 3186 5148 3204
rect 5130 3204 5148 3222
rect 5130 3222 5148 3240
rect 5130 3240 5148 3258
rect 5130 3258 5148 3276
rect 5130 3276 5148 3294
rect 5130 3294 5148 3312
rect 5130 3312 5148 3330
rect 5130 3330 5148 3348
rect 5130 3348 5148 3366
rect 5130 3366 5148 3384
rect 5130 3384 5148 3402
rect 5130 3402 5148 3420
rect 5130 3420 5148 3438
rect 5130 3438 5148 3456
rect 5130 3456 5148 3474
rect 5130 3474 5148 3492
rect 5130 3492 5148 3510
rect 5130 3510 5148 3528
rect 5130 3528 5148 3546
rect 5130 3546 5148 3564
rect 5130 3564 5148 3582
rect 5130 3582 5148 3600
rect 5130 3600 5148 3618
rect 5130 3618 5148 3636
rect 5130 3636 5148 3654
rect 5130 3654 5148 3672
rect 5130 3672 5148 3690
rect 5130 3690 5148 3708
rect 5130 3708 5148 3726
rect 5130 3726 5148 3744
rect 5130 3744 5148 3762
rect 5130 3762 5148 3780
rect 5130 3780 5148 3798
rect 5130 3798 5148 3816
rect 5130 3816 5148 3834
rect 5130 3834 5148 3852
rect 5130 3852 5148 3870
rect 5130 3870 5148 3888
rect 5130 3888 5148 3906
rect 5130 3906 5148 3924
rect 5130 3924 5148 3942
rect 5130 3942 5148 3960
rect 5130 3960 5148 3978
rect 5130 3978 5148 3996
rect 5130 3996 5148 4014
rect 5130 4014 5148 4032
rect 5130 4032 5148 4050
rect 5130 4050 5148 4068
rect 5130 4068 5148 4086
rect 5130 4086 5148 4104
rect 5130 4104 5148 4122
rect 5130 4122 5148 4140
rect 5130 4140 5148 4158
rect 5130 4158 5148 4176
rect 5130 4176 5148 4194
rect 5130 4194 5148 4212
rect 5130 4212 5148 4230
rect 5130 4230 5148 4248
rect 5130 4248 5148 4266
rect 5130 4266 5148 4284
rect 5130 4284 5148 4302
rect 5130 4302 5148 4320
rect 5130 4320 5148 4338
rect 5130 4338 5148 4356
rect 5130 4356 5148 4374
rect 5130 4374 5148 4392
rect 5130 4392 5148 4410
rect 5130 4410 5148 4428
rect 5130 4428 5148 4446
rect 5130 4446 5148 4464
rect 5130 4464 5148 4482
rect 5130 4482 5148 4500
rect 5130 4500 5148 4518
rect 5130 4734 5148 4752
rect 5130 4752 5148 4770
rect 5130 4770 5148 4788
rect 5130 4788 5148 4806
rect 5130 4806 5148 4824
rect 5130 4824 5148 4842
rect 5130 4842 5148 4860
rect 5130 4860 5148 4878
rect 5130 4878 5148 4896
rect 5130 4896 5148 4914
rect 5130 4914 5148 4932
rect 5130 4932 5148 4950
rect 5130 4950 5148 4968
rect 5130 4968 5148 4986
rect 5130 4986 5148 5004
rect 5130 5004 5148 5022
rect 5130 5022 5148 5040
rect 5130 5040 5148 5058
rect 5130 5058 5148 5076
rect 5130 5076 5148 5094
rect 5130 5094 5148 5112
rect 5130 5112 5148 5130
rect 5130 5130 5148 5148
rect 5130 5148 5148 5166
rect 5130 5166 5148 5184
rect 5130 5184 5148 5202
rect 5130 5202 5148 5220
rect 5130 5220 5148 5238
rect 5130 5238 5148 5256
rect 5130 5256 5148 5274
rect 5130 5274 5148 5292
rect 5130 5292 5148 5310
rect 5130 5310 5148 5328
rect 5130 5328 5148 5346
rect 5130 5346 5148 5364
rect 5130 5364 5148 5382
rect 5130 5382 5148 5400
rect 5130 5400 5148 5418
rect 5130 5418 5148 5436
rect 5130 5436 5148 5454
rect 5130 5454 5148 5472
rect 5130 5472 5148 5490
rect 5130 5490 5148 5508
rect 5130 5508 5148 5526
rect 5130 5526 5148 5544
rect 5130 5544 5148 5562
rect 5130 5562 5148 5580
rect 5130 5580 5148 5598
rect 5130 5598 5148 5616
rect 5130 5616 5148 5634
rect 5130 5634 5148 5652
rect 5130 5652 5148 5670
rect 5130 5670 5148 5688
rect 5130 5688 5148 5706
rect 5130 5706 5148 5724
rect 5130 5724 5148 5742
rect 5130 5742 5148 5760
rect 5130 5760 5148 5778
rect 5130 5778 5148 5796
rect 5130 5796 5148 5814
rect 5130 5814 5148 5832
rect 5130 5832 5148 5850
rect 5130 5850 5148 5868
rect 5130 5868 5148 5886
rect 5130 5886 5148 5904
rect 5130 5904 5148 5922
rect 5130 5922 5148 5940
rect 5130 5940 5148 5958
rect 5130 5958 5148 5976
rect 5130 5976 5148 5994
rect 5130 5994 5148 6012
rect 5130 6012 5148 6030
rect 5130 6030 5148 6048
rect 5130 6048 5148 6066
rect 5130 6066 5148 6084
rect 5130 6084 5148 6102
rect 5130 6102 5148 6120
rect 5130 6120 5148 6138
rect 5130 6138 5148 6156
rect 5130 6156 5148 6174
rect 5130 6174 5148 6192
rect 5130 6192 5148 6210
rect 5130 6210 5148 6228
rect 5130 6228 5148 6246
rect 5130 6246 5148 6264
rect 5130 6264 5148 6282
rect 5130 6282 5148 6300
rect 5130 6300 5148 6318
rect 5130 6318 5148 6336
rect 5130 6336 5148 6354
rect 5130 6354 5148 6372
rect 5130 6372 5148 6390
rect 5130 6390 5148 6408
rect 5130 6408 5148 6426
rect 5130 6426 5148 6444
rect 5130 6444 5148 6462
rect 5130 6462 5148 6480
rect 5130 6480 5148 6498
rect 5130 6498 5148 6516
rect 5130 6516 5148 6534
rect 5130 6534 5148 6552
rect 5130 6552 5148 6570
rect 5130 6570 5148 6588
rect 5130 6588 5148 6606
rect 5130 6606 5148 6624
rect 5130 6624 5148 6642
rect 5130 6642 5148 6660
rect 5130 6660 5148 6678
rect 5130 6678 5148 6696
rect 5130 6696 5148 6714
rect 5130 6714 5148 6732
rect 5130 6732 5148 6750
rect 5130 6750 5148 6768
rect 5130 6768 5148 6786
rect 5130 6786 5148 6804
rect 5130 6804 5148 6822
rect 5130 6822 5148 6840
rect 5130 6840 5148 6858
rect 5130 6858 5148 6876
rect 5130 6876 5148 6894
rect 5130 6894 5148 6912
rect 5130 6912 5148 6930
rect 5130 6930 5148 6948
rect 5130 6948 5148 6966
rect 5130 6966 5148 6984
rect 5130 6984 5148 7002
rect 5130 7002 5148 7020
rect 5130 7020 5148 7038
rect 5130 7038 5148 7056
rect 5130 7056 5148 7074
rect 5130 7074 5148 7092
rect 5130 7092 5148 7110
rect 5130 7110 5148 7128
rect 5130 7128 5148 7146
rect 5130 7146 5148 7164
rect 5130 7164 5148 7182
rect 5130 7182 5148 7200
rect 5130 7200 5148 7218
rect 5130 7218 5148 7236
rect 5130 7236 5148 7254
rect 5130 7254 5148 7272
rect 5130 7272 5148 7290
rect 5130 7290 5148 7308
rect 5130 7308 5148 7326
rect 5130 7326 5148 7344
rect 5130 7344 5148 7362
rect 5130 7362 5148 7380
rect 5130 7380 5148 7398
rect 5130 7398 5148 7416
rect 5130 7416 5148 7434
rect 5130 7434 5148 7452
rect 5130 7452 5148 7470
rect 5130 7470 5148 7488
rect 5130 7488 5148 7506
rect 5130 7506 5148 7524
rect 5130 7524 5148 7542
rect 5130 7542 5148 7560
rect 5130 7560 5148 7578
rect 5130 7578 5148 7596
rect 5130 7596 5148 7614
rect 5130 7614 5148 7632
rect 5130 7632 5148 7650
rect 5130 7650 5148 7668
rect 5130 7668 5148 7686
rect 5130 7686 5148 7704
rect 5130 7704 5148 7722
rect 5130 7722 5148 7740
rect 5130 7740 5148 7758
rect 5130 7758 5148 7776
rect 5130 7776 5148 7794
rect 5130 7794 5148 7812
rect 5130 7812 5148 7830
rect 5130 7830 5148 7848
rect 5130 7848 5148 7866
rect 5130 7866 5148 7884
rect 5130 7884 5148 7902
rect 5130 7902 5148 7920
rect 5130 7920 5148 7938
rect 5130 7938 5148 7956
rect 5130 7956 5148 7974
rect 5130 7974 5148 7992
rect 5130 7992 5148 8010
rect 5130 8010 5148 8028
rect 5130 8028 5148 8046
rect 5148 324 5166 342
rect 5148 342 5166 360
rect 5148 360 5166 378
rect 5148 378 5166 396
rect 5148 396 5166 414
rect 5148 414 5166 432
rect 5148 432 5166 450
rect 5148 450 5166 468
rect 5148 468 5166 486
rect 5148 486 5166 504
rect 5148 504 5166 522
rect 5148 522 5166 540
rect 5148 540 5166 558
rect 5148 558 5166 576
rect 5148 576 5166 594
rect 5148 594 5166 612
rect 5148 612 5166 630
rect 5148 630 5166 648
rect 5148 648 5166 666
rect 5148 666 5166 684
rect 5148 684 5166 702
rect 5148 702 5166 720
rect 5148 720 5166 738
rect 5148 738 5166 756
rect 5148 756 5166 774
rect 5148 774 5166 792
rect 5148 918 5166 936
rect 5148 936 5166 954
rect 5148 954 5166 972
rect 5148 972 5166 990
rect 5148 990 5166 1008
rect 5148 1008 5166 1026
rect 5148 1026 5166 1044
rect 5148 1044 5166 1062
rect 5148 1062 5166 1080
rect 5148 1080 5166 1098
rect 5148 1098 5166 1116
rect 5148 1116 5166 1134
rect 5148 1134 5166 1152
rect 5148 1152 5166 1170
rect 5148 1170 5166 1188
rect 5148 1188 5166 1206
rect 5148 1206 5166 1224
rect 5148 1224 5166 1242
rect 5148 1242 5166 1260
rect 5148 1260 5166 1278
rect 5148 1278 5166 1296
rect 5148 1296 5166 1314
rect 5148 1314 5166 1332
rect 5148 1332 5166 1350
rect 5148 1350 5166 1368
rect 5148 1368 5166 1386
rect 5148 1386 5166 1404
rect 5148 1404 5166 1422
rect 5148 1422 5166 1440
rect 5148 1440 5166 1458
rect 5148 1458 5166 1476
rect 5148 1476 5166 1494
rect 5148 1494 5166 1512
rect 5148 1512 5166 1530
rect 5148 1530 5166 1548
rect 5148 1548 5166 1566
rect 5148 1566 5166 1584
rect 5148 1584 5166 1602
rect 5148 1602 5166 1620
rect 5148 1620 5166 1638
rect 5148 1638 5166 1656
rect 5148 1656 5166 1674
rect 5148 1674 5166 1692
rect 5148 1692 5166 1710
rect 5148 1710 5166 1728
rect 5148 1728 5166 1746
rect 5148 1746 5166 1764
rect 5148 1764 5166 1782
rect 5148 1782 5166 1800
rect 5148 1800 5166 1818
rect 5148 1818 5166 1836
rect 5148 1836 5166 1854
rect 5148 1854 5166 1872
rect 5148 1872 5166 1890
rect 5148 1890 5166 1908
rect 5148 1908 5166 1926
rect 5148 1926 5166 1944
rect 5148 1944 5166 1962
rect 5148 1962 5166 1980
rect 5148 1980 5166 1998
rect 5148 1998 5166 2016
rect 5148 2016 5166 2034
rect 5148 2034 5166 2052
rect 5148 2052 5166 2070
rect 5148 2070 5166 2088
rect 5148 2088 5166 2106
rect 5148 2106 5166 2124
rect 5148 2124 5166 2142
rect 5148 2142 5166 2160
rect 5148 2160 5166 2178
rect 5148 2178 5166 2196
rect 5148 2196 5166 2214
rect 5148 2214 5166 2232
rect 5148 2232 5166 2250
rect 5148 2250 5166 2268
rect 5148 2268 5166 2286
rect 5148 2286 5166 2304
rect 5148 2304 5166 2322
rect 5148 2538 5166 2556
rect 5148 2556 5166 2574
rect 5148 2574 5166 2592
rect 5148 2592 5166 2610
rect 5148 2610 5166 2628
rect 5148 2628 5166 2646
rect 5148 2646 5166 2664
rect 5148 2664 5166 2682
rect 5148 2682 5166 2700
rect 5148 2700 5166 2718
rect 5148 2718 5166 2736
rect 5148 2736 5166 2754
rect 5148 2754 5166 2772
rect 5148 2772 5166 2790
rect 5148 2790 5166 2808
rect 5148 2808 5166 2826
rect 5148 2826 5166 2844
rect 5148 2844 5166 2862
rect 5148 2862 5166 2880
rect 5148 2880 5166 2898
rect 5148 2898 5166 2916
rect 5148 2916 5166 2934
rect 5148 2934 5166 2952
rect 5148 2952 5166 2970
rect 5148 2970 5166 2988
rect 5148 2988 5166 3006
rect 5148 3006 5166 3024
rect 5148 3024 5166 3042
rect 5148 3042 5166 3060
rect 5148 3060 5166 3078
rect 5148 3078 5166 3096
rect 5148 3096 5166 3114
rect 5148 3114 5166 3132
rect 5148 3132 5166 3150
rect 5148 3150 5166 3168
rect 5148 3168 5166 3186
rect 5148 3186 5166 3204
rect 5148 3204 5166 3222
rect 5148 3222 5166 3240
rect 5148 3240 5166 3258
rect 5148 3258 5166 3276
rect 5148 3276 5166 3294
rect 5148 3294 5166 3312
rect 5148 3312 5166 3330
rect 5148 3330 5166 3348
rect 5148 3348 5166 3366
rect 5148 3366 5166 3384
rect 5148 3384 5166 3402
rect 5148 3402 5166 3420
rect 5148 3420 5166 3438
rect 5148 3438 5166 3456
rect 5148 3456 5166 3474
rect 5148 3474 5166 3492
rect 5148 3492 5166 3510
rect 5148 3510 5166 3528
rect 5148 3528 5166 3546
rect 5148 3546 5166 3564
rect 5148 3564 5166 3582
rect 5148 3582 5166 3600
rect 5148 3600 5166 3618
rect 5148 3618 5166 3636
rect 5148 3636 5166 3654
rect 5148 3654 5166 3672
rect 5148 3672 5166 3690
rect 5148 3690 5166 3708
rect 5148 3708 5166 3726
rect 5148 3726 5166 3744
rect 5148 3744 5166 3762
rect 5148 3762 5166 3780
rect 5148 3780 5166 3798
rect 5148 3798 5166 3816
rect 5148 3816 5166 3834
rect 5148 3834 5166 3852
rect 5148 3852 5166 3870
rect 5148 3870 5166 3888
rect 5148 3888 5166 3906
rect 5148 3906 5166 3924
rect 5148 3924 5166 3942
rect 5148 3942 5166 3960
rect 5148 3960 5166 3978
rect 5148 3978 5166 3996
rect 5148 3996 5166 4014
rect 5148 4014 5166 4032
rect 5148 4032 5166 4050
rect 5148 4050 5166 4068
rect 5148 4068 5166 4086
rect 5148 4086 5166 4104
rect 5148 4104 5166 4122
rect 5148 4122 5166 4140
rect 5148 4140 5166 4158
rect 5148 4158 5166 4176
rect 5148 4176 5166 4194
rect 5148 4194 5166 4212
rect 5148 4212 5166 4230
rect 5148 4230 5166 4248
rect 5148 4248 5166 4266
rect 5148 4266 5166 4284
rect 5148 4284 5166 4302
rect 5148 4302 5166 4320
rect 5148 4320 5166 4338
rect 5148 4338 5166 4356
rect 5148 4356 5166 4374
rect 5148 4374 5166 4392
rect 5148 4392 5166 4410
rect 5148 4410 5166 4428
rect 5148 4428 5166 4446
rect 5148 4446 5166 4464
rect 5148 4464 5166 4482
rect 5148 4482 5166 4500
rect 5148 4500 5166 4518
rect 5148 4518 5166 4536
rect 5148 4752 5166 4770
rect 5148 4770 5166 4788
rect 5148 4788 5166 4806
rect 5148 4806 5166 4824
rect 5148 4824 5166 4842
rect 5148 4842 5166 4860
rect 5148 4860 5166 4878
rect 5148 4878 5166 4896
rect 5148 4896 5166 4914
rect 5148 4914 5166 4932
rect 5148 4932 5166 4950
rect 5148 4950 5166 4968
rect 5148 4968 5166 4986
rect 5148 4986 5166 5004
rect 5148 5004 5166 5022
rect 5148 5022 5166 5040
rect 5148 5040 5166 5058
rect 5148 5058 5166 5076
rect 5148 5076 5166 5094
rect 5148 5094 5166 5112
rect 5148 5112 5166 5130
rect 5148 5130 5166 5148
rect 5148 5148 5166 5166
rect 5148 5166 5166 5184
rect 5148 5184 5166 5202
rect 5148 5202 5166 5220
rect 5148 5220 5166 5238
rect 5148 5238 5166 5256
rect 5148 5256 5166 5274
rect 5148 5274 5166 5292
rect 5148 5292 5166 5310
rect 5148 5310 5166 5328
rect 5148 5328 5166 5346
rect 5148 5346 5166 5364
rect 5148 5364 5166 5382
rect 5148 5382 5166 5400
rect 5148 5400 5166 5418
rect 5148 5418 5166 5436
rect 5148 5436 5166 5454
rect 5148 5454 5166 5472
rect 5148 5472 5166 5490
rect 5148 5490 5166 5508
rect 5148 5508 5166 5526
rect 5148 5526 5166 5544
rect 5148 5544 5166 5562
rect 5148 5562 5166 5580
rect 5148 5580 5166 5598
rect 5148 5598 5166 5616
rect 5148 5616 5166 5634
rect 5148 5634 5166 5652
rect 5148 5652 5166 5670
rect 5148 5670 5166 5688
rect 5148 5688 5166 5706
rect 5148 5706 5166 5724
rect 5148 5724 5166 5742
rect 5148 5742 5166 5760
rect 5148 5760 5166 5778
rect 5148 5778 5166 5796
rect 5148 5796 5166 5814
rect 5148 5814 5166 5832
rect 5148 5832 5166 5850
rect 5148 5850 5166 5868
rect 5148 5868 5166 5886
rect 5148 5886 5166 5904
rect 5148 5904 5166 5922
rect 5148 5922 5166 5940
rect 5148 5940 5166 5958
rect 5148 5958 5166 5976
rect 5148 5976 5166 5994
rect 5148 5994 5166 6012
rect 5148 6012 5166 6030
rect 5148 6030 5166 6048
rect 5148 6048 5166 6066
rect 5148 6066 5166 6084
rect 5148 6084 5166 6102
rect 5148 6102 5166 6120
rect 5148 6120 5166 6138
rect 5148 6138 5166 6156
rect 5148 6156 5166 6174
rect 5148 6174 5166 6192
rect 5148 6192 5166 6210
rect 5148 6210 5166 6228
rect 5148 6228 5166 6246
rect 5148 6246 5166 6264
rect 5148 6264 5166 6282
rect 5148 6282 5166 6300
rect 5148 6300 5166 6318
rect 5148 6318 5166 6336
rect 5148 6336 5166 6354
rect 5148 6354 5166 6372
rect 5148 6372 5166 6390
rect 5148 6390 5166 6408
rect 5148 6408 5166 6426
rect 5148 6426 5166 6444
rect 5148 6444 5166 6462
rect 5148 6462 5166 6480
rect 5148 6480 5166 6498
rect 5148 6498 5166 6516
rect 5148 6516 5166 6534
rect 5148 6534 5166 6552
rect 5148 6552 5166 6570
rect 5148 6570 5166 6588
rect 5148 6588 5166 6606
rect 5148 6606 5166 6624
rect 5148 6624 5166 6642
rect 5148 6642 5166 6660
rect 5148 6660 5166 6678
rect 5148 6678 5166 6696
rect 5148 6696 5166 6714
rect 5148 6714 5166 6732
rect 5148 6732 5166 6750
rect 5148 6750 5166 6768
rect 5148 6768 5166 6786
rect 5148 6786 5166 6804
rect 5148 6804 5166 6822
rect 5148 6822 5166 6840
rect 5148 6840 5166 6858
rect 5148 6858 5166 6876
rect 5148 6876 5166 6894
rect 5148 6894 5166 6912
rect 5148 6912 5166 6930
rect 5148 6930 5166 6948
rect 5148 6948 5166 6966
rect 5148 6966 5166 6984
rect 5148 6984 5166 7002
rect 5148 7002 5166 7020
rect 5148 7020 5166 7038
rect 5148 7038 5166 7056
rect 5148 7056 5166 7074
rect 5148 7074 5166 7092
rect 5148 7092 5166 7110
rect 5148 7110 5166 7128
rect 5148 7128 5166 7146
rect 5148 7146 5166 7164
rect 5148 7164 5166 7182
rect 5148 7182 5166 7200
rect 5148 7200 5166 7218
rect 5148 7218 5166 7236
rect 5148 7236 5166 7254
rect 5148 7254 5166 7272
rect 5148 7272 5166 7290
rect 5148 7290 5166 7308
rect 5148 7308 5166 7326
rect 5148 7326 5166 7344
rect 5148 7344 5166 7362
rect 5148 7362 5166 7380
rect 5148 7380 5166 7398
rect 5148 7398 5166 7416
rect 5148 7416 5166 7434
rect 5148 7434 5166 7452
rect 5148 7452 5166 7470
rect 5148 7470 5166 7488
rect 5148 7488 5166 7506
rect 5148 7506 5166 7524
rect 5148 7524 5166 7542
rect 5148 7542 5166 7560
rect 5148 7560 5166 7578
rect 5148 7578 5166 7596
rect 5148 7596 5166 7614
rect 5148 7614 5166 7632
rect 5148 7632 5166 7650
rect 5148 7650 5166 7668
rect 5148 7668 5166 7686
rect 5148 7686 5166 7704
rect 5148 7704 5166 7722
rect 5148 7722 5166 7740
rect 5148 7740 5166 7758
rect 5148 7758 5166 7776
rect 5148 7776 5166 7794
rect 5148 7794 5166 7812
rect 5148 7812 5166 7830
rect 5148 7830 5166 7848
rect 5148 7848 5166 7866
rect 5148 7866 5166 7884
rect 5148 7884 5166 7902
rect 5148 7902 5166 7920
rect 5148 7920 5166 7938
rect 5148 7938 5166 7956
rect 5148 7956 5166 7974
rect 5148 7974 5166 7992
rect 5148 7992 5166 8010
rect 5148 8010 5166 8028
rect 5148 8028 5166 8046
rect 5148 8046 5166 8064
rect 5166 342 5184 360
rect 5166 360 5184 378
rect 5166 378 5184 396
rect 5166 396 5184 414
rect 5166 414 5184 432
rect 5166 432 5184 450
rect 5166 450 5184 468
rect 5166 468 5184 486
rect 5166 486 5184 504
rect 5166 504 5184 522
rect 5166 522 5184 540
rect 5166 540 5184 558
rect 5166 558 5184 576
rect 5166 576 5184 594
rect 5166 594 5184 612
rect 5166 612 5184 630
rect 5166 630 5184 648
rect 5166 648 5184 666
rect 5166 666 5184 684
rect 5166 684 5184 702
rect 5166 702 5184 720
rect 5166 720 5184 738
rect 5166 738 5184 756
rect 5166 756 5184 774
rect 5166 774 5184 792
rect 5166 918 5184 936
rect 5166 936 5184 954
rect 5166 954 5184 972
rect 5166 972 5184 990
rect 5166 990 5184 1008
rect 5166 1008 5184 1026
rect 5166 1026 5184 1044
rect 5166 1044 5184 1062
rect 5166 1062 5184 1080
rect 5166 1080 5184 1098
rect 5166 1098 5184 1116
rect 5166 1116 5184 1134
rect 5166 1134 5184 1152
rect 5166 1152 5184 1170
rect 5166 1170 5184 1188
rect 5166 1188 5184 1206
rect 5166 1206 5184 1224
rect 5166 1224 5184 1242
rect 5166 1242 5184 1260
rect 5166 1260 5184 1278
rect 5166 1278 5184 1296
rect 5166 1296 5184 1314
rect 5166 1314 5184 1332
rect 5166 1332 5184 1350
rect 5166 1350 5184 1368
rect 5166 1368 5184 1386
rect 5166 1386 5184 1404
rect 5166 1404 5184 1422
rect 5166 1422 5184 1440
rect 5166 1440 5184 1458
rect 5166 1458 5184 1476
rect 5166 1476 5184 1494
rect 5166 1494 5184 1512
rect 5166 1512 5184 1530
rect 5166 1530 5184 1548
rect 5166 1548 5184 1566
rect 5166 1566 5184 1584
rect 5166 1584 5184 1602
rect 5166 1602 5184 1620
rect 5166 1620 5184 1638
rect 5166 1638 5184 1656
rect 5166 1656 5184 1674
rect 5166 1674 5184 1692
rect 5166 1692 5184 1710
rect 5166 1710 5184 1728
rect 5166 1728 5184 1746
rect 5166 1746 5184 1764
rect 5166 1764 5184 1782
rect 5166 1782 5184 1800
rect 5166 1800 5184 1818
rect 5166 1818 5184 1836
rect 5166 1836 5184 1854
rect 5166 1854 5184 1872
rect 5166 1872 5184 1890
rect 5166 1890 5184 1908
rect 5166 1908 5184 1926
rect 5166 1926 5184 1944
rect 5166 1944 5184 1962
rect 5166 1962 5184 1980
rect 5166 1980 5184 1998
rect 5166 1998 5184 2016
rect 5166 2016 5184 2034
rect 5166 2034 5184 2052
rect 5166 2052 5184 2070
rect 5166 2070 5184 2088
rect 5166 2088 5184 2106
rect 5166 2106 5184 2124
rect 5166 2124 5184 2142
rect 5166 2142 5184 2160
rect 5166 2160 5184 2178
rect 5166 2178 5184 2196
rect 5166 2196 5184 2214
rect 5166 2214 5184 2232
rect 5166 2232 5184 2250
rect 5166 2250 5184 2268
rect 5166 2268 5184 2286
rect 5166 2286 5184 2304
rect 5166 2304 5184 2322
rect 5166 2322 5184 2340
rect 5166 2538 5184 2556
rect 5166 2556 5184 2574
rect 5166 2574 5184 2592
rect 5166 2592 5184 2610
rect 5166 2610 5184 2628
rect 5166 2628 5184 2646
rect 5166 2646 5184 2664
rect 5166 2664 5184 2682
rect 5166 2682 5184 2700
rect 5166 2700 5184 2718
rect 5166 2718 5184 2736
rect 5166 2736 5184 2754
rect 5166 2754 5184 2772
rect 5166 2772 5184 2790
rect 5166 2790 5184 2808
rect 5166 2808 5184 2826
rect 5166 2826 5184 2844
rect 5166 2844 5184 2862
rect 5166 2862 5184 2880
rect 5166 2880 5184 2898
rect 5166 2898 5184 2916
rect 5166 2916 5184 2934
rect 5166 2934 5184 2952
rect 5166 2952 5184 2970
rect 5166 2970 5184 2988
rect 5166 2988 5184 3006
rect 5166 3006 5184 3024
rect 5166 3024 5184 3042
rect 5166 3042 5184 3060
rect 5166 3060 5184 3078
rect 5166 3078 5184 3096
rect 5166 3096 5184 3114
rect 5166 3114 5184 3132
rect 5166 3132 5184 3150
rect 5166 3150 5184 3168
rect 5166 3168 5184 3186
rect 5166 3186 5184 3204
rect 5166 3204 5184 3222
rect 5166 3222 5184 3240
rect 5166 3240 5184 3258
rect 5166 3258 5184 3276
rect 5166 3276 5184 3294
rect 5166 3294 5184 3312
rect 5166 3312 5184 3330
rect 5166 3330 5184 3348
rect 5166 3348 5184 3366
rect 5166 3366 5184 3384
rect 5166 3384 5184 3402
rect 5166 3402 5184 3420
rect 5166 3420 5184 3438
rect 5166 3438 5184 3456
rect 5166 3456 5184 3474
rect 5166 3474 5184 3492
rect 5166 3492 5184 3510
rect 5166 3510 5184 3528
rect 5166 3528 5184 3546
rect 5166 3546 5184 3564
rect 5166 3564 5184 3582
rect 5166 3582 5184 3600
rect 5166 3600 5184 3618
rect 5166 3618 5184 3636
rect 5166 3636 5184 3654
rect 5166 3654 5184 3672
rect 5166 3672 5184 3690
rect 5166 3690 5184 3708
rect 5166 3708 5184 3726
rect 5166 3726 5184 3744
rect 5166 3744 5184 3762
rect 5166 3762 5184 3780
rect 5166 3780 5184 3798
rect 5166 3798 5184 3816
rect 5166 3816 5184 3834
rect 5166 3834 5184 3852
rect 5166 3852 5184 3870
rect 5166 3870 5184 3888
rect 5166 3888 5184 3906
rect 5166 3906 5184 3924
rect 5166 3924 5184 3942
rect 5166 3942 5184 3960
rect 5166 3960 5184 3978
rect 5166 3978 5184 3996
rect 5166 3996 5184 4014
rect 5166 4014 5184 4032
rect 5166 4032 5184 4050
rect 5166 4050 5184 4068
rect 5166 4068 5184 4086
rect 5166 4086 5184 4104
rect 5166 4104 5184 4122
rect 5166 4122 5184 4140
rect 5166 4140 5184 4158
rect 5166 4158 5184 4176
rect 5166 4176 5184 4194
rect 5166 4194 5184 4212
rect 5166 4212 5184 4230
rect 5166 4230 5184 4248
rect 5166 4248 5184 4266
rect 5166 4266 5184 4284
rect 5166 4284 5184 4302
rect 5166 4302 5184 4320
rect 5166 4320 5184 4338
rect 5166 4338 5184 4356
rect 5166 4356 5184 4374
rect 5166 4374 5184 4392
rect 5166 4392 5184 4410
rect 5166 4410 5184 4428
rect 5166 4428 5184 4446
rect 5166 4446 5184 4464
rect 5166 4464 5184 4482
rect 5166 4482 5184 4500
rect 5166 4500 5184 4518
rect 5166 4518 5184 4536
rect 5166 4536 5184 4554
rect 5166 4770 5184 4788
rect 5166 4788 5184 4806
rect 5166 4806 5184 4824
rect 5166 4824 5184 4842
rect 5166 4842 5184 4860
rect 5166 4860 5184 4878
rect 5166 4878 5184 4896
rect 5166 4896 5184 4914
rect 5166 4914 5184 4932
rect 5166 4932 5184 4950
rect 5166 4950 5184 4968
rect 5166 4968 5184 4986
rect 5166 4986 5184 5004
rect 5166 5004 5184 5022
rect 5166 5022 5184 5040
rect 5166 5040 5184 5058
rect 5166 5058 5184 5076
rect 5166 5076 5184 5094
rect 5166 5094 5184 5112
rect 5166 5112 5184 5130
rect 5166 5130 5184 5148
rect 5166 5148 5184 5166
rect 5166 5166 5184 5184
rect 5166 5184 5184 5202
rect 5166 5202 5184 5220
rect 5166 5220 5184 5238
rect 5166 5238 5184 5256
rect 5166 5256 5184 5274
rect 5166 5274 5184 5292
rect 5166 5292 5184 5310
rect 5166 5310 5184 5328
rect 5166 5328 5184 5346
rect 5166 5346 5184 5364
rect 5166 5364 5184 5382
rect 5166 5382 5184 5400
rect 5166 5400 5184 5418
rect 5166 5418 5184 5436
rect 5166 5436 5184 5454
rect 5166 5454 5184 5472
rect 5166 5472 5184 5490
rect 5166 5490 5184 5508
rect 5166 5508 5184 5526
rect 5166 5526 5184 5544
rect 5166 5544 5184 5562
rect 5166 5562 5184 5580
rect 5166 5580 5184 5598
rect 5166 5598 5184 5616
rect 5166 5616 5184 5634
rect 5166 5634 5184 5652
rect 5166 5652 5184 5670
rect 5166 5670 5184 5688
rect 5166 5688 5184 5706
rect 5166 5706 5184 5724
rect 5166 5724 5184 5742
rect 5166 5742 5184 5760
rect 5166 5760 5184 5778
rect 5166 5778 5184 5796
rect 5166 5796 5184 5814
rect 5166 5814 5184 5832
rect 5166 5832 5184 5850
rect 5166 5850 5184 5868
rect 5166 5868 5184 5886
rect 5166 5886 5184 5904
rect 5166 5904 5184 5922
rect 5166 5922 5184 5940
rect 5166 5940 5184 5958
rect 5166 5958 5184 5976
rect 5166 5976 5184 5994
rect 5166 5994 5184 6012
rect 5166 6012 5184 6030
rect 5166 6030 5184 6048
rect 5166 6048 5184 6066
rect 5166 6066 5184 6084
rect 5166 6084 5184 6102
rect 5166 6102 5184 6120
rect 5166 6120 5184 6138
rect 5166 6138 5184 6156
rect 5166 6156 5184 6174
rect 5166 6174 5184 6192
rect 5166 6192 5184 6210
rect 5166 6210 5184 6228
rect 5166 6228 5184 6246
rect 5166 6246 5184 6264
rect 5166 6264 5184 6282
rect 5166 6282 5184 6300
rect 5166 6300 5184 6318
rect 5166 6318 5184 6336
rect 5166 6336 5184 6354
rect 5166 6354 5184 6372
rect 5166 6372 5184 6390
rect 5166 6390 5184 6408
rect 5166 6408 5184 6426
rect 5166 6426 5184 6444
rect 5166 6444 5184 6462
rect 5166 6462 5184 6480
rect 5166 6480 5184 6498
rect 5166 6498 5184 6516
rect 5166 6516 5184 6534
rect 5166 6534 5184 6552
rect 5166 6552 5184 6570
rect 5166 6570 5184 6588
rect 5166 6588 5184 6606
rect 5166 6606 5184 6624
rect 5166 6624 5184 6642
rect 5166 6642 5184 6660
rect 5166 6660 5184 6678
rect 5166 6678 5184 6696
rect 5166 6696 5184 6714
rect 5166 6714 5184 6732
rect 5166 6732 5184 6750
rect 5166 6750 5184 6768
rect 5166 6768 5184 6786
rect 5166 6786 5184 6804
rect 5166 6804 5184 6822
rect 5166 6822 5184 6840
rect 5166 6840 5184 6858
rect 5166 6858 5184 6876
rect 5166 6876 5184 6894
rect 5166 6894 5184 6912
rect 5166 6912 5184 6930
rect 5166 6930 5184 6948
rect 5166 6948 5184 6966
rect 5166 6966 5184 6984
rect 5166 6984 5184 7002
rect 5166 7002 5184 7020
rect 5166 7020 5184 7038
rect 5166 7038 5184 7056
rect 5166 7056 5184 7074
rect 5166 7074 5184 7092
rect 5166 7092 5184 7110
rect 5166 7110 5184 7128
rect 5166 7128 5184 7146
rect 5166 7146 5184 7164
rect 5166 7164 5184 7182
rect 5166 7182 5184 7200
rect 5166 7200 5184 7218
rect 5166 7218 5184 7236
rect 5166 7236 5184 7254
rect 5166 7254 5184 7272
rect 5166 7272 5184 7290
rect 5166 7290 5184 7308
rect 5166 7308 5184 7326
rect 5166 7326 5184 7344
rect 5166 7344 5184 7362
rect 5166 7362 5184 7380
rect 5166 7380 5184 7398
rect 5166 7398 5184 7416
rect 5166 7416 5184 7434
rect 5166 7434 5184 7452
rect 5166 7452 5184 7470
rect 5166 7470 5184 7488
rect 5166 7488 5184 7506
rect 5166 7506 5184 7524
rect 5166 7524 5184 7542
rect 5166 7542 5184 7560
rect 5166 7560 5184 7578
rect 5166 7578 5184 7596
rect 5166 7596 5184 7614
rect 5166 7614 5184 7632
rect 5166 7632 5184 7650
rect 5166 7650 5184 7668
rect 5166 7668 5184 7686
rect 5166 7686 5184 7704
rect 5166 7704 5184 7722
rect 5166 7722 5184 7740
rect 5166 7740 5184 7758
rect 5166 7758 5184 7776
rect 5166 7776 5184 7794
rect 5166 7794 5184 7812
rect 5166 7812 5184 7830
rect 5166 7830 5184 7848
rect 5166 7848 5184 7866
rect 5166 7866 5184 7884
rect 5166 7884 5184 7902
rect 5166 7902 5184 7920
rect 5166 7920 5184 7938
rect 5166 7938 5184 7956
rect 5166 7956 5184 7974
rect 5166 7974 5184 7992
rect 5166 7992 5184 8010
rect 5166 8010 5184 8028
rect 5166 8028 5184 8046
rect 5166 8046 5184 8064
rect 5166 8064 5184 8082
rect 5184 342 5202 360
rect 5184 360 5202 378
rect 5184 378 5202 396
rect 5184 396 5202 414
rect 5184 414 5202 432
rect 5184 432 5202 450
rect 5184 450 5202 468
rect 5184 468 5202 486
rect 5184 486 5202 504
rect 5184 504 5202 522
rect 5184 522 5202 540
rect 5184 540 5202 558
rect 5184 558 5202 576
rect 5184 576 5202 594
rect 5184 594 5202 612
rect 5184 612 5202 630
rect 5184 630 5202 648
rect 5184 648 5202 666
rect 5184 666 5202 684
rect 5184 684 5202 702
rect 5184 702 5202 720
rect 5184 720 5202 738
rect 5184 738 5202 756
rect 5184 756 5202 774
rect 5184 774 5202 792
rect 5184 792 5202 810
rect 5184 936 5202 954
rect 5184 954 5202 972
rect 5184 972 5202 990
rect 5184 990 5202 1008
rect 5184 1008 5202 1026
rect 5184 1026 5202 1044
rect 5184 1044 5202 1062
rect 5184 1062 5202 1080
rect 5184 1080 5202 1098
rect 5184 1098 5202 1116
rect 5184 1116 5202 1134
rect 5184 1134 5202 1152
rect 5184 1152 5202 1170
rect 5184 1170 5202 1188
rect 5184 1188 5202 1206
rect 5184 1206 5202 1224
rect 5184 1224 5202 1242
rect 5184 1242 5202 1260
rect 5184 1260 5202 1278
rect 5184 1278 5202 1296
rect 5184 1296 5202 1314
rect 5184 1314 5202 1332
rect 5184 1332 5202 1350
rect 5184 1350 5202 1368
rect 5184 1368 5202 1386
rect 5184 1386 5202 1404
rect 5184 1404 5202 1422
rect 5184 1422 5202 1440
rect 5184 1440 5202 1458
rect 5184 1458 5202 1476
rect 5184 1476 5202 1494
rect 5184 1494 5202 1512
rect 5184 1512 5202 1530
rect 5184 1530 5202 1548
rect 5184 1548 5202 1566
rect 5184 1566 5202 1584
rect 5184 1584 5202 1602
rect 5184 1602 5202 1620
rect 5184 1620 5202 1638
rect 5184 1638 5202 1656
rect 5184 1656 5202 1674
rect 5184 1674 5202 1692
rect 5184 1692 5202 1710
rect 5184 1710 5202 1728
rect 5184 1728 5202 1746
rect 5184 1746 5202 1764
rect 5184 1764 5202 1782
rect 5184 1782 5202 1800
rect 5184 1800 5202 1818
rect 5184 1818 5202 1836
rect 5184 1836 5202 1854
rect 5184 1854 5202 1872
rect 5184 1872 5202 1890
rect 5184 1890 5202 1908
rect 5184 1908 5202 1926
rect 5184 1926 5202 1944
rect 5184 1944 5202 1962
rect 5184 1962 5202 1980
rect 5184 1980 5202 1998
rect 5184 1998 5202 2016
rect 5184 2016 5202 2034
rect 5184 2034 5202 2052
rect 5184 2052 5202 2070
rect 5184 2070 5202 2088
rect 5184 2088 5202 2106
rect 5184 2106 5202 2124
rect 5184 2124 5202 2142
rect 5184 2142 5202 2160
rect 5184 2160 5202 2178
rect 5184 2178 5202 2196
rect 5184 2196 5202 2214
rect 5184 2214 5202 2232
rect 5184 2232 5202 2250
rect 5184 2250 5202 2268
rect 5184 2268 5202 2286
rect 5184 2286 5202 2304
rect 5184 2304 5202 2322
rect 5184 2322 5202 2340
rect 5184 2556 5202 2574
rect 5184 2574 5202 2592
rect 5184 2592 5202 2610
rect 5184 2610 5202 2628
rect 5184 2628 5202 2646
rect 5184 2646 5202 2664
rect 5184 2664 5202 2682
rect 5184 2682 5202 2700
rect 5184 2700 5202 2718
rect 5184 2718 5202 2736
rect 5184 2736 5202 2754
rect 5184 2754 5202 2772
rect 5184 2772 5202 2790
rect 5184 2790 5202 2808
rect 5184 2808 5202 2826
rect 5184 2826 5202 2844
rect 5184 2844 5202 2862
rect 5184 2862 5202 2880
rect 5184 2880 5202 2898
rect 5184 2898 5202 2916
rect 5184 2916 5202 2934
rect 5184 2934 5202 2952
rect 5184 2952 5202 2970
rect 5184 2970 5202 2988
rect 5184 2988 5202 3006
rect 5184 3006 5202 3024
rect 5184 3024 5202 3042
rect 5184 3042 5202 3060
rect 5184 3060 5202 3078
rect 5184 3078 5202 3096
rect 5184 3096 5202 3114
rect 5184 3114 5202 3132
rect 5184 3132 5202 3150
rect 5184 3150 5202 3168
rect 5184 3168 5202 3186
rect 5184 3186 5202 3204
rect 5184 3204 5202 3222
rect 5184 3222 5202 3240
rect 5184 3240 5202 3258
rect 5184 3258 5202 3276
rect 5184 3276 5202 3294
rect 5184 3294 5202 3312
rect 5184 3312 5202 3330
rect 5184 3330 5202 3348
rect 5184 3348 5202 3366
rect 5184 3366 5202 3384
rect 5184 3384 5202 3402
rect 5184 3402 5202 3420
rect 5184 3420 5202 3438
rect 5184 3438 5202 3456
rect 5184 3456 5202 3474
rect 5184 3474 5202 3492
rect 5184 3492 5202 3510
rect 5184 3510 5202 3528
rect 5184 3528 5202 3546
rect 5184 3546 5202 3564
rect 5184 3564 5202 3582
rect 5184 3582 5202 3600
rect 5184 3600 5202 3618
rect 5184 3618 5202 3636
rect 5184 3636 5202 3654
rect 5184 3654 5202 3672
rect 5184 3672 5202 3690
rect 5184 3690 5202 3708
rect 5184 3708 5202 3726
rect 5184 3726 5202 3744
rect 5184 3744 5202 3762
rect 5184 3762 5202 3780
rect 5184 3780 5202 3798
rect 5184 3798 5202 3816
rect 5184 3816 5202 3834
rect 5184 3834 5202 3852
rect 5184 3852 5202 3870
rect 5184 3870 5202 3888
rect 5184 3888 5202 3906
rect 5184 3906 5202 3924
rect 5184 3924 5202 3942
rect 5184 3942 5202 3960
rect 5184 3960 5202 3978
rect 5184 3978 5202 3996
rect 5184 3996 5202 4014
rect 5184 4014 5202 4032
rect 5184 4032 5202 4050
rect 5184 4050 5202 4068
rect 5184 4068 5202 4086
rect 5184 4086 5202 4104
rect 5184 4104 5202 4122
rect 5184 4122 5202 4140
rect 5184 4140 5202 4158
rect 5184 4158 5202 4176
rect 5184 4176 5202 4194
rect 5184 4194 5202 4212
rect 5184 4212 5202 4230
rect 5184 4230 5202 4248
rect 5184 4248 5202 4266
rect 5184 4266 5202 4284
rect 5184 4284 5202 4302
rect 5184 4302 5202 4320
rect 5184 4320 5202 4338
rect 5184 4338 5202 4356
rect 5184 4356 5202 4374
rect 5184 4374 5202 4392
rect 5184 4392 5202 4410
rect 5184 4410 5202 4428
rect 5184 4428 5202 4446
rect 5184 4446 5202 4464
rect 5184 4464 5202 4482
rect 5184 4482 5202 4500
rect 5184 4500 5202 4518
rect 5184 4518 5202 4536
rect 5184 4536 5202 4554
rect 5184 4554 5202 4572
rect 5184 4788 5202 4806
rect 5184 4806 5202 4824
rect 5184 4824 5202 4842
rect 5184 4842 5202 4860
rect 5184 4860 5202 4878
rect 5184 4878 5202 4896
rect 5184 4896 5202 4914
rect 5184 4914 5202 4932
rect 5184 4932 5202 4950
rect 5184 4950 5202 4968
rect 5184 4968 5202 4986
rect 5184 4986 5202 5004
rect 5184 5004 5202 5022
rect 5184 5022 5202 5040
rect 5184 5040 5202 5058
rect 5184 5058 5202 5076
rect 5184 5076 5202 5094
rect 5184 5094 5202 5112
rect 5184 5112 5202 5130
rect 5184 5130 5202 5148
rect 5184 5148 5202 5166
rect 5184 5166 5202 5184
rect 5184 5184 5202 5202
rect 5184 5202 5202 5220
rect 5184 5220 5202 5238
rect 5184 5238 5202 5256
rect 5184 5256 5202 5274
rect 5184 5274 5202 5292
rect 5184 5292 5202 5310
rect 5184 5310 5202 5328
rect 5184 5328 5202 5346
rect 5184 5346 5202 5364
rect 5184 5364 5202 5382
rect 5184 5382 5202 5400
rect 5184 5400 5202 5418
rect 5184 5418 5202 5436
rect 5184 5436 5202 5454
rect 5184 5454 5202 5472
rect 5184 5472 5202 5490
rect 5184 5490 5202 5508
rect 5184 5508 5202 5526
rect 5184 5526 5202 5544
rect 5184 5544 5202 5562
rect 5184 5562 5202 5580
rect 5184 5580 5202 5598
rect 5184 5598 5202 5616
rect 5184 5616 5202 5634
rect 5184 5634 5202 5652
rect 5184 5652 5202 5670
rect 5184 5670 5202 5688
rect 5184 5688 5202 5706
rect 5184 5706 5202 5724
rect 5184 5724 5202 5742
rect 5184 5742 5202 5760
rect 5184 5760 5202 5778
rect 5184 5778 5202 5796
rect 5184 5796 5202 5814
rect 5184 5814 5202 5832
rect 5184 5832 5202 5850
rect 5184 5850 5202 5868
rect 5184 5868 5202 5886
rect 5184 5886 5202 5904
rect 5184 5904 5202 5922
rect 5184 5922 5202 5940
rect 5184 5940 5202 5958
rect 5184 5958 5202 5976
rect 5184 5976 5202 5994
rect 5184 5994 5202 6012
rect 5184 6012 5202 6030
rect 5184 6030 5202 6048
rect 5184 6048 5202 6066
rect 5184 6066 5202 6084
rect 5184 6084 5202 6102
rect 5184 6102 5202 6120
rect 5184 6120 5202 6138
rect 5184 6138 5202 6156
rect 5184 6156 5202 6174
rect 5184 6174 5202 6192
rect 5184 6192 5202 6210
rect 5184 6210 5202 6228
rect 5184 6228 5202 6246
rect 5184 6246 5202 6264
rect 5184 6264 5202 6282
rect 5184 6282 5202 6300
rect 5184 6300 5202 6318
rect 5184 6318 5202 6336
rect 5184 6336 5202 6354
rect 5184 6354 5202 6372
rect 5184 6372 5202 6390
rect 5184 6390 5202 6408
rect 5184 6408 5202 6426
rect 5184 6426 5202 6444
rect 5184 6444 5202 6462
rect 5184 6462 5202 6480
rect 5184 6480 5202 6498
rect 5184 6498 5202 6516
rect 5184 6516 5202 6534
rect 5184 6534 5202 6552
rect 5184 6552 5202 6570
rect 5184 6570 5202 6588
rect 5184 6588 5202 6606
rect 5184 6606 5202 6624
rect 5184 6624 5202 6642
rect 5184 6642 5202 6660
rect 5184 6660 5202 6678
rect 5184 6678 5202 6696
rect 5184 6696 5202 6714
rect 5184 6714 5202 6732
rect 5184 6732 5202 6750
rect 5184 6750 5202 6768
rect 5184 6768 5202 6786
rect 5184 6786 5202 6804
rect 5184 6804 5202 6822
rect 5184 6822 5202 6840
rect 5184 6840 5202 6858
rect 5184 6858 5202 6876
rect 5184 6876 5202 6894
rect 5184 6894 5202 6912
rect 5184 6912 5202 6930
rect 5184 6930 5202 6948
rect 5184 6948 5202 6966
rect 5184 6966 5202 6984
rect 5184 6984 5202 7002
rect 5184 7002 5202 7020
rect 5184 7020 5202 7038
rect 5184 7038 5202 7056
rect 5184 7056 5202 7074
rect 5184 7074 5202 7092
rect 5184 7092 5202 7110
rect 5184 7110 5202 7128
rect 5184 7128 5202 7146
rect 5184 7146 5202 7164
rect 5184 7164 5202 7182
rect 5184 7182 5202 7200
rect 5184 7200 5202 7218
rect 5184 7218 5202 7236
rect 5184 7236 5202 7254
rect 5184 7254 5202 7272
rect 5184 7272 5202 7290
rect 5184 7290 5202 7308
rect 5184 7308 5202 7326
rect 5184 7326 5202 7344
rect 5184 7344 5202 7362
rect 5184 7362 5202 7380
rect 5184 7380 5202 7398
rect 5184 7398 5202 7416
rect 5184 7416 5202 7434
rect 5184 7434 5202 7452
rect 5184 7452 5202 7470
rect 5184 7470 5202 7488
rect 5184 7488 5202 7506
rect 5184 7506 5202 7524
rect 5184 7524 5202 7542
rect 5184 7542 5202 7560
rect 5184 7560 5202 7578
rect 5184 7578 5202 7596
rect 5184 7596 5202 7614
rect 5184 7614 5202 7632
rect 5184 7632 5202 7650
rect 5184 7650 5202 7668
rect 5184 7668 5202 7686
rect 5184 7686 5202 7704
rect 5184 7704 5202 7722
rect 5184 7722 5202 7740
rect 5184 7740 5202 7758
rect 5184 7758 5202 7776
rect 5184 7776 5202 7794
rect 5184 7794 5202 7812
rect 5184 7812 5202 7830
rect 5184 7830 5202 7848
rect 5184 7848 5202 7866
rect 5184 7866 5202 7884
rect 5184 7884 5202 7902
rect 5184 7902 5202 7920
rect 5184 7920 5202 7938
rect 5184 7938 5202 7956
rect 5184 7956 5202 7974
rect 5184 7974 5202 7992
rect 5184 7992 5202 8010
rect 5184 8010 5202 8028
rect 5184 8028 5202 8046
rect 5184 8046 5202 8064
rect 5184 8064 5202 8082
rect 5184 8082 5202 8100
rect 5184 8100 5202 8118
rect 5202 360 5220 378
rect 5202 378 5220 396
rect 5202 396 5220 414
rect 5202 414 5220 432
rect 5202 432 5220 450
rect 5202 450 5220 468
rect 5202 468 5220 486
rect 5202 486 5220 504
rect 5202 504 5220 522
rect 5202 522 5220 540
rect 5202 540 5220 558
rect 5202 558 5220 576
rect 5202 576 5220 594
rect 5202 594 5220 612
rect 5202 612 5220 630
rect 5202 630 5220 648
rect 5202 648 5220 666
rect 5202 666 5220 684
rect 5202 684 5220 702
rect 5202 702 5220 720
rect 5202 720 5220 738
rect 5202 738 5220 756
rect 5202 756 5220 774
rect 5202 774 5220 792
rect 5202 792 5220 810
rect 5202 936 5220 954
rect 5202 954 5220 972
rect 5202 972 5220 990
rect 5202 990 5220 1008
rect 5202 1008 5220 1026
rect 5202 1026 5220 1044
rect 5202 1044 5220 1062
rect 5202 1062 5220 1080
rect 5202 1080 5220 1098
rect 5202 1098 5220 1116
rect 5202 1116 5220 1134
rect 5202 1134 5220 1152
rect 5202 1152 5220 1170
rect 5202 1170 5220 1188
rect 5202 1188 5220 1206
rect 5202 1206 5220 1224
rect 5202 1224 5220 1242
rect 5202 1242 5220 1260
rect 5202 1260 5220 1278
rect 5202 1278 5220 1296
rect 5202 1296 5220 1314
rect 5202 1314 5220 1332
rect 5202 1332 5220 1350
rect 5202 1350 5220 1368
rect 5202 1368 5220 1386
rect 5202 1386 5220 1404
rect 5202 1404 5220 1422
rect 5202 1422 5220 1440
rect 5202 1440 5220 1458
rect 5202 1458 5220 1476
rect 5202 1476 5220 1494
rect 5202 1494 5220 1512
rect 5202 1512 5220 1530
rect 5202 1530 5220 1548
rect 5202 1548 5220 1566
rect 5202 1566 5220 1584
rect 5202 1584 5220 1602
rect 5202 1602 5220 1620
rect 5202 1620 5220 1638
rect 5202 1638 5220 1656
rect 5202 1656 5220 1674
rect 5202 1674 5220 1692
rect 5202 1692 5220 1710
rect 5202 1710 5220 1728
rect 5202 1728 5220 1746
rect 5202 1746 5220 1764
rect 5202 1764 5220 1782
rect 5202 1782 5220 1800
rect 5202 1800 5220 1818
rect 5202 1818 5220 1836
rect 5202 1836 5220 1854
rect 5202 1854 5220 1872
rect 5202 1872 5220 1890
rect 5202 1890 5220 1908
rect 5202 1908 5220 1926
rect 5202 1926 5220 1944
rect 5202 1944 5220 1962
rect 5202 1962 5220 1980
rect 5202 1980 5220 1998
rect 5202 1998 5220 2016
rect 5202 2016 5220 2034
rect 5202 2034 5220 2052
rect 5202 2052 5220 2070
rect 5202 2070 5220 2088
rect 5202 2088 5220 2106
rect 5202 2106 5220 2124
rect 5202 2124 5220 2142
rect 5202 2142 5220 2160
rect 5202 2160 5220 2178
rect 5202 2178 5220 2196
rect 5202 2196 5220 2214
rect 5202 2214 5220 2232
rect 5202 2232 5220 2250
rect 5202 2250 5220 2268
rect 5202 2268 5220 2286
rect 5202 2286 5220 2304
rect 5202 2304 5220 2322
rect 5202 2322 5220 2340
rect 5202 2340 5220 2358
rect 5202 2556 5220 2574
rect 5202 2574 5220 2592
rect 5202 2592 5220 2610
rect 5202 2610 5220 2628
rect 5202 2628 5220 2646
rect 5202 2646 5220 2664
rect 5202 2664 5220 2682
rect 5202 2682 5220 2700
rect 5202 2700 5220 2718
rect 5202 2718 5220 2736
rect 5202 2736 5220 2754
rect 5202 2754 5220 2772
rect 5202 2772 5220 2790
rect 5202 2790 5220 2808
rect 5202 2808 5220 2826
rect 5202 2826 5220 2844
rect 5202 2844 5220 2862
rect 5202 2862 5220 2880
rect 5202 2880 5220 2898
rect 5202 2898 5220 2916
rect 5202 2916 5220 2934
rect 5202 2934 5220 2952
rect 5202 2952 5220 2970
rect 5202 2970 5220 2988
rect 5202 2988 5220 3006
rect 5202 3006 5220 3024
rect 5202 3024 5220 3042
rect 5202 3042 5220 3060
rect 5202 3060 5220 3078
rect 5202 3078 5220 3096
rect 5202 3096 5220 3114
rect 5202 3114 5220 3132
rect 5202 3132 5220 3150
rect 5202 3150 5220 3168
rect 5202 3168 5220 3186
rect 5202 3186 5220 3204
rect 5202 3204 5220 3222
rect 5202 3222 5220 3240
rect 5202 3240 5220 3258
rect 5202 3258 5220 3276
rect 5202 3276 5220 3294
rect 5202 3294 5220 3312
rect 5202 3312 5220 3330
rect 5202 3330 5220 3348
rect 5202 3348 5220 3366
rect 5202 3366 5220 3384
rect 5202 3384 5220 3402
rect 5202 3402 5220 3420
rect 5202 3420 5220 3438
rect 5202 3438 5220 3456
rect 5202 3456 5220 3474
rect 5202 3474 5220 3492
rect 5202 3492 5220 3510
rect 5202 3510 5220 3528
rect 5202 3528 5220 3546
rect 5202 3546 5220 3564
rect 5202 3564 5220 3582
rect 5202 3582 5220 3600
rect 5202 3600 5220 3618
rect 5202 3618 5220 3636
rect 5202 3636 5220 3654
rect 5202 3654 5220 3672
rect 5202 3672 5220 3690
rect 5202 3690 5220 3708
rect 5202 3708 5220 3726
rect 5202 3726 5220 3744
rect 5202 3744 5220 3762
rect 5202 3762 5220 3780
rect 5202 3780 5220 3798
rect 5202 3798 5220 3816
rect 5202 3816 5220 3834
rect 5202 3834 5220 3852
rect 5202 3852 5220 3870
rect 5202 3870 5220 3888
rect 5202 3888 5220 3906
rect 5202 3906 5220 3924
rect 5202 3924 5220 3942
rect 5202 3942 5220 3960
rect 5202 3960 5220 3978
rect 5202 3978 5220 3996
rect 5202 3996 5220 4014
rect 5202 4014 5220 4032
rect 5202 4032 5220 4050
rect 5202 4050 5220 4068
rect 5202 4068 5220 4086
rect 5202 4086 5220 4104
rect 5202 4104 5220 4122
rect 5202 4122 5220 4140
rect 5202 4140 5220 4158
rect 5202 4158 5220 4176
rect 5202 4176 5220 4194
rect 5202 4194 5220 4212
rect 5202 4212 5220 4230
rect 5202 4230 5220 4248
rect 5202 4248 5220 4266
rect 5202 4266 5220 4284
rect 5202 4284 5220 4302
rect 5202 4302 5220 4320
rect 5202 4320 5220 4338
rect 5202 4338 5220 4356
rect 5202 4356 5220 4374
rect 5202 4374 5220 4392
rect 5202 4392 5220 4410
rect 5202 4410 5220 4428
rect 5202 4428 5220 4446
rect 5202 4446 5220 4464
rect 5202 4464 5220 4482
rect 5202 4482 5220 4500
rect 5202 4500 5220 4518
rect 5202 4518 5220 4536
rect 5202 4536 5220 4554
rect 5202 4554 5220 4572
rect 5202 4572 5220 4590
rect 5202 4590 5220 4608
rect 5202 4806 5220 4824
rect 5202 4824 5220 4842
rect 5202 4842 5220 4860
rect 5202 4860 5220 4878
rect 5202 4878 5220 4896
rect 5202 4896 5220 4914
rect 5202 4914 5220 4932
rect 5202 4932 5220 4950
rect 5202 4950 5220 4968
rect 5202 4968 5220 4986
rect 5202 4986 5220 5004
rect 5202 5004 5220 5022
rect 5202 5022 5220 5040
rect 5202 5040 5220 5058
rect 5202 5058 5220 5076
rect 5202 5076 5220 5094
rect 5202 5094 5220 5112
rect 5202 5112 5220 5130
rect 5202 5130 5220 5148
rect 5202 5148 5220 5166
rect 5202 5166 5220 5184
rect 5202 5184 5220 5202
rect 5202 5202 5220 5220
rect 5202 5220 5220 5238
rect 5202 5238 5220 5256
rect 5202 5256 5220 5274
rect 5202 5274 5220 5292
rect 5202 5292 5220 5310
rect 5202 5310 5220 5328
rect 5202 5328 5220 5346
rect 5202 5346 5220 5364
rect 5202 5364 5220 5382
rect 5202 5382 5220 5400
rect 5202 5400 5220 5418
rect 5202 5418 5220 5436
rect 5202 5436 5220 5454
rect 5202 5454 5220 5472
rect 5202 5472 5220 5490
rect 5202 5490 5220 5508
rect 5202 5508 5220 5526
rect 5202 5526 5220 5544
rect 5202 5544 5220 5562
rect 5202 5562 5220 5580
rect 5202 5580 5220 5598
rect 5202 5598 5220 5616
rect 5202 5616 5220 5634
rect 5202 5634 5220 5652
rect 5202 5652 5220 5670
rect 5202 5670 5220 5688
rect 5202 5688 5220 5706
rect 5202 5706 5220 5724
rect 5202 5724 5220 5742
rect 5202 5742 5220 5760
rect 5202 5760 5220 5778
rect 5202 5778 5220 5796
rect 5202 5796 5220 5814
rect 5202 5814 5220 5832
rect 5202 5832 5220 5850
rect 5202 5850 5220 5868
rect 5202 5868 5220 5886
rect 5202 5886 5220 5904
rect 5202 5904 5220 5922
rect 5202 5922 5220 5940
rect 5202 5940 5220 5958
rect 5202 5958 5220 5976
rect 5202 5976 5220 5994
rect 5202 5994 5220 6012
rect 5202 6012 5220 6030
rect 5202 6030 5220 6048
rect 5202 6048 5220 6066
rect 5202 6066 5220 6084
rect 5202 6084 5220 6102
rect 5202 6102 5220 6120
rect 5202 6120 5220 6138
rect 5202 6138 5220 6156
rect 5202 6156 5220 6174
rect 5202 6174 5220 6192
rect 5202 6192 5220 6210
rect 5202 6210 5220 6228
rect 5202 6228 5220 6246
rect 5202 6246 5220 6264
rect 5202 6264 5220 6282
rect 5202 6282 5220 6300
rect 5202 6300 5220 6318
rect 5202 6318 5220 6336
rect 5202 6336 5220 6354
rect 5202 6354 5220 6372
rect 5202 6372 5220 6390
rect 5202 6390 5220 6408
rect 5202 6408 5220 6426
rect 5202 6426 5220 6444
rect 5202 6444 5220 6462
rect 5202 6462 5220 6480
rect 5202 6480 5220 6498
rect 5202 6498 5220 6516
rect 5202 6516 5220 6534
rect 5202 6534 5220 6552
rect 5202 6552 5220 6570
rect 5202 6570 5220 6588
rect 5202 6588 5220 6606
rect 5202 6606 5220 6624
rect 5202 6624 5220 6642
rect 5202 6642 5220 6660
rect 5202 6660 5220 6678
rect 5202 6678 5220 6696
rect 5202 6696 5220 6714
rect 5202 6714 5220 6732
rect 5202 6732 5220 6750
rect 5202 6750 5220 6768
rect 5202 6768 5220 6786
rect 5202 6786 5220 6804
rect 5202 6804 5220 6822
rect 5202 6822 5220 6840
rect 5202 6840 5220 6858
rect 5202 6858 5220 6876
rect 5202 6876 5220 6894
rect 5202 6894 5220 6912
rect 5202 6912 5220 6930
rect 5202 6930 5220 6948
rect 5202 6948 5220 6966
rect 5202 6966 5220 6984
rect 5202 6984 5220 7002
rect 5202 7002 5220 7020
rect 5202 7020 5220 7038
rect 5202 7038 5220 7056
rect 5202 7056 5220 7074
rect 5202 7074 5220 7092
rect 5202 7092 5220 7110
rect 5202 7110 5220 7128
rect 5202 7128 5220 7146
rect 5202 7146 5220 7164
rect 5202 7164 5220 7182
rect 5202 7182 5220 7200
rect 5202 7200 5220 7218
rect 5202 7218 5220 7236
rect 5202 7236 5220 7254
rect 5202 7254 5220 7272
rect 5202 7272 5220 7290
rect 5202 7290 5220 7308
rect 5202 7308 5220 7326
rect 5202 7326 5220 7344
rect 5202 7344 5220 7362
rect 5202 7362 5220 7380
rect 5202 7380 5220 7398
rect 5202 7398 5220 7416
rect 5202 7416 5220 7434
rect 5202 7434 5220 7452
rect 5202 7452 5220 7470
rect 5202 7470 5220 7488
rect 5202 7488 5220 7506
rect 5202 7506 5220 7524
rect 5202 7524 5220 7542
rect 5202 7542 5220 7560
rect 5202 7560 5220 7578
rect 5202 7578 5220 7596
rect 5202 7596 5220 7614
rect 5202 7614 5220 7632
rect 5202 7632 5220 7650
rect 5202 7650 5220 7668
rect 5202 7668 5220 7686
rect 5202 7686 5220 7704
rect 5202 7704 5220 7722
rect 5202 7722 5220 7740
rect 5202 7740 5220 7758
rect 5202 7758 5220 7776
rect 5202 7776 5220 7794
rect 5202 7794 5220 7812
rect 5202 7812 5220 7830
rect 5202 7830 5220 7848
rect 5202 7848 5220 7866
rect 5202 7866 5220 7884
rect 5202 7884 5220 7902
rect 5202 7902 5220 7920
rect 5202 7920 5220 7938
rect 5202 7938 5220 7956
rect 5202 7956 5220 7974
rect 5202 7974 5220 7992
rect 5202 7992 5220 8010
rect 5202 8010 5220 8028
rect 5202 8028 5220 8046
rect 5202 8046 5220 8064
rect 5202 8064 5220 8082
rect 5202 8082 5220 8100
rect 5202 8100 5220 8118
rect 5202 8118 5220 8136
rect 5220 360 5238 378
rect 5220 378 5238 396
rect 5220 396 5238 414
rect 5220 414 5238 432
rect 5220 432 5238 450
rect 5220 450 5238 468
rect 5220 468 5238 486
rect 5220 486 5238 504
rect 5220 504 5238 522
rect 5220 522 5238 540
rect 5220 540 5238 558
rect 5220 558 5238 576
rect 5220 576 5238 594
rect 5220 594 5238 612
rect 5220 612 5238 630
rect 5220 630 5238 648
rect 5220 648 5238 666
rect 5220 666 5238 684
rect 5220 684 5238 702
rect 5220 702 5238 720
rect 5220 720 5238 738
rect 5220 738 5238 756
rect 5220 756 5238 774
rect 5220 774 5238 792
rect 5220 792 5238 810
rect 5220 954 5238 972
rect 5220 972 5238 990
rect 5220 990 5238 1008
rect 5220 1008 5238 1026
rect 5220 1026 5238 1044
rect 5220 1044 5238 1062
rect 5220 1062 5238 1080
rect 5220 1080 5238 1098
rect 5220 1098 5238 1116
rect 5220 1116 5238 1134
rect 5220 1134 5238 1152
rect 5220 1152 5238 1170
rect 5220 1170 5238 1188
rect 5220 1188 5238 1206
rect 5220 1206 5238 1224
rect 5220 1224 5238 1242
rect 5220 1242 5238 1260
rect 5220 1260 5238 1278
rect 5220 1278 5238 1296
rect 5220 1296 5238 1314
rect 5220 1314 5238 1332
rect 5220 1332 5238 1350
rect 5220 1350 5238 1368
rect 5220 1368 5238 1386
rect 5220 1386 5238 1404
rect 5220 1404 5238 1422
rect 5220 1422 5238 1440
rect 5220 1440 5238 1458
rect 5220 1458 5238 1476
rect 5220 1476 5238 1494
rect 5220 1494 5238 1512
rect 5220 1512 5238 1530
rect 5220 1530 5238 1548
rect 5220 1548 5238 1566
rect 5220 1566 5238 1584
rect 5220 1584 5238 1602
rect 5220 1602 5238 1620
rect 5220 1620 5238 1638
rect 5220 1638 5238 1656
rect 5220 1656 5238 1674
rect 5220 1674 5238 1692
rect 5220 1692 5238 1710
rect 5220 1710 5238 1728
rect 5220 1728 5238 1746
rect 5220 1746 5238 1764
rect 5220 1764 5238 1782
rect 5220 1782 5238 1800
rect 5220 1800 5238 1818
rect 5220 1818 5238 1836
rect 5220 1836 5238 1854
rect 5220 1854 5238 1872
rect 5220 1872 5238 1890
rect 5220 1890 5238 1908
rect 5220 1908 5238 1926
rect 5220 1926 5238 1944
rect 5220 1944 5238 1962
rect 5220 1962 5238 1980
rect 5220 1980 5238 1998
rect 5220 1998 5238 2016
rect 5220 2016 5238 2034
rect 5220 2034 5238 2052
rect 5220 2052 5238 2070
rect 5220 2070 5238 2088
rect 5220 2088 5238 2106
rect 5220 2106 5238 2124
rect 5220 2124 5238 2142
rect 5220 2142 5238 2160
rect 5220 2160 5238 2178
rect 5220 2178 5238 2196
rect 5220 2196 5238 2214
rect 5220 2214 5238 2232
rect 5220 2232 5238 2250
rect 5220 2250 5238 2268
rect 5220 2268 5238 2286
rect 5220 2286 5238 2304
rect 5220 2304 5238 2322
rect 5220 2322 5238 2340
rect 5220 2340 5238 2358
rect 5220 2574 5238 2592
rect 5220 2592 5238 2610
rect 5220 2610 5238 2628
rect 5220 2628 5238 2646
rect 5220 2646 5238 2664
rect 5220 2664 5238 2682
rect 5220 2682 5238 2700
rect 5220 2700 5238 2718
rect 5220 2718 5238 2736
rect 5220 2736 5238 2754
rect 5220 2754 5238 2772
rect 5220 2772 5238 2790
rect 5220 2790 5238 2808
rect 5220 2808 5238 2826
rect 5220 2826 5238 2844
rect 5220 2844 5238 2862
rect 5220 2862 5238 2880
rect 5220 2880 5238 2898
rect 5220 2898 5238 2916
rect 5220 2916 5238 2934
rect 5220 2934 5238 2952
rect 5220 2952 5238 2970
rect 5220 2970 5238 2988
rect 5220 2988 5238 3006
rect 5220 3006 5238 3024
rect 5220 3024 5238 3042
rect 5220 3042 5238 3060
rect 5220 3060 5238 3078
rect 5220 3078 5238 3096
rect 5220 3096 5238 3114
rect 5220 3114 5238 3132
rect 5220 3132 5238 3150
rect 5220 3150 5238 3168
rect 5220 3168 5238 3186
rect 5220 3186 5238 3204
rect 5220 3204 5238 3222
rect 5220 3222 5238 3240
rect 5220 3240 5238 3258
rect 5220 3258 5238 3276
rect 5220 3276 5238 3294
rect 5220 3294 5238 3312
rect 5220 3312 5238 3330
rect 5220 3330 5238 3348
rect 5220 3348 5238 3366
rect 5220 3366 5238 3384
rect 5220 3384 5238 3402
rect 5220 3402 5238 3420
rect 5220 3420 5238 3438
rect 5220 3438 5238 3456
rect 5220 3456 5238 3474
rect 5220 3474 5238 3492
rect 5220 3492 5238 3510
rect 5220 3510 5238 3528
rect 5220 3528 5238 3546
rect 5220 3546 5238 3564
rect 5220 3564 5238 3582
rect 5220 3582 5238 3600
rect 5220 3600 5238 3618
rect 5220 3618 5238 3636
rect 5220 3636 5238 3654
rect 5220 3654 5238 3672
rect 5220 3672 5238 3690
rect 5220 3690 5238 3708
rect 5220 3708 5238 3726
rect 5220 3726 5238 3744
rect 5220 3744 5238 3762
rect 5220 3762 5238 3780
rect 5220 3780 5238 3798
rect 5220 3798 5238 3816
rect 5220 3816 5238 3834
rect 5220 3834 5238 3852
rect 5220 3852 5238 3870
rect 5220 3870 5238 3888
rect 5220 3888 5238 3906
rect 5220 3906 5238 3924
rect 5220 3924 5238 3942
rect 5220 3942 5238 3960
rect 5220 3960 5238 3978
rect 5220 3978 5238 3996
rect 5220 3996 5238 4014
rect 5220 4014 5238 4032
rect 5220 4032 5238 4050
rect 5220 4050 5238 4068
rect 5220 4068 5238 4086
rect 5220 4086 5238 4104
rect 5220 4104 5238 4122
rect 5220 4122 5238 4140
rect 5220 4140 5238 4158
rect 5220 4158 5238 4176
rect 5220 4176 5238 4194
rect 5220 4194 5238 4212
rect 5220 4212 5238 4230
rect 5220 4230 5238 4248
rect 5220 4248 5238 4266
rect 5220 4266 5238 4284
rect 5220 4284 5238 4302
rect 5220 4302 5238 4320
rect 5220 4320 5238 4338
rect 5220 4338 5238 4356
rect 5220 4356 5238 4374
rect 5220 4374 5238 4392
rect 5220 4392 5238 4410
rect 5220 4410 5238 4428
rect 5220 4428 5238 4446
rect 5220 4446 5238 4464
rect 5220 4464 5238 4482
rect 5220 4482 5238 4500
rect 5220 4500 5238 4518
rect 5220 4518 5238 4536
rect 5220 4536 5238 4554
rect 5220 4554 5238 4572
rect 5220 4572 5238 4590
rect 5220 4590 5238 4608
rect 5220 4608 5238 4626
rect 5220 4824 5238 4842
rect 5220 4842 5238 4860
rect 5220 4860 5238 4878
rect 5220 4878 5238 4896
rect 5220 4896 5238 4914
rect 5220 4914 5238 4932
rect 5220 4932 5238 4950
rect 5220 4950 5238 4968
rect 5220 4968 5238 4986
rect 5220 4986 5238 5004
rect 5220 5004 5238 5022
rect 5220 5022 5238 5040
rect 5220 5040 5238 5058
rect 5220 5058 5238 5076
rect 5220 5076 5238 5094
rect 5220 5094 5238 5112
rect 5220 5112 5238 5130
rect 5220 5130 5238 5148
rect 5220 5148 5238 5166
rect 5220 5166 5238 5184
rect 5220 5184 5238 5202
rect 5220 5202 5238 5220
rect 5220 5220 5238 5238
rect 5220 5238 5238 5256
rect 5220 5256 5238 5274
rect 5220 5274 5238 5292
rect 5220 5292 5238 5310
rect 5220 5310 5238 5328
rect 5220 5328 5238 5346
rect 5220 5346 5238 5364
rect 5220 5364 5238 5382
rect 5220 5382 5238 5400
rect 5220 5400 5238 5418
rect 5220 5418 5238 5436
rect 5220 5436 5238 5454
rect 5220 5454 5238 5472
rect 5220 5472 5238 5490
rect 5220 5490 5238 5508
rect 5220 5508 5238 5526
rect 5220 5526 5238 5544
rect 5220 5544 5238 5562
rect 5220 5562 5238 5580
rect 5220 5580 5238 5598
rect 5220 5598 5238 5616
rect 5220 5616 5238 5634
rect 5220 5634 5238 5652
rect 5220 5652 5238 5670
rect 5220 5670 5238 5688
rect 5220 5688 5238 5706
rect 5220 5706 5238 5724
rect 5220 5724 5238 5742
rect 5220 5742 5238 5760
rect 5220 5760 5238 5778
rect 5220 5778 5238 5796
rect 5220 5796 5238 5814
rect 5220 5814 5238 5832
rect 5220 5832 5238 5850
rect 5220 5850 5238 5868
rect 5220 5868 5238 5886
rect 5220 5886 5238 5904
rect 5220 5904 5238 5922
rect 5220 5922 5238 5940
rect 5220 5940 5238 5958
rect 5220 5958 5238 5976
rect 5220 5976 5238 5994
rect 5220 5994 5238 6012
rect 5220 6012 5238 6030
rect 5220 6030 5238 6048
rect 5220 6048 5238 6066
rect 5220 6066 5238 6084
rect 5220 6084 5238 6102
rect 5220 6102 5238 6120
rect 5220 6120 5238 6138
rect 5220 6138 5238 6156
rect 5220 6156 5238 6174
rect 5220 6174 5238 6192
rect 5220 6192 5238 6210
rect 5220 6210 5238 6228
rect 5220 6228 5238 6246
rect 5220 6246 5238 6264
rect 5220 6264 5238 6282
rect 5220 6282 5238 6300
rect 5220 6300 5238 6318
rect 5220 6318 5238 6336
rect 5220 6336 5238 6354
rect 5220 6354 5238 6372
rect 5220 6372 5238 6390
rect 5220 6390 5238 6408
rect 5220 6408 5238 6426
rect 5220 6426 5238 6444
rect 5220 6444 5238 6462
rect 5220 6462 5238 6480
rect 5220 6480 5238 6498
rect 5220 6498 5238 6516
rect 5220 6516 5238 6534
rect 5220 6534 5238 6552
rect 5220 6552 5238 6570
rect 5220 6570 5238 6588
rect 5220 6588 5238 6606
rect 5220 6606 5238 6624
rect 5220 6624 5238 6642
rect 5220 6642 5238 6660
rect 5220 6660 5238 6678
rect 5220 6678 5238 6696
rect 5220 6696 5238 6714
rect 5220 6714 5238 6732
rect 5220 6732 5238 6750
rect 5220 6750 5238 6768
rect 5220 6768 5238 6786
rect 5220 6786 5238 6804
rect 5220 6804 5238 6822
rect 5220 6822 5238 6840
rect 5220 6840 5238 6858
rect 5220 6858 5238 6876
rect 5220 6876 5238 6894
rect 5220 6894 5238 6912
rect 5220 6912 5238 6930
rect 5220 6930 5238 6948
rect 5220 6948 5238 6966
rect 5220 6966 5238 6984
rect 5220 6984 5238 7002
rect 5220 7002 5238 7020
rect 5220 7020 5238 7038
rect 5220 7038 5238 7056
rect 5220 7056 5238 7074
rect 5220 7074 5238 7092
rect 5220 7092 5238 7110
rect 5220 7110 5238 7128
rect 5220 7128 5238 7146
rect 5220 7146 5238 7164
rect 5220 7164 5238 7182
rect 5220 7182 5238 7200
rect 5220 7200 5238 7218
rect 5220 7218 5238 7236
rect 5220 7236 5238 7254
rect 5220 7254 5238 7272
rect 5220 7272 5238 7290
rect 5220 7290 5238 7308
rect 5220 7308 5238 7326
rect 5220 7326 5238 7344
rect 5220 7344 5238 7362
rect 5220 7362 5238 7380
rect 5220 7380 5238 7398
rect 5220 7398 5238 7416
rect 5220 7416 5238 7434
rect 5220 7434 5238 7452
rect 5220 7452 5238 7470
rect 5220 7470 5238 7488
rect 5220 7488 5238 7506
rect 5220 7506 5238 7524
rect 5220 7524 5238 7542
rect 5220 7542 5238 7560
rect 5220 7560 5238 7578
rect 5220 7578 5238 7596
rect 5220 7596 5238 7614
rect 5220 7614 5238 7632
rect 5220 7632 5238 7650
rect 5220 7650 5238 7668
rect 5220 7668 5238 7686
rect 5220 7686 5238 7704
rect 5220 7704 5238 7722
rect 5220 7722 5238 7740
rect 5220 7740 5238 7758
rect 5220 7758 5238 7776
rect 5220 7776 5238 7794
rect 5220 7794 5238 7812
rect 5220 7812 5238 7830
rect 5220 7830 5238 7848
rect 5220 7848 5238 7866
rect 5220 7866 5238 7884
rect 5220 7884 5238 7902
rect 5220 7902 5238 7920
rect 5220 7920 5238 7938
rect 5220 7938 5238 7956
rect 5220 7956 5238 7974
rect 5220 7974 5238 7992
rect 5220 7992 5238 8010
rect 5220 8010 5238 8028
rect 5220 8028 5238 8046
rect 5220 8046 5238 8064
rect 5220 8064 5238 8082
rect 5220 8082 5238 8100
rect 5220 8100 5238 8118
rect 5220 8118 5238 8136
rect 5220 8136 5238 8154
rect 5220 8154 5238 8172
rect 5238 378 5256 396
rect 5238 396 5256 414
rect 5238 414 5256 432
rect 5238 432 5256 450
rect 5238 450 5256 468
rect 5238 468 5256 486
rect 5238 486 5256 504
rect 5238 504 5256 522
rect 5238 522 5256 540
rect 5238 540 5256 558
rect 5238 558 5256 576
rect 5238 576 5256 594
rect 5238 594 5256 612
rect 5238 612 5256 630
rect 5238 630 5256 648
rect 5238 648 5256 666
rect 5238 666 5256 684
rect 5238 684 5256 702
rect 5238 702 5256 720
rect 5238 720 5256 738
rect 5238 738 5256 756
rect 5238 756 5256 774
rect 5238 774 5256 792
rect 5238 792 5256 810
rect 5238 810 5256 828
rect 5238 954 5256 972
rect 5238 972 5256 990
rect 5238 990 5256 1008
rect 5238 1008 5256 1026
rect 5238 1026 5256 1044
rect 5238 1044 5256 1062
rect 5238 1062 5256 1080
rect 5238 1080 5256 1098
rect 5238 1098 5256 1116
rect 5238 1116 5256 1134
rect 5238 1134 5256 1152
rect 5238 1152 5256 1170
rect 5238 1170 5256 1188
rect 5238 1188 5256 1206
rect 5238 1206 5256 1224
rect 5238 1224 5256 1242
rect 5238 1242 5256 1260
rect 5238 1260 5256 1278
rect 5238 1278 5256 1296
rect 5238 1296 5256 1314
rect 5238 1314 5256 1332
rect 5238 1332 5256 1350
rect 5238 1350 5256 1368
rect 5238 1368 5256 1386
rect 5238 1386 5256 1404
rect 5238 1404 5256 1422
rect 5238 1422 5256 1440
rect 5238 1440 5256 1458
rect 5238 1458 5256 1476
rect 5238 1476 5256 1494
rect 5238 1494 5256 1512
rect 5238 1512 5256 1530
rect 5238 1530 5256 1548
rect 5238 1548 5256 1566
rect 5238 1566 5256 1584
rect 5238 1584 5256 1602
rect 5238 1602 5256 1620
rect 5238 1620 5256 1638
rect 5238 1638 5256 1656
rect 5238 1656 5256 1674
rect 5238 1674 5256 1692
rect 5238 1692 5256 1710
rect 5238 1710 5256 1728
rect 5238 1728 5256 1746
rect 5238 1746 5256 1764
rect 5238 1764 5256 1782
rect 5238 1782 5256 1800
rect 5238 1800 5256 1818
rect 5238 1818 5256 1836
rect 5238 1836 5256 1854
rect 5238 1854 5256 1872
rect 5238 1872 5256 1890
rect 5238 1890 5256 1908
rect 5238 1908 5256 1926
rect 5238 1926 5256 1944
rect 5238 1944 5256 1962
rect 5238 1962 5256 1980
rect 5238 1980 5256 1998
rect 5238 1998 5256 2016
rect 5238 2016 5256 2034
rect 5238 2034 5256 2052
rect 5238 2052 5256 2070
rect 5238 2070 5256 2088
rect 5238 2088 5256 2106
rect 5238 2106 5256 2124
rect 5238 2124 5256 2142
rect 5238 2142 5256 2160
rect 5238 2160 5256 2178
rect 5238 2178 5256 2196
rect 5238 2196 5256 2214
rect 5238 2214 5256 2232
rect 5238 2232 5256 2250
rect 5238 2250 5256 2268
rect 5238 2268 5256 2286
rect 5238 2286 5256 2304
rect 5238 2304 5256 2322
rect 5238 2322 5256 2340
rect 5238 2340 5256 2358
rect 5238 2358 5256 2376
rect 5238 2574 5256 2592
rect 5238 2592 5256 2610
rect 5238 2610 5256 2628
rect 5238 2628 5256 2646
rect 5238 2646 5256 2664
rect 5238 2664 5256 2682
rect 5238 2682 5256 2700
rect 5238 2700 5256 2718
rect 5238 2718 5256 2736
rect 5238 2736 5256 2754
rect 5238 2754 5256 2772
rect 5238 2772 5256 2790
rect 5238 2790 5256 2808
rect 5238 2808 5256 2826
rect 5238 2826 5256 2844
rect 5238 2844 5256 2862
rect 5238 2862 5256 2880
rect 5238 2880 5256 2898
rect 5238 2898 5256 2916
rect 5238 2916 5256 2934
rect 5238 2934 5256 2952
rect 5238 2952 5256 2970
rect 5238 2970 5256 2988
rect 5238 2988 5256 3006
rect 5238 3006 5256 3024
rect 5238 3024 5256 3042
rect 5238 3042 5256 3060
rect 5238 3060 5256 3078
rect 5238 3078 5256 3096
rect 5238 3096 5256 3114
rect 5238 3114 5256 3132
rect 5238 3132 5256 3150
rect 5238 3150 5256 3168
rect 5238 3168 5256 3186
rect 5238 3186 5256 3204
rect 5238 3204 5256 3222
rect 5238 3222 5256 3240
rect 5238 3240 5256 3258
rect 5238 3258 5256 3276
rect 5238 3276 5256 3294
rect 5238 3294 5256 3312
rect 5238 3312 5256 3330
rect 5238 3330 5256 3348
rect 5238 3348 5256 3366
rect 5238 3366 5256 3384
rect 5238 3384 5256 3402
rect 5238 3402 5256 3420
rect 5238 3420 5256 3438
rect 5238 3438 5256 3456
rect 5238 3456 5256 3474
rect 5238 3474 5256 3492
rect 5238 3492 5256 3510
rect 5238 3510 5256 3528
rect 5238 3528 5256 3546
rect 5238 3546 5256 3564
rect 5238 3564 5256 3582
rect 5238 3582 5256 3600
rect 5238 3600 5256 3618
rect 5238 3618 5256 3636
rect 5238 3636 5256 3654
rect 5238 3654 5256 3672
rect 5238 3672 5256 3690
rect 5238 3690 5256 3708
rect 5238 3708 5256 3726
rect 5238 3726 5256 3744
rect 5238 3744 5256 3762
rect 5238 3762 5256 3780
rect 5238 3780 5256 3798
rect 5238 3798 5256 3816
rect 5238 3816 5256 3834
rect 5238 3834 5256 3852
rect 5238 3852 5256 3870
rect 5238 3870 5256 3888
rect 5238 3888 5256 3906
rect 5238 3906 5256 3924
rect 5238 3924 5256 3942
rect 5238 3942 5256 3960
rect 5238 3960 5256 3978
rect 5238 3978 5256 3996
rect 5238 3996 5256 4014
rect 5238 4014 5256 4032
rect 5238 4032 5256 4050
rect 5238 4050 5256 4068
rect 5238 4068 5256 4086
rect 5238 4086 5256 4104
rect 5238 4104 5256 4122
rect 5238 4122 5256 4140
rect 5238 4140 5256 4158
rect 5238 4158 5256 4176
rect 5238 4176 5256 4194
rect 5238 4194 5256 4212
rect 5238 4212 5256 4230
rect 5238 4230 5256 4248
rect 5238 4248 5256 4266
rect 5238 4266 5256 4284
rect 5238 4284 5256 4302
rect 5238 4302 5256 4320
rect 5238 4320 5256 4338
rect 5238 4338 5256 4356
rect 5238 4356 5256 4374
rect 5238 4374 5256 4392
rect 5238 4392 5256 4410
rect 5238 4410 5256 4428
rect 5238 4428 5256 4446
rect 5238 4446 5256 4464
rect 5238 4464 5256 4482
rect 5238 4482 5256 4500
rect 5238 4500 5256 4518
rect 5238 4518 5256 4536
rect 5238 4536 5256 4554
rect 5238 4554 5256 4572
rect 5238 4572 5256 4590
rect 5238 4590 5256 4608
rect 5238 4608 5256 4626
rect 5238 4626 5256 4644
rect 5238 4842 5256 4860
rect 5238 4860 5256 4878
rect 5238 4878 5256 4896
rect 5238 4896 5256 4914
rect 5238 4914 5256 4932
rect 5238 4932 5256 4950
rect 5238 4950 5256 4968
rect 5238 4968 5256 4986
rect 5238 4986 5256 5004
rect 5238 5004 5256 5022
rect 5238 5022 5256 5040
rect 5238 5040 5256 5058
rect 5238 5058 5256 5076
rect 5238 5076 5256 5094
rect 5238 5094 5256 5112
rect 5238 5112 5256 5130
rect 5238 5130 5256 5148
rect 5238 5148 5256 5166
rect 5238 5166 5256 5184
rect 5238 5184 5256 5202
rect 5238 5202 5256 5220
rect 5238 5220 5256 5238
rect 5238 5238 5256 5256
rect 5238 5256 5256 5274
rect 5238 5274 5256 5292
rect 5238 5292 5256 5310
rect 5238 5310 5256 5328
rect 5238 5328 5256 5346
rect 5238 5346 5256 5364
rect 5238 5364 5256 5382
rect 5238 5382 5256 5400
rect 5238 5400 5256 5418
rect 5238 5418 5256 5436
rect 5238 5436 5256 5454
rect 5238 5454 5256 5472
rect 5238 5472 5256 5490
rect 5238 5490 5256 5508
rect 5238 5508 5256 5526
rect 5238 5526 5256 5544
rect 5238 5544 5256 5562
rect 5238 5562 5256 5580
rect 5238 5580 5256 5598
rect 5238 5598 5256 5616
rect 5238 5616 5256 5634
rect 5238 5634 5256 5652
rect 5238 5652 5256 5670
rect 5238 5670 5256 5688
rect 5238 5688 5256 5706
rect 5238 5706 5256 5724
rect 5238 5724 5256 5742
rect 5238 5742 5256 5760
rect 5238 5760 5256 5778
rect 5238 5778 5256 5796
rect 5238 5796 5256 5814
rect 5238 5814 5256 5832
rect 5238 5832 5256 5850
rect 5238 5850 5256 5868
rect 5238 5868 5256 5886
rect 5238 5886 5256 5904
rect 5238 5904 5256 5922
rect 5238 5922 5256 5940
rect 5238 5940 5256 5958
rect 5238 5958 5256 5976
rect 5238 5976 5256 5994
rect 5238 5994 5256 6012
rect 5238 6012 5256 6030
rect 5238 6030 5256 6048
rect 5238 6048 5256 6066
rect 5238 6066 5256 6084
rect 5238 6084 5256 6102
rect 5238 6102 5256 6120
rect 5238 6120 5256 6138
rect 5238 6138 5256 6156
rect 5238 6156 5256 6174
rect 5238 6174 5256 6192
rect 5238 6192 5256 6210
rect 5238 6210 5256 6228
rect 5238 6228 5256 6246
rect 5238 6246 5256 6264
rect 5238 6264 5256 6282
rect 5238 6282 5256 6300
rect 5238 6300 5256 6318
rect 5238 6318 5256 6336
rect 5238 6336 5256 6354
rect 5238 6354 5256 6372
rect 5238 6372 5256 6390
rect 5238 6390 5256 6408
rect 5238 6408 5256 6426
rect 5238 6426 5256 6444
rect 5238 6444 5256 6462
rect 5238 6462 5256 6480
rect 5238 6480 5256 6498
rect 5238 6498 5256 6516
rect 5238 6516 5256 6534
rect 5238 6534 5256 6552
rect 5238 6552 5256 6570
rect 5238 6570 5256 6588
rect 5238 6588 5256 6606
rect 5238 6606 5256 6624
rect 5238 6624 5256 6642
rect 5238 6642 5256 6660
rect 5238 6660 5256 6678
rect 5238 6678 5256 6696
rect 5238 6696 5256 6714
rect 5238 6714 5256 6732
rect 5238 6732 5256 6750
rect 5238 6750 5256 6768
rect 5238 6768 5256 6786
rect 5238 6786 5256 6804
rect 5238 6804 5256 6822
rect 5238 6822 5256 6840
rect 5238 6840 5256 6858
rect 5238 6858 5256 6876
rect 5238 6876 5256 6894
rect 5238 6894 5256 6912
rect 5238 6912 5256 6930
rect 5238 6930 5256 6948
rect 5238 6948 5256 6966
rect 5238 6966 5256 6984
rect 5238 6984 5256 7002
rect 5238 7002 5256 7020
rect 5238 7020 5256 7038
rect 5238 7038 5256 7056
rect 5238 7056 5256 7074
rect 5238 7074 5256 7092
rect 5238 7092 5256 7110
rect 5238 7110 5256 7128
rect 5238 7128 5256 7146
rect 5238 7146 5256 7164
rect 5238 7164 5256 7182
rect 5238 7182 5256 7200
rect 5238 7200 5256 7218
rect 5238 7218 5256 7236
rect 5238 7236 5256 7254
rect 5238 7254 5256 7272
rect 5238 7272 5256 7290
rect 5238 7290 5256 7308
rect 5238 7308 5256 7326
rect 5238 7326 5256 7344
rect 5238 7344 5256 7362
rect 5238 7362 5256 7380
rect 5238 7380 5256 7398
rect 5238 7398 5256 7416
rect 5238 7416 5256 7434
rect 5238 7434 5256 7452
rect 5238 7452 5256 7470
rect 5238 7470 5256 7488
rect 5238 7488 5256 7506
rect 5238 7506 5256 7524
rect 5238 7524 5256 7542
rect 5238 7542 5256 7560
rect 5238 7560 5256 7578
rect 5238 7578 5256 7596
rect 5238 7596 5256 7614
rect 5238 7614 5256 7632
rect 5238 7632 5256 7650
rect 5238 7650 5256 7668
rect 5238 7668 5256 7686
rect 5238 7686 5256 7704
rect 5238 7704 5256 7722
rect 5238 7722 5256 7740
rect 5238 7740 5256 7758
rect 5238 7758 5256 7776
rect 5238 7776 5256 7794
rect 5238 7794 5256 7812
rect 5238 7812 5256 7830
rect 5238 7830 5256 7848
rect 5238 7848 5256 7866
rect 5238 7866 5256 7884
rect 5238 7884 5256 7902
rect 5238 7902 5256 7920
rect 5238 7920 5256 7938
rect 5238 7938 5256 7956
rect 5238 7956 5256 7974
rect 5238 7974 5256 7992
rect 5238 7992 5256 8010
rect 5238 8010 5256 8028
rect 5238 8028 5256 8046
rect 5238 8046 5256 8064
rect 5238 8064 5256 8082
rect 5238 8082 5256 8100
rect 5238 8100 5256 8118
rect 5238 8118 5256 8136
rect 5238 8136 5256 8154
rect 5238 8154 5256 8172
rect 5238 8172 5256 8190
rect 5256 378 5274 396
rect 5256 396 5274 414
rect 5256 414 5274 432
rect 5256 432 5274 450
rect 5256 450 5274 468
rect 5256 468 5274 486
rect 5256 486 5274 504
rect 5256 504 5274 522
rect 5256 522 5274 540
rect 5256 540 5274 558
rect 5256 558 5274 576
rect 5256 576 5274 594
rect 5256 594 5274 612
rect 5256 612 5274 630
rect 5256 630 5274 648
rect 5256 648 5274 666
rect 5256 666 5274 684
rect 5256 684 5274 702
rect 5256 702 5274 720
rect 5256 720 5274 738
rect 5256 738 5274 756
rect 5256 756 5274 774
rect 5256 774 5274 792
rect 5256 792 5274 810
rect 5256 810 5274 828
rect 5256 954 5274 972
rect 5256 972 5274 990
rect 5256 990 5274 1008
rect 5256 1008 5274 1026
rect 5256 1026 5274 1044
rect 5256 1044 5274 1062
rect 5256 1062 5274 1080
rect 5256 1080 5274 1098
rect 5256 1098 5274 1116
rect 5256 1116 5274 1134
rect 5256 1134 5274 1152
rect 5256 1152 5274 1170
rect 5256 1170 5274 1188
rect 5256 1188 5274 1206
rect 5256 1206 5274 1224
rect 5256 1224 5274 1242
rect 5256 1242 5274 1260
rect 5256 1260 5274 1278
rect 5256 1278 5274 1296
rect 5256 1296 5274 1314
rect 5256 1314 5274 1332
rect 5256 1332 5274 1350
rect 5256 1350 5274 1368
rect 5256 1368 5274 1386
rect 5256 1386 5274 1404
rect 5256 1404 5274 1422
rect 5256 1422 5274 1440
rect 5256 1440 5274 1458
rect 5256 1458 5274 1476
rect 5256 1476 5274 1494
rect 5256 1494 5274 1512
rect 5256 1512 5274 1530
rect 5256 1530 5274 1548
rect 5256 1548 5274 1566
rect 5256 1566 5274 1584
rect 5256 1584 5274 1602
rect 5256 1602 5274 1620
rect 5256 1620 5274 1638
rect 5256 1638 5274 1656
rect 5256 1656 5274 1674
rect 5256 1674 5274 1692
rect 5256 1692 5274 1710
rect 5256 1710 5274 1728
rect 5256 1728 5274 1746
rect 5256 1746 5274 1764
rect 5256 1764 5274 1782
rect 5256 1782 5274 1800
rect 5256 1800 5274 1818
rect 5256 1818 5274 1836
rect 5256 1836 5274 1854
rect 5256 1854 5274 1872
rect 5256 1872 5274 1890
rect 5256 1890 5274 1908
rect 5256 1908 5274 1926
rect 5256 1926 5274 1944
rect 5256 1944 5274 1962
rect 5256 1962 5274 1980
rect 5256 1980 5274 1998
rect 5256 1998 5274 2016
rect 5256 2016 5274 2034
rect 5256 2034 5274 2052
rect 5256 2052 5274 2070
rect 5256 2070 5274 2088
rect 5256 2088 5274 2106
rect 5256 2106 5274 2124
rect 5256 2124 5274 2142
rect 5256 2142 5274 2160
rect 5256 2160 5274 2178
rect 5256 2178 5274 2196
rect 5256 2196 5274 2214
rect 5256 2214 5274 2232
rect 5256 2232 5274 2250
rect 5256 2250 5274 2268
rect 5256 2268 5274 2286
rect 5256 2286 5274 2304
rect 5256 2304 5274 2322
rect 5256 2322 5274 2340
rect 5256 2340 5274 2358
rect 5256 2358 5274 2376
rect 5256 2592 5274 2610
rect 5256 2610 5274 2628
rect 5256 2628 5274 2646
rect 5256 2646 5274 2664
rect 5256 2664 5274 2682
rect 5256 2682 5274 2700
rect 5256 2700 5274 2718
rect 5256 2718 5274 2736
rect 5256 2736 5274 2754
rect 5256 2754 5274 2772
rect 5256 2772 5274 2790
rect 5256 2790 5274 2808
rect 5256 2808 5274 2826
rect 5256 2826 5274 2844
rect 5256 2844 5274 2862
rect 5256 2862 5274 2880
rect 5256 2880 5274 2898
rect 5256 2898 5274 2916
rect 5256 2916 5274 2934
rect 5256 2934 5274 2952
rect 5256 2952 5274 2970
rect 5256 2970 5274 2988
rect 5256 2988 5274 3006
rect 5256 3006 5274 3024
rect 5256 3024 5274 3042
rect 5256 3042 5274 3060
rect 5256 3060 5274 3078
rect 5256 3078 5274 3096
rect 5256 3096 5274 3114
rect 5256 3114 5274 3132
rect 5256 3132 5274 3150
rect 5256 3150 5274 3168
rect 5256 3168 5274 3186
rect 5256 3186 5274 3204
rect 5256 3204 5274 3222
rect 5256 3222 5274 3240
rect 5256 3240 5274 3258
rect 5256 3258 5274 3276
rect 5256 3276 5274 3294
rect 5256 3294 5274 3312
rect 5256 3312 5274 3330
rect 5256 3330 5274 3348
rect 5256 3348 5274 3366
rect 5256 3366 5274 3384
rect 5256 3384 5274 3402
rect 5256 3402 5274 3420
rect 5256 3420 5274 3438
rect 5256 3438 5274 3456
rect 5256 3456 5274 3474
rect 5256 3474 5274 3492
rect 5256 3492 5274 3510
rect 5256 3510 5274 3528
rect 5256 3528 5274 3546
rect 5256 3546 5274 3564
rect 5256 3564 5274 3582
rect 5256 3582 5274 3600
rect 5256 3600 5274 3618
rect 5256 3618 5274 3636
rect 5256 3636 5274 3654
rect 5256 3654 5274 3672
rect 5256 3672 5274 3690
rect 5256 3690 5274 3708
rect 5256 3708 5274 3726
rect 5256 3726 5274 3744
rect 5256 3744 5274 3762
rect 5256 3762 5274 3780
rect 5256 3780 5274 3798
rect 5256 3798 5274 3816
rect 5256 3816 5274 3834
rect 5256 3834 5274 3852
rect 5256 3852 5274 3870
rect 5256 3870 5274 3888
rect 5256 3888 5274 3906
rect 5256 3906 5274 3924
rect 5256 3924 5274 3942
rect 5256 3942 5274 3960
rect 5256 3960 5274 3978
rect 5256 3978 5274 3996
rect 5256 3996 5274 4014
rect 5256 4014 5274 4032
rect 5256 4032 5274 4050
rect 5256 4050 5274 4068
rect 5256 4068 5274 4086
rect 5256 4086 5274 4104
rect 5256 4104 5274 4122
rect 5256 4122 5274 4140
rect 5256 4140 5274 4158
rect 5256 4158 5274 4176
rect 5256 4176 5274 4194
rect 5256 4194 5274 4212
rect 5256 4212 5274 4230
rect 5256 4230 5274 4248
rect 5256 4248 5274 4266
rect 5256 4266 5274 4284
rect 5256 4284 5274 4302
rect 5256 4302 5274 4320
rect 5256 4320 5274 4338
rect 5256 4338 5274 4356
rect 5256 4356 5274 4374
rect 5256 4374 5274 4392
rect 5256 4392 5274 4410
rect 5256 4410 5274 4428
rect 5256 4428 5274 4446
rect 5256 4446 5274 4464
rect 5256 4464 5274 4482
rect 5256 4482 5274 4500
rect 5256 4500 5274 4518
rect 5256 4518 5274 4536
rect 5256 4536 5274 4554
rect 5256 4554 5274 4572
rect 5256 4572 5274 4590
rect 5256 4590 5274 4608
rect 5256 4608 5274 4626
rect 5256 4626 5274 4644
rect 5256 4644 5274 4662
rect 5256 4878 5274 4896
rect 5256 4896 5274 4914
rect 5256 4914 5274 4932
rect 5256 4932 5274 4950
rect 5256 4950 5274 4968
rect 5256 4968 5274 4986
rect 5256 4986 5274 5004
rect 5256 5004 5274 5022
rect 5256 5022 5274 5040
rect 5256 5040 5274 5058
rect 5256 5058 5274 5076
rect 5256 5076 5274 5094
rect 5256 5094 5274 5112
rect 5256 5112 5274 5130
rect 5256 5130 5274 5148
rect 5256 5148 5274 5166
rect 5256 5166 5274 5184
rect 5256 5184 5274 5202
rect 5256 5202 5274 5220
rect 5256 5220 5274 5238
rect 5256 5238 5274 5256
rect 5256 5256 5274 5274
rect 5256 5274 5274 5292
rect 5256 5292 5274 5310
rect 5256 5310 5274 5328
rect 5256 5328 5274 5346
rect 5256 5346 5274 5364
rect 5256 5364 5274 5382
rect 5256 5382 5274 5400
rect 5256 5400 5274 5418
rect 5256 5418 5274 5436
rect 5256 5436 5274 5454
rect 5256 5454 5274 5472
rect 5256 5472 5274 5490
rect 5256 5490 5274 5508
rect 5256 5508 5274 5526
rect 5256 5526 5274 5544
rect 5256 5544 5274 5562
rect 5256 5562 5274 5580
rect 5256 5580 5274 5598
rect 5256 5598 5274 5616
rect 5256 5616 5274 5634
rect 5256 5634 5274 5652
rect 5256 5652 5274 5670
rect 5256 5670 5274 5688
rect 5256 5688 5274 5706
rect 5256 5706 5274 5724
rect 5256 5724 5274 5742
rect 5256 5742 5274 5760
rect 5256 5760 5274 5778
rect 5256 5778 5274 5796
rect 5256 5796 5274 5814
rect 5256 5814 5274 5832
rect 5256 5832 5274 5850
rect 5256 5850 5274 5868
rect 5256 5868 5274 5886
rect 5256 5886 5274 5904
rect 5256 5904 5274 5922
rect 5256 5922 5274 5940
rect 5256 5940 5274 5958
rect 5256 5958 5274 5976
rect 5256 5976 5274 5994
rect 5256 5994 5274 6012
rect 5256 6012 5274 6030
rect 5256 6030 5274 6048
rect 5256 6048 5274 6066
rect 5256 6066 5274 6084
rect 5256 6084 5274 6102
rect 5256 6102 5274 6120
rect 5256 6120 5274 6138
rect 5256 6138 5274 6156
rect 5256 6156 5274 6174
rect 5256 6174 5274 6192
rect 5256 6192 5274 6210
rect 5256 6210 5274 6228
rect 5256 6228 5274 6246
rect 5256 6246 5274 6264
rect 5256 6264 5274 6282
rect 5256 6282 5274 6300
rect 5256 6300 5274 6318
rect 5256 6318 5274 6336
rect 5256 6336 5274 6354
rect 5256 6354 5274 6372
rect 5256 6372 5274 6390
rect 5256 6390 5274 6408
rect 5256 6408 5274 6426
rect 5256 6426 5274 6444
rect 5256 6444 5274 6462
rect 5256 6462 5274 6480
rect 5256 6480 5274 6498
rect 5256 6498 5274 6516
rect 5256 6516 5274 6534
rect 5256 6534 5274 6552
rect 5256 6552 5274 6570
rect 5256 6570 5274 6588
rect 5256 6588 5274 6606
rect 5256 6606 5274 6624
rect 5256 6624 5274 6642
rect 5256 6642 5274 6660
rect 5256 6660 5274 6678
rect 5256 6678 5274 6696
rect 5256 6696 5274 6714
rect 5256 6714 5274 6732
rect 5256 6732 5274 6750
rect 5256 6750 5274 6768
rect 5256 6768 5274 6786
rect 5256 6786 5274 6804
rect 5256 6804 5274 6822
rect 5256 6822 5274 6840
rect 5256 6840 5274 6858
rect 5256 6858 5274 6876
rect 5256 6876 5274 6894
rect 5256 6894 5274 6912
rect 5256 6912 5274 6930
rect 5256 6930 5274 6948
rect 5256 6948 5274 6966
rect 5256 6966 5274 6984
rect 5256 6984 5274 7002
rect 5256 7002 5274 7020
rect 5256 7020 5274 7038
rect 5256 7038 5274 7056
rect 5256 7056 5274 7074
rect 5256 7074 5274 7092
rect 5256 7092 5274 7110
rect 5256 7110 5274 7128
rect 5256 7128 5274 7146
rect 5256 7146 5274 7164
rect 5256 7164 5274 7182
rect 5256 7182 5274 7200
rect 5256 7200 5274 7218
rect 5256 7218 5274 7236
rect 5256 7236 5274 7254
rect 5256 7254 5274 7272
rect 5256 7272 5274 7290
rect 5256 7290 5274 7308
rect 5256 7308 5274 7326
rect 5256 7326 5274 7344
rect 5256 7344 5274 7362
rect 5256 7362 5274 7380
rect 5256 7380 5274 7398
rect 5256 7398 5274 7416
rect 5256 7416 5274 7434
rect 5256 7434 5274 7452
rect 5256 7452 5274 7470
rect 5256 7470 5274 7488
rect 5256 7488 5274 7506
rect 5256 7506 5274 7524
rect 5256 7524 5274 7542
rect 5256 7542 5274 7560
rect 5256 7560 5274 7578
rect 5256 7578 5274 7596
rect 5256 7596 5274 7614
rect 5256 7614 5274 7632
rect 5256 7632 5274 7650
rect 5256 7650 5274 7668
rect 5256 7668 5274 7686
rect 5256 7686 5274 7704
rect 5256 7704 5274 7722
rect 5256 7722 5274 7740
rect 5256 7740 5274 7758
rect 5256 7758 5274 7776
rect 5256 7776 5274 7794
rect 5256 7794 5274 7812
rect 5256 7812 5274 7830
rect 5256 7830 5274 7848
rect 5256 7848 5274 7866
rect 5256 7866 5274 7884
rect 5256 7884 5274 7902
rect 5256 7902 5274 7920
rect 5256 7920 5274 7938
rect 5256 7938 5274 7956
rect 5256 7956 5274 7974
rect 5256 7974 5274 7992
rect 5256 7992 5274 8010
rect 5256 8010 5274 8028
rect 5256 8028 5274 8046
rect 5256 8046 5274 8064
rect 5256 8064 5274 8082
rect 5256 8082 5274 8100
rect 5256 8100 5274 8118
rect 5256 8118 5274 8136
rect 5256 8136 5274 8154
rect 5256 8154 5274 8172
rect 5256 8172 5274 8190
rect 5256 8190 5274 8208
rect 5256 8208 5274 8226
rect 5274 396 5292 414
rect 5274 414 5292 432
rect 5274 432 5292 450
rect 5274 450 5292 468
rect 5274 468 5292 486
rect 5274 486 5292 504
rect 5274 504 5292 522
rect 5274 522 5292 540
rect 5274 540 5292 558
rect 5274 558 5292 576
rect 5274 576 5292 594
rect 5274 594 5292 612
rect 5274 612 5292 630
rect 5274 630 5292 648
rect 5274 648 5292 666
rect 5274 666 5292 684
rect 5274 684 5292 702
rect 5274 702 5292 720
rect 5274 720 5292 738
rect 5274 738 5292 756
rect 5274 756 5292 774
rect 5274 774 5292 792
rect 5274 792 5292 810
rect 5274 810 5292 828
rect 5274 972 5292 990
rect 5274 990 5292 1008
rect 5274 1008 5292 1026
rect 5274 1026 5292 1044
rect 5274 1044 5292 1062
rect 5274 1062 5292 1080
rect 5274 1080 5292 1098
rect 5274 1098 5292 1116
rect 5274 1116 5292 1134
rect 5274 1134 5292 1152
rect 5274 1152 5292 1170
rect 5274 1170 5292 1188
rect 5274 1188 5292 1206
rect 5274 1206 5292 1224
rect 5274 1224 5292 1242
rect 5274 1242 5292 1260
rect 5274 1260 5292 1278
rect 5274 1278 5292 1296
rect 5274 1296 5292 1314
rect 5274 1314 5292 1332
rect 5274 1332 5292 1350
rect 5274 1350 5292 1368
rect 5274 1368 5292 1386
rect 5274 1386 5292 1404
rect 5274 1404 5292 1422
rect 5274 1422 5292 1440
rect 5274 1440 5292 1458
rect 5274 1458 5292 1476
rect 5274 1476 5292 1494
rect 5274 1494 5292 1512
rect 5274 1512 5292 1530
rect 5274 1530 5292 1548
rect 5274 1548 5292 1566
rect 5274 1566 5292 1584
rect 5274 1584 5292 1602
rect 5274 1602 5292 1620
rect 5274 1620 5292 1638
rect 5274 1638 5292 1656
rect 5274 1656 5292 1674
rect 5274 1674 5292 1692
rect 5274 1692 5292 1710
rect 5274 1710 5292 1728
rect 5274 1728 5292 1746
rect 5274 1746 5292 1764
rect 5274 1764 5292 1782
rect 5274 1782 5292 1800
rect 5274 1800 5292 1818
rect 5274 1818 5292 1836
rect 5274 1836 5292 1854
rect 5274 1854 5292 1872
rect 5274 1872 5292 1890
rect 5274 1890 5292 1908
rect 5274 1908 5292 1926
rect 5274 1926 5292 1944
rect 5274 1944 5292 1962
rect 5274 1962 5292 1980
rect 5274 1980 5292 1998
rect 5274 1998 5292 2016
rect 5274 2016 5292 2034
rect 5274 2034 5292 2052
rect 5274 2052 5292 2070
rect 5274 2070 5292 2088
rect 5274 2088 5292 2106
rect 5274 2106 5292 2124
rect 5274 2124 5292 2142
rect 5274 2142 5292 2160
rect 5274 2160 5292 2178
rect 5274 2178 5292 2196
rect 5274 2196 5292 2214
rect 5274 2214 5292 2232
rect 5274 2232 5292 2250
rect 5274 2250 5292 2268
rect 5274 2268 5292 2286
rect 5274 2286 5292 2304
rect 5274 2304 5292 2322
rect 5274 2322 5292 2340
rect 5274 2340 5292 2358
rect 5274 2358 5292 2376
rect 5274 2376 5292 2394
rect 5274 2592 5292 2610
rect 5274 2610 5292 2628
rect 5274 2628 5292 2646
rect 5274 2646 5292 2664
rect 5274 2664 5292 2682
rect 5274 2682 5292 2700
rect 5274 2700 5292 2718
rect 5274 2718 5292 2736
rect 5274 2736 5292 2754
rect 5274 2754 5292 2772
rect 5274 2772 5292 2790
rect 5274 2790 5292 2808
rect 5274 2808 5292 2826
rect 5274 2826 5292 2844
rect 5274 2844 5292 2862
rect 5274 2862 5292 2880
rect 5274 2880 5292 2898
rect 5274 2898 5292 2916
rect 5274 2916 5292 2934
rect 5274 2934 5292 2952
rect 5274 2952 5292 2970
rect 5274 2970 5292 2988
rect 5274 2988 5292 3006
rect 5274 3006 5292 3024
rect 5274 3024 5292 3042
rect 5274 3042 5292 3060
rect 5274 3060 5292 3078
rect 5274 3078 5292 3096
rect 5274 3096 5292 3114
rect 5274 3114 5292 3132
rect 5274 3132 5292 3150
rect 5274 3150 5292 3168
rect 5274 3168 5292 3186
rect 5274 3186 5292 3204
rect 5274 3204 5292 3222
rect 5274 3222 5292 3240
rect 5274 3240 5292 3258
rect 5274 3258 5292 3276
rect 5274 3276 5292 3294
rect 5274 3294 5292 3312
rect 5274 3312 5292 3330
rect 5274 3330 5292 3348
rect 5274 3348 5292 3366
rect 5274 3366 5292 3384
rect 5274 3384 5292 3402
rect 5274 3402 5292 3420
rect 5274 3420 5292 3438
rect 5274 3438 5292 3456
rect 5274 3456 5292 3474
rect 5274 3474 5292 3492
rect 5274 3492 5292 3510
rect 5274 3510 5292 3528
rect 5274 3528 5292 3546
rect 5274 3546 5292 3564
rect 5274 3564 5292 3582
rect 5274 3582 5292 3600
rect 5274 3600 5292 3618
rect 5274 3618 5292 3636
rect 5274 3636 5292 3654
rect 5274 3654 5292 3672
rect 5274 3672 5292 3690
rect 5274 3690 5292 3708
rect 5274 3708 5292 3726
rect 5274 3726 5292 3744
rect 5274 3744 5292 3762
rect 5274 3762 5292 3780
rect 5274 3780 5292 3798
rect 5274 3798 5292 3816
rect 5274 3816 5292 3834
rect 5274 3834 5292 3852
rect 5274 3852 5292 3870
rect 5274 3870 5292 3888
rect 5274 3888 5292 3906
rect 5274 3906 5292 3924
rect 5274 3924 5292 3942
rect 5274 3942 5292 3960
rect 5274 3960 5292 3978
rect 5274 3978 5292 3996
rect 5274 3996 5292 4014
rect 5274 4014 5292 4032
rect 5274 4032 5292 4050
rect 5274 4050 5292 4068
rect 5274 4068 5292 4086
rect 5274 4086 5292 4104
rect 5274 4104 5292 4122
rect 5274 4122 5292 4140
rect 5274 4140 5292 4158
rect 5274 4158 5292 4176
rect 5274 4176 5292 4194
rect 5274 4194 5292 4212
rect 5274 4212 5292 4230
rect 5274 4230 5292 4248
rect 5274 4248 5292 4266
rect 5274 4266 5292 4284
rect 5274 4284 5292 4302
rect 5274 4302 5292 4320
rect 5274 4320 5292 4338
rect 5274 4338 5292 4356
rect 5274 4356 5292 4374
rect 5274 4374 5292 4392
rect 5274 4392 5292 4410
rect 5274 4410 5292 4428
rect 5274 4428 5292 4446
rect 5274 4446 5292 4464
rect 5274 4464 5292 4482
rect 5274 4482 5292 4500
rect 5274 4500 5292 4518
rect 5274 4518 5292 4536
rect 5274 4536 5292 4554
rect 5274 4554 5292 4572
rect 5274 4572 5292 4590
rect 5274 4590 5292 4608
rect 5274 4608 5292 4626
rect 5274 4626 5292 4644
rect 5274 4644 5292 4662
rect 5274 4662 5292 4680
rect 5274 4896 5292 4914
rect 5274 4914 5292 4932
rect 5274 4932 5292 4950
rect 5274 4950 5292 4968
rect 5274 4968 5292 4986
rect 5274 4986 5292 5004
rect 5274 5004 5292 5022
rect 5274 5022 5292 5040
rect 5274 5040 5292 5058
rect 5274 5058 5292 5076
rect 5274 5076 5292 5094
rect 5274 5094 5292 5112
rect 5274 5112 5292 5130
rect 5274 5130 5292 5148
rect 5274 5148 5292 5166
rect 5274 5166 5292 5184
rect 5274 5184 5292 5202
rect 5274 5202 5292 5220
rect 5274 5220 5292 5238
rect 5274 5238 5292 5256
rect 5274 5256 5292 5274
rect 5274 5274 5292 5292
rect 5274 5292 5292 5310
rect 5274 5310 5292 5328
rect 5274 5328 5292 5346
rect 5274 5346 5292 5364
rect 5274 5364 5292 5382
rect 5274 5382 5292 5400
rect 5274 5400 5292 5418
rect 5274 5418 5292 5436
rect 5274 5436 5292 5454
rect 5274 5454 5292 5472
rect 5274 5472 5292 5490
rect 5274 5490 5292 5508
rect 5274 5508 5292 5526
rect 5274 5526 5292 5544
rect 5274 5544 5292 5562
rect 5274 5562 5292 5580
rect 5274 5580 5292 5598
rect 5274 5598 5292 5616
rect 5274 5616 5292 5634
rect 5274 5634 5292 5652
rect 5274 5652 5292 5670
rect 5274 5670 5292 5688
rect 5274 5688 5292 5706
rect 5274 5706 5292 5724
rect 5274 5724 5292 5742
rect 5274 5742 5292 5760
rect 5274 5760 5292 5778
rect 5274 5778 5292 5796
rect 5274 5796 5292 5814
rect 5274 5814 5292 5832
rect 5274 5832 5292 5850
rect 5274 5850 5292 5868
rect 5274 5868 5292 5886
rect 5274 5886 5292 5904
rect 5274 5904 5292 5922
rect 5274 5922 5292 5940
rect 5274 5940 5292 5958
rect 5274 5958 5292 5976
rect 5274 5976 5292 5994
rect 5274 5994 5292 6012
rect 5274 6012 5292 6030
rect 5274 6030 5292 6048
rect 5274 6048 5292 6066
rect 5274 6066 5292 6084
rect 5274 6084 5292 6102
rect 5274 6102 5292 6120
rect 5274 6120 5292 6138
rect 5274 6138 5292 6156
rect 5274 6156 5292 6174
rect 5274 6174 5292 6192
rect 5274 6192 5292 6210
rect 5274 6210 5292 6228
rect 5274 6228 5292 6246
rect 5274 6246 5292 6264
rect 5274 6264 5292 6282
rect 5274 6282 5292 6300
rect 5274 6300 5292 6318
rect 5274 6318 5292 6336
rect 5274 6336 5292 6354
rect 5274 6354 5292 6372
rect 5274 6372 5292 6390
rect 5274 6390 5292 6408
rect 5274 6408 5292 6426
rect 5274 6426 5292 6444
rect 5274 6444 5292 6462
rect 5274 6462 5292 6480
rect 5274 6480 5292 6498
rect 5274 6498 5292 6516
rect 5274 6516 5292 6534
rect 5274 6534 5292 6552
rect 5274 6552 5292 6570
rect 5274 6570 5292 6588
rect 5274 6588 5292 6606
rect 5274 6606 5292 6624
rect 5274 6624 5292 6642
rect 5274 6642 5292 6660
rect 5274 6660 5292 6678
rect 5274 6678 5292 6696
rect 5274 6696 5292 6714
rect 5274 6714 5292 6732
rect 5274 6732 5292 6750
rect 5274 6750 5292 6768
rect 5274 6768 5292 6786
rect 5274 6786 5292 6804
rect 5274 6804 5292 6822
rect 5274 6822 5292 6840
rect 5274 6840 5292 6858
rect 5274 6858 5292 6876
rect 5274 6876 5292 6894
rect 5274 6894 5292 6912
rect 5274 6912 5292 6930
rect 5274 6930 5292 6948
rect 5274 6948 5292 6966
rect 5274 6966 5292 6984
rect 5274 6984 5292 7002
rect 5274 7002 5292 7020
rect 5274 7020 5292 7038
rect 5274 7038 5292 7056
rect 5274 7056 5292 7074
rect 5274 7074 5292 7092
rect 5274 7092 5292 7110
rect 5274 7110 5292 7128
rect 5274 7128 5292 7146
rect 5274 7146 5292 7164
rect 5274 7164 5292 7182
rect 5274 7182 5292 7200
rect 5274 7200 5292 7218
rect 5274 7218 5292 7236
rect 5274 7236 5292 7254
rect 5274 7254 5292 7272
rect 5274 7272 5292 7290
rect 5274 7290 5292 7308
rect 5274 7308 5292 7326
rect 5274 7326 5292 7344
rect 5274 7344 5292 7362
rect 5274 7362 5292 7380
rect 5274 7380 5292 7398
rect 5274 7398 5292 7416
rect 5274 7416 5292 7434
rect 5274 7434 5292 7452
rect 5274 7452 5292 7470
rect 5274 7470 5292 7488
rect 5274 7488 5292 7506
rect 5274 7506 5292 7524
rect 5274 7524 5292 7542
rect 5274 7542 5292 7560
rect 5274 7560 5292 7578
rect 5274 7578 5292 7596
rect 5274 7596 5292 7614
rect 5274 7614 5292 7632
rect 5274 7632 5292 7650
rect 5274 7650 5292 7668
rect 5274 7668 5292 7686
rect 5274 7686 5292 7704
rect 5274 7704 5292 7722
rect 5274 7722 5292 7740
rect 5274 7740 5292 7758
rect 5274 7758 5292 7776
rect 5274 7776 5292 7794
rect 5274 7794 5292 7812
rect 5274 7812 5292 7830
rect 5274 7830 5292 7848
rect 5274 7848 5292 7866
rect 5274 7866 5292 7884
rect 5274 7884 5292 7902
rect 5274 7902 5292 7920
rect 5274 7920 5292 7938
rect 5274 7938 5292 7956
rect 5274 7956 5292 7974
rect 5274 7974 5292 7992
rect 5274 7992 5292 8010
rect 5274 8010 5292 8028
rect 5274 8028 5292 8046
rect 5274 8046 5292 8064
rect 5274 8064 5292 8082
rect 5274 8082 5292 8100
rect 5274 8100 5292 8118
rect 5274 8118 5292 8136
rect 5274 8136 5292 8154
rect 5274 8154 5292 8172
rect 5274 8172 5292 8190
rect 5274 8190 5292 8208
rect 5274 8208 5292 8226
rect 5274 8226 5292 8244
rect 5292 396 5310 414
rect 5292 414 5310 432
rect 5292 432 5310 450
rect 5292 450 5310 468
rect 5292 468 5310 486
rect 5292 486 5310 504
rect 5292 504 5310 522
rect 5292 522 5310 540
rect 5292 540 5310 558
rect 5292 558 5310 576
rect 5292 576 5310 594
rect 5292 594 5310 612
rect 5292 612 5310 630
rect 5292 630 5310 648
rect 5292 648 5310 666
rect 5292 666 5310 684
rect 5292 684 5310 702
rect 5292 702 5310 720
rect 5292 720 5310 738
rect 5292 738 5310 756
rect 5292 756 5310 774
rect 5292 774 5310 792
rect 5292 792 5310 810
rect 5292 810 5310 828
rect 5292 828 5310 846
rect 5292 972 5310 990
rect 5292 990 5310 1008
rect 5292 1008 5310 1026
rect 5292 1026 5310 1044
rect 5292 1044 5310 1062
rect 5292 1062 5310 1080
rect 5292 1080 5310 1098
rect 5292 1098 5310 1116
rect 5292 1116 5310 1134
rect 5292 1134 5310 1152
rect 5292 1152 5310 1170
rect 5292 1170 5310 1188
rect 5292 1188 5310 1206
rect 5292 1206 5310 1224
rect 5292 1224 5310 1242
rect 5292 1242 5310 1260
rect 5292 1260 5310 1278
rect 5292 1278 5310 1296
rect 5292 1296 5310 1314
rect 5292 1314 5310 1332
rect 5292 1332 5310 1350
rect 5292 1350 5310 1368
rect 5292 1368 5310 1386
rect 5292 1386 5310 1404
rect 5292 1404 5310 1422
rect 5292 1422 5310 1440
rect 5292 1440 5310 1458
rect 5292 1458 5310 1476
rect 5292 1476 5310 1494
rect 5292 1494 5310 1512
rect 5292 1512 5310 1530
rect 5292 1530 5310 1548
rect 5292 1548 5310 1566
rect 5292 1566 5310 1584
rect 5292 1584 5310 1602
rect 5292 1602 5310 1620
rect 5292 1620 5310 1638
rect 5292 1638 5310 1656
rect 5292 1656 5310 1674
rect 5292 1674 5310 1692
rect 5292 1692 5310 1710
rect 5292 1710 5310 1728
rect 5292 1728 5310 1746
rect 5292 1746 5310 1764
rect 5292 1764 5310 1782
rect 5292 1782 5310 1800
rect 5292 1800 5310 1818
rect 5292 1818 5310 1836
rect 5292 1836 5310 1854
rect 5292 1854 5310 1872
rect 5292 1872 5310 1890
rect 5292 1890 5310 1908
rect 5292 1908 5310 1926
rect 5292 1926 5310 1944
rect 5292 1944 5310 1962
rect 5292 1962 5310 1980
rect 5292 1980 5310 1998
rect 5292 1998 5310 2016
rect 5292 2016 5310 2034
rect 5292 2034 5310 2052
rect 5292 2052 5310 2070
rect 5292 2070 5310 2088
rect 5292 2088 5310 2106
rect 5292 2106 5310 2124
rect 5292 2124 5310 2142
rect 5292 2142 5310 2160
rect 5292 2160 5310 2178
rect 5292 2178 5310 2196
rect 5292 2196 5310 2214
rect 5292 2214 5310 2232
rect 5292 2232 5310 2250
rect 5292 2250 5310 2268
rect 5292 2268 5310 2286
rect 5292 2286 5310 2304
rect 5292 2304 5310 2322
rect 5292 2322 5310 2340
rect 5292 2340 5310 2358
rect 5292 2358 5310 2376
rect 5292 2376 5310 2394
rect 5292 2394 5310 2412
rect 5292 2610 5310 2628
rect 5292 2628 5310 2646
rect 5292 2646 5310 2664
rect 5292 2664 5310 2682
rect 5292 2682 5310 2700
rect 5292 2700 5310 2718
rect 5292 2718 5310 2736
rect 5292 2736 5310 2754
rect 5292 2754 5310 2772
rect 5292 2772 5310 2790
rect 5292 2790 5310 2808
rect 5292 2808 5310 2826
rect 5292 2826 5310 2844
rect 5292 2844 5310 2862
rect 5292 2862 5310 2880
rect 5292 2880 5310 2898
rect 5292 2898 5310 2916
rect 5292 2916 5310 2934
rect 5292 2934 5310 2952
rect 5292 2952 5310 2970
rect 5292 2970 5310 2988
rect 5292 2988 5310 3006
rect 5292 3006 5310 3024
rect 5292 3024 5310 3042
rect 5292 3042 5310 3060
rect 5292 3060 5310 3078
rect 5292 3078 5310 3096
rect 5292 3096 5310 3114
rect 5292 3114 5310 3132
rect 5292 3132 5310 3150
rect 5292 3150 5310 3168
rect 5292 3168 5310 3186
rect 5292 3186 5310 3204
rect 5292 3204 5310 3222
rect 5292 3222 5310 3240
rect 5292 3240 5310 3258
rect 5292 3258 5310 3276
rect 5292 3276 5310 3294
rect 5292 3294 5310 3312
rect 5292 3312 5310 3330
rect 5292 3330 5310 3348
rect 5292 3348 5310 3366
rect 5292 3366 5310 3384
rect 5292 3384 5310 3402
rect 5292 3402 5310 3420
rect 5292 3420 5310 3438
rect 5292 3438 5310 3456
rect 5292 3456 5310 3474
rect 5292 3474 5310 3492
rect 5292 3492 5310 3510
rect 5292 3510 5310 3528
rect 5292 3528 5310 3546
rect 5292 3546 5310 3564
rect 5292 3564 5310 3582
rect 5292 3582 5310 3600
rect 5292 3600 5310 3618
rect 5292 3618 5310 3636
rect 5292 3636 5310 3654
rect 5292 3654 5310 3672
rect 5292 3672 5310 3690
rect 5292 3690 5310 3708
rect 5292 3708 5310 3726
rect 5292 3726 5310 3744
rect 5292 3744 5310 3762
rect 5292 3762 5310 3780
rect 5292 3780 5310 3798
rect 5292 3798 5310 3816
rect 5292 3816 5310 3834
rect 5292 3834 5310 3852
rect 5292 3852 5310 3870
rect 5292 3870 5310 3888
rect 5292 3888 5310 3906
rect 5292 3906 5310 3924
rect 5292 3924 5310 3942
rect 5292 3942 5310 3960
rect 5292 3960 5310 3978
rect 5292 3978 5310 3996
rect 5292 3996 5310 4014
rect 5292 4014 5310 4032
rect 5292 4032 5310 4050
rect 5292 4050 5310 4068
rect 5292 4068 5310 4086
rect 5292 4086 5310 4104
rect 5292 4104 5310 4122
rect 5292 4122 5310 4140
rect 5292 4140 5310 4158
rect 5292 4158 5310 4176
rect 5292 4176 5310 4194
rect 5292 4194 5310 4212
rect 5292 4212 5310 4230
rect 5292 4230 5310 4248
rect 5292 4248 5310 4266
rect 5292 4266 5310 4284
rect 5292 4284 5310 4302
rect 5292 4302 5310 4320
rect 5292 4320 5310 4338
rect 5292 4338 5310 4356
rect 5292 4356 5310 4374
rect 5292 4374 5310 4392
rect 5292 4392 5310 4410
rect 5292 4410 5310 4428
rect 5292 4428 5310 4446
rect 5292 4446 5310 4464
rect 5292 4464 5310 4482
rect 5292 4482 5310 4500
rect 5292 4500 5310 4518
rect 5292 4518 5310 4536
rect 5292 4536 5310 4554
rect 5292 4554 5310 4572
rect 5292 4572 5310 4590
rect 5292 4590 5310 4608
rect 5292 4608 5310 4626
rect 5292 4626 5310 4644
rect 5292 4644 5310 4662
rect 5292 4662 5310 4680
rect 5292 4680 5310 4698
rect 5292 4914 5310 4932
rect 5292 4932 5310 4950
rect 5292 4950 5310 4968
rect 5292 4968 5310 4986
rect 5292 4986 5310 5004
rect 5292 5004 5310 5022
rect 5292 5022 5310 5040
rect 5292 5040 5310 5058
rect 5292 5058 5310 5076
rect 5292 5076 5310 5094
rect 5292 5094 5310 5112
rect 5292 5112 5310 5130
rect 5292 5130 5310 5148
rect 5292 5148 5310 5166
rect 5292 5166 5310 5184
rect 5292 5184 5310 5202
rect 5292 5202 5310 5220
rect 5292 5220 5310 5238
rect 5292 5238 5310 5256
rect 5292 5256 5310 5274
rect 5292 5274 5310 5292
rect 5292 5292 5310 5310
rect 5292 5310 5310 5328
rect 5292 5328 5310 5346
rect 5292 5346 5310 5364
rect 5292 5364 5310 5382
rect 5292 5382 5310 5400
rect 5292 5400 5310 5418
rect 5292 5418 5310 5436
rect 5292 5436 5310 5454
rect 5292 5454 5310 5472
rect 5292 5472 5310 5490
rect 5292 5490 5310 5508
rect 5292 5508 5310 5526
rect 5292 5526 5310 5544
rect 5292 5544 5310 5562
rect 5292 5562 5310 5580
rect 5292 5580 5310 5598
rect 5292 5598 5310 5616
rect 5292 5616 5310 5634
rect 5292 5634 5310 5652
rect 5292 5652 5310 5670
rect 5292 5670 5310 5688
rect 5292 5688 5310 5706
rect 5292 5706 5310 5724
rect 5292 5724 5310 5742
rect 5292 5742 5310 5760
rect 5292 5760 5310 5778
rect 5292 5778 5310 5796
rect 5292 5796 5310 5814
rect 5292 5814 5310 5832
rect 5292 5832 5310 5850
rect 5292 5850 5310 5868
rect 5292 5868 5310 5886
rect 5292 5886 5310 5904
rect 5292 5904 5310 5922
rect 5292 5922 5310 5940
rect 5292 5940 5310 5958
rect 5292 5958 5310 5976
rect 5292 5976 5310 5994
rect 5292 5994 5310 6012
rect 5292 6012 5310 6030
rect 5292 6030 5310 6048
rect 5292 6048 5310 6066
rect 5292 6066 5310 6084
rect 5292 6084 5310 6102
rect 5292 6102 5310 6120
rect 5292 6120 5310 6138
rect 5292 6138 5310 6156
rect 5292 6156 5310 6174
rect 5292 6174 5310 6192
rect 5292 6192 5310 6210
rect 5292 6210 5310 6228
rect 5292 6228 5310 6246
rect 5292 6246 5310 6264
rect 5292 6264 5310 6282
rect 5292 6282 5310 6300
rect 5292 6300 5310 6318
rect 5292 6318 5310 6336
rect 5292 6336 5310 6354
rect 5292 6354 5310 6372
rect 5292 6372 5310 6390
rect 5292 6390 5310 6408
rect 5292 6408 5310 6426
rect 5292 6426 5310 6444
rect 5292 6444 5310 6462
rect 5292 6462 5310 6480
rect 5292 6480 5310 6498
rect 5292 6498 5310 6516
rect 5292 6516 5310 6534
rect 5292 6534 5310 6552
rect 5292 6552 5310 6570
rect 5292 6570 5310 6588
rect 5292 6588 5310 6606
rect 5292 6606 5310 6624
rect 5292 6624 5310 6642
rect 5292 6642 5310 6660
rect 5292 6660 5310 6678
rect 5292 6678 5310 6696
rect 5292 6696 5310 6714
rect 5292 6714 5310 6732
rect 5292 6732 5310 6750
rect 5292 6750 5310 6768
rect 5292 6768 5310 6786
rect 5292 6786 5310 6804
rect 5292 6804 5310 6822
rect 5292 6822 5310 6840
rect 5292 6840 5310 6858
rect 5292 6858 5310 6876
rect 5292 6876 5310 6894
rect 5292 6894 5310 6912
rect 5292 6912 5310 6930
rect 5292 6930 5310 6948
rect 5292 6948 5310 6966
rect 5292 6966 5310 6984
rect 5292 6984 5310 7002
rect 5292 7002 5310 7020
rect 5292 7020 5310 7038
rect 5292 7038 5310 7056
rect 5292 7056 5310 7074
rect 5292 7074 5310 7092
rect 5292 7092 5310 7110
rect 5292 7110 5310 7128
rect 5292 7128 5310 7146
rect 5292 7146 5310 7164
rect 5292 7164 5310 7182
rect 5292 7182 5310 7200
rect 5292 7200 5310 7218
rect 5292 7218 5310 7236
rect 5292 7236 5310 7254
rect 5292 7254 5310 7272
rect 5292 7272 5310 7290
rect 5292 7290 5310 7308
rect 5292 7308 5310 7326
rect 5292 7326 5310 7344
rect 5292 7344 5310 7362
rect 5292 7362 5310 7380
rect 5292 7380 5310 7398
rect 5292 7398 5310 7416
rect 5292 7416 5310 7434
rect 5292 7434 5310 7452
rect 5292 7452 5310 7470
rect 5292 7470 5310 7488
rect 5292 7488 5310 7506
rect 5292 7506 5310 7524
rect 5292 7524 5310 7542
rect 5292 7542 5310 7560
rect 5292 7560 5310 7578
rect 5292 7578 5310 7596
rect 5292 7596 5310 7614
rect 5292 7614 5310 7632
rect 5292 7632 5310 7650
rect 5292 7650 5310 7668
rect 5292 7668 5310 7686
rect 5292 7686 5310 7704
rect 5292 7704 5310 7722
rect 5292 7722 5310 7740
rect 5292 7740 5310 7758
rect 5292 7758 5310 7776
rect 5292 7776 5310 7794
rect 5292 7794 5310 7812
rect 5292 7812 5310 7830
rect 5292 7830 5310 7848
rect 5292 7848 5310 7866
rect 5292 7866 5310 7884
rect 5292 7884 5310 7902
rect 5292 7902 5310 7920
rect 5292 7920 5310 7938
rect 5292 7938 5310 7956
rect 5292 7956 5310 7974
rect 5292 7974 5310 7992
rect 5292 7992 5310 8010
rect 5292 8010 5310 8028
rect 5292 8028 5310 8046
rect 5292 8046 5310 8064
rect 5292 8064 5310 8082
rect 5292 8082 5310 8100
rect 5292 8100 5310 8118
rect 5292 8118 5310 8136
rect 5292 8136 5310 8154
rect 5292 8154 5310 8172
rect 5292 8172 5310 8190
rect 5292 8190 5310 8208
rect 5292 8208 5310 8226
rect 5292 8226 5310 8244
rect 5292 8244 5310 8262
rect 5292 8262 5310 8280
rect 5310 414 5328 432
rect 5310 432 5328 450
rect 5310 450 5328 468
rect 5310 468 5328 486
rect 5310 486 5328 504
rect 5310 504 5328 522
rect 5310 522 5328 540
rect 5310 540 5328 558
rect 5310 558 5328 576
rect 5310 576 5328 594
rect 5310 594 5328 612
rect 5310 612 5328 630
rect 5310 630 5328 648
rect 5310 648 5328 666
rect 5310 666 5328 684
rect 5310 684 5328 702
rect 5310 702 5328 720
rect 5310 720 5328 738
rect 5310 738 5328 756
rect 5310 756 5328 774
rect 5310 774 5328 792
rect 5310 792 5328 810
rect 5310 810 5328 828
rect 5310 828 5328 846
rect 5310 990 5328 1008
rect 5310 1008 5328 1026
rect 5310 1026 5328 1044
rect 5310 1044 5328 1062
rect 5310 1062 5328 1080
rect 5310 1080 5328 1098
rect 5310 1098 5328 1116
rect 5310 1116 5328 1134
rect 5310 1134 5328 1152
rect 5310 1152 5328 1170
rect 5310 1170 5328 1188
rect 5310 1188 5328 1206
rect 5310 1206 5328 1224
rect 5310 1224 5328 1242
rect 5310 1242 5328 1260
rect 5310 1260 5328 1278
rect 5310 1278 5328 1296
rect 5310 1296 5328 1314
rect 5310 1314 5328 1332
rect 5310 1332 5328 1350
rect 5310 1350 5328 1368
rect 5310 1368 5328 1386
rect 5310 1386 5328 1404
rect 5310 1404 5328 1422
rect 5310 1422 5328 1440
rect 5310 1440 5328 1458
rect 5310 1458 5328 1476
rect 5310 1476 5328 1494
rect 5310 1494 5328 1512
rect 5310 1512 5328 1530
rect 5310 1530 5328 1548
rect 5310 1548 5328 1566
rect 5310 1566 5328 1584
rect 5310 1584 5328 1602
rect 5310 1602 5328 1620
rect 5310 1620 5328 1638
rect 5310 1638 5328 1656
rect 5310 1656 5328 1674
rect 5310 1674 5328 1692
rect 5310 1692 5328 1710
rect 5310 1710 5328 1728
rect 5310 1728 5328 1746
rect 5310 1746 5328 1764
rect 5310 1764 5328 1782
rect 5310 1782 5328 1800
rect 5310 1800 5328 1818
rect 5310 1818 5328 1836
rect 5310 1836 5328 1854
rect 5310 1854 5328 1872
rect 5310 1872 5328 1890
rect 5310 1890 5328 1908
rect 5310 1908 5328 1926
rect 5310 1926 5328 1944
rect 5310 1944 5328 1962
rect 5310 1962 5328 1980
rect 5310 1980 5328 1998
rect 5310 1998 5328 2016
rect 5310 2016 5328 2034
rect 5310 2034 5328 2052
rect 5310 2052 5328 2070
rect 5310 2070 5328 2088
rect 5310 2088 5328 2106
rect 5310 2106 5328 2124
rect 5310 2124 5328 2142
rect 5310 2142 5328 2160
rect 5310 2160 5328 2178
rect 5310 2178 5328 2196
rect 5310 2196 5328 2214
rect 5310 2214 5328 2232
rect 5310 2232 5328 2250
rect 5310 2250 5328 2268
rect 5310 2268 5328 2286
rect 5310 2286 5328 2304
rect 5310 2304 5328 2322
rect 5310 2322 5328 2340
rect 5310 2340 5328 2358
rect 5310 2358 5328 2376
rect 5310 2376 5328 2394
rect 5310 2394 5328 2412
rect 5310 2628 5328 2646
rect 5310 2646 5328 2664
rect 5310 2664 5328 2682
rect 5310 2682 5328 2700
rect 5310 2700 5328 2718
rect 5310 2718 5328 2736
rect 5310 2736 5328 2754
rect 5310 2754 5328 2772
rect 5310 2772 5328 2790
rect 5310 2790 5328 2808
rect 5310 2808 5328 2826
rect 5310 2826 5328 2844
rect 5310 2844 5328 2862
rect 5310 2862 5328 2880
rect 5310 2880 5328 2898
rect 5310 2898 5328 2916
rect 5310 2916 5328 2934
rect 5310 2934 5328 2952
rect 5310 2952 5328 2970
rect 5310 2970 5328 2988
rect 5310 2988 5328 3006
rect 5310 3006 5328 3024
rect 5310 3024 5328 3042
rect 5310 3042 5328 3060
rect 5310 3060 5328 3078
rect 5310 3078 5328 3096
rect 5310 3096 5328 3114
rect 5310 3114 5328 3132
rect 5310 3132 5328 3150
rect 5310 3150 5328 3168
rect 5310 3168 5328 3186
rect 5310 3186 5328 3204
rect 5310 3204 5328 3222
rect 5310 3222 5328 3240
rect 5310 3240 5328 3258
rect 5310 3258 5328 3276
rect 5310 3276 5328 3294
rect 5310 3294 5328 3312
rect 5310 3312 5328 3330
rect 5310 3330 5328 3348
rect 5310 3348 5328 3366
rect 5310 3366 5328 3384
rect 5310 3384 5328 3402
rect 5310 3402 5328 3420
rect 5310 3420 5328 3438
rect 5310 3438 5328 3456
rect 5310 3456 5328 3474
rect 5310 3474 5328 3492
rect 5310 3492 5328 3510
rect 5310 3510 5328 3528
rect 5310 3528 5328 3546
rect 5310 3546 5328 3564
rect 5310 3564 5328 3582
rect 5310 3582 5328 3600
rect 5310 3600 5328 3618
rect 5310 3618 5328 3636
rect 5310 3636 5328 3654
rect 5310 3654 5328 3672
rect 5310 3672 5328 3690
rect 5310 3690 5328 3708
rect 5310 3708 5328 3726
rect 5310 3726 5328 3744
rect 5310 3744 5328 3762
rect 5310 3762 5328 3780
rect 5310 3780 5328 3798
rect 5310 3798 5328 3816
rect 5310 3816 5328 3834
rect 5310 3834 5328 3852
rect 5310 3852 5328 3870
rect 5310 3870 5328 3888
rect 5310 3888 5328 3906
rect 5310 3906 5328 3924
rect 5310 3924 5328 3942
rect 5310 3942 5328 3960
rect 5310 3960 5328 3978
rect 5310 3978 5328 3996
rect 5310 3996 5328 4014
rect 5310 4014 5328 4032
rect 5310 4032 5328 4050
rect 5310 4050 5328 4068
rect 5310 4068 5328 4086
rect 5310 4086 5328 4104
rect 5310 4104 5328 4122
rect 5310 4122 5328 4140
rect 5310 4140 5328 4158
rect 5310 4158 5328 4176
rect 5310 4176 5328 4194
rect 5310 4194 5328 4212
rect 5310 4212 5328 4230
rect 5310 4230 5328 4248
rect 5310 4248 5328 4266
rect 5310 4266 5328 4284
rect 5310 4284 5328 4302
rect 5310 4302 5328 4320
rect 5310 4320 5328 4338
rect 5310 4338 5328 4356
rect 5310 4356 5328 4374
rect 5310 4374 5328 4392
rect 5310 4392 5328 4410
rect 5310 4410 5328 4428
rect 5310 4428 5328 4446
rect 5310 4446 5328 4464
rect 5310 4464 5328 4482
rect 5310 4482 5328 4500
rect 5310 4500 5328 4518
rect 5310 4518 5328 4536
rect 5310 4536 5328 4554
rect 5310 4554 5328 4572
rect 5310 4572 5328 4590
rect 5310 4590 5328 4608
rect 5310 4608 5328 4626
rect 5310 4626 5328 4644
rect 5310 4644 5328 4662
rect 5310 4662 5328 4680
rect 5310 4680 5328 4698
rect 5310 4698 5328 4716
rect 5310 4932 5328 4950
rect 5310 4950 5328 4968
rect 5310 4968 5328 4986
rect 5310 4986 5328 5004
rect 5310 5004 5328 5022
rect 5310 5022 5328 5040
rect 5310 5040 5328 5058
rect 5310 5058 5328 5076
rect 5310 5076 5328 5094
rect 5310 5094 5328 5112
rect 5310 5112 5328 5130
rect 5310 5130 5328 5148
rect 5310 5148 5328 5166
rect 5310 5166 5328 5184
rect 5310 5184 5328 5202
rect 5310 5202 5328 5220
rect 5310 5220 5328 5238
rect 5310 5238 5328 5256
rect 5310 5256 5328 5274
rect 5310 5274 5328 5292
rect 5310 5292 5328 5310
rect 5310 5310 5328 5328
rect 5310 5328 5328 5346
rect 5310 5346 5328 5364
rect 5310 5364 5328 5382
rect 5310 5382 5328 5400
rect 5310 5400 5328 5418
rect 5310 5418 5328 5436
rect 5310 5436 5328 5454
rect 5310 5454 5328 5472
rect 5310 5472 5328 5490
rect 5310 5490 5328 5508
rect 5310 5508 5328 5526
rect 5310 5526 5328 5544
rect 5310 5544 5328 5562
rect 5310 5562 5328 5580
rect 5310 5580 5328 5598
rect 5310 5598 5328 5616
rect 5310 5616 5328 5634
rect 5310 5634 5328 5652
rect 5310 5652 5328 5670
rect 5310 5670 5328 5688
rect 5310 5688 5328 5706
rect 5310 5706 5328 5724
rect 5310 5724 5328 5742
rect 5310 5742 5328 5760
rect 5310 5760 5328 5778
rect 5310 5778 5328 5796
rect 5310 5796 5328 5814
rect 5310 5814 5328 5832
rect 5310 5832 5328 5850
rect 5310 5850 5328 5868
rect 5310 5868 5328 5886
rect 5310 5886 5328 5904
rect 5310 5904 5328 5922
rect 5310 5922 5328 5940
rect 5310 5940 5328 5958
rect 5310 5958 5328 5976
rect 5310 5976 5328 5994
rect 5310 5994 5328 6012
rect 5310 6012 5328 6030
rect 5310 6030 5328 6048
rect 5310 6048 5328 6066
rect 5310 6066 5328 6084
rect 5310 6084 5328 6102
rect 5310 6102 5328 6120
rect 5310 6120 5328 6138
rect 5310 6138 5328 6156
rect 5310 6156 5328 6174
rect 5310 6174 5328 6192
rect 5310 6192 5328 6210
rect 5310 6210 5328 6228
rect 5310 6228 5328 6246
rect 5310 6246 5328 6264
rect 5310 6264 5328 6282
rect 5310 6282 5328 6300
rect 5310 6300 5328 6318
rect 5310 6318 5328 6336
rect 5310 6336 5328 6354
rect 5310 6354 5328 6372
rect 5310 6372 5328 6390
rect 5310 6390 5328 6408
rect 5310 6408 5328 6426
rect 5310 6426 5328 6444
rect 5310 6444 5328 6462
rect 5310 6462 5328 6480
rect 5310 6480 5328 6498
rect 5310 6498 5328 6516
rect 5310 6516 5328 6534
rect 5310 6534 5328 6552
rect 5310 6552 5328 6570
rect 5310 6570 5328 6588
rect 5310 6588 5328 6606
rect 5310 6606 5328 6624
rect 5310 6624 5328 6642
rect 5310 6642 5328 6660
rect 5310 6660 5328 6678
rect 5310 6678 5328 6696
rect 5310 6696 5328 6714
rect 5310 6714 5328 6732
rect 5310 6732 5328 6750
rect 5310 6750 5328 6768
rect 5310 6768 5328 6786
rect 5310 6786 5328 6804
rect 5310 6804 5328 6822
rect 5310 6822 5328 6840
rect 5310 6840 5328 6858
rect 5310 6858 5328 6876
rect 5310 6876 5328 6894
rect 5310 6894 5328 6912
rect 5310 6912 5328 6930
rect 5310 6930 5328 6948
rect 5310 6948 5328 6966
rect 5310 6966 5328 6984
rect 5310 6984 5328 7002
rect 5310 7002 5328 7020
rect 5310 7020 5328 7038
rect 5310 7038 5328 7056
rect 5310 7056 5328 7074
rect 5310 7074 5328 7092
rect 5310 7092 5328 7110
rect 5310 7110 5328 7128
rect 5310 7128 5328 7146
rect 5310 7146 5328 7164
rect 5310 7164 5328 7182
rect 5310 7182 5328 7200
rect 5310 7200 5328 7218
rect 5310 7218 5328 7236
rect 5310 7236 5328 7254
rect 5310 7254 5328 7272
rect 5310 7272 5328 7290
rect 5310 7290 5328 7308
rect 5310 7308 5328 7326
rect 5310 7326 5328 7344
rect 5310 7344 5328 7362
rect 5310 7362 5328 7380
rect 5310 7380 5328 7398
rect 5310 7398 5328 7416
rect 5310 7416 5328 7434
rect 5310 7434 5328 7452
rect 5310 7452 5328 7470
rect 5310 7470 5328 7488
rect 5310 7488 5328 7506
rect 5310 7506 5328 7524
rect 5310 7524 5328 7542
rect 5310 7542 5328 7560
rect 5310 7560 5328 7578
rect 5310 7578 5328 7596
rect 5310 7596 5328 7614
rect 5310 7614 5328 7632
rect 5310 7632 5328 7650
rect 5310 7650 5328 7668
rect 5310 7668 5328 7686
rect 5310 7686 5328 7704
rect 5310 7704 5328 7722
rect 5310 7722 5328 7740
rect 5310 7740 5328 7758
rect 5310 7758 5328 7776
rect 5310 7776 5328 7794
rect 5310 7794 5328 7812
rect 5310 7812 5328 7830
rect 5310 7830 5328 7848
rect 5310 7848 5328 7866
rect 5310 7866 5328 7884
rect 5310 7884 5328 7902
rect 5310 7902 5328 7920
rect 5310 7920 5328 7938
rect 5310 7938 5328 7956
rect 5310 7956 5328 7974
rect 5310 7974 5328 7992
rect 5310 7992 5328 8010
rect 5310 8010 5328 8028
rect 5310 8028 5328 8046
rect 5310 8046 5328 8064
rect 5310 8064 5328 8082
rect 5310 8082 5328 8100
rect 5310 8100 5328 8118
rect 5310 8118 5328 8136
rect 5310 8136 5328 8154
rect 5310 8154 5328 8172
rect 5310 8172 5328 8190
rect 5310 8190 5328 8208
rect 5310 8208 5328 8226
rect 5310 8226 5328 8244
rect 5310 8244 5328 8262
rect 5310 8262 5328 8280
rect 5310 8280 5328 8298
rect 5328 414 5346 432
rect 5328 432 5346 450
rect 5328 450 5346 468
rect 5328 468 5346 486
rect 5328 486 5346 504
rect 5328 504 5346 522
rect 5328 522 5346 540
rect 5328 540 5346 558
rect 5328 558 5346 576
rect 5328 576 5346 594
rect 5328 594 5346 612
rect 5328 612 5346 630
rect 5328 630 5346 648
rect 5328 648 5346 666
rect 5328 666 5346 684
rect 5328 684 5346 702
rect 5328 702 5346 720
rect 5328 720 5346 738
rect 5328 738 5346 756
rect 5328 756 5346 774
rect 5328 774 5346 792
rect 5328 792 5346 810
rect 5328 810 5346 828
rect 5328 828 5346 846
rect 5328 846 5346 864
rect 5328 990 5346 1008
rect 5328 1008 5346 1026
rect 5328 1026 5346 1044
rect 5328 1044 5346 1062
rect 5328 1062 5346 1080
rect 5328 1080 5346 1098
rect 5328 1098 5346 1116
rect 5328 1116 5346 1134
rect 5328 1134 5346 1152
rect 5328 1152 5346 1170
rect 5328 1170 5346 1188
rect 5328 1188 5346 1206
rect 5328 1206 5346 1224
rect 5328 1224 5346 1242
rect 5328 1242 5346 1260
rect 5328 1260 5346 1278
rect 5328 1278 5346 1296
rect 5328 1296 5346 1314
rect 5328 1314 5346 1332
rect 5328 1332 5346 1350
rect 5328 1350 5346 1368
rect 5328 1368 5346 1386
rect 5328 1386 5346 1404
rect 5328 1404 5346 1422
rect 5328 1422 5346 1440
rect 5328 1440 5346 1458
rect 5328 1458 5346 1476
rect 5328 1476 5346 1494
rect 5328 1494 5346 1512
rect 5328 1512 5346 1530
rect 5328 1530 5346 1548
rect 5328 1548 5346 1566
rect 5328 1566 5346 1584
rect 5328 1584 5346 1602
rect 5328 1602 5346 1620
rect 5328 1620 5346 1638
rect 5328 1638 5346 1656
rect 5328 1656 5346 1674
rect 5328 1674 5346 1692
rect 5328 1692 5346 1710
rect 5328 1710 5346 1728
rect 5328 1728 5346 1746
rect 5328 1746 5346 1764
rect 5328 1764 5346 1782
rect 5328 1782 5346 1800
rect 5328 1800 5346 1818
rect 5328 1818 5346 1836
rect 5328 1836 5346 1854
rect 5328 1854 5346 1872
rect 5328 1872 5346 1890
rect 5328 1890 5346 1908
rect 5328 1908 5346 1926
rect 5328 1926 5346 1944
rect 5328 1944 5346 1962
rect 5328 1962 5346 1980
rect 5328 1980 5346 1998
rect 5328 1998 5346 2016
rect 5328 2016 5346 2034
rect 5328 2034 5346 2052
rect 5328 2052 5346 2070
rect 5328 2070 5346 2088
rect 5328 2088 5346 2106
rect 5328 2106 5346 2124
rect 5328 2124 5346 2142
rect 5328 2142 5346 2160
rect 5328 2160 5346 2178
rect 5328 2178 5346 2196
rect 5328 2196 5346 2214
rect 5328 2214 5346 2232
rect 5328 2232 5346 2250
rect 5328 2250 5346 2268
rect 5328 2268 5346 2286
rect 5328 2286 5346 2304
rect 5328 2304 5346 2322
rect 5328 2322 5346 2340
rect 5328 2340 5346 2358
rect 5328 2358 5346 2376
rect 5328 2376 5346 2394
rect 5328 2394 5346 2412
rect 5328 2412 5346 2430
rect 5328 2628 5346 2646
rect 5328 2646 5346 2664
rect 5328 2664 5346 2682
rect 5328 2682 5346 2700
rect 5328 2700 5346 2718
rect 5328 2718 5346 2736
rect 5328 2736 5346 2754
rect 5328 2754 5346 2772
rect 5328 2772 5346 2790
rect 5328 2790 5346 2808
rect 5328 2808 5346 2826
rect 5328 2826 5346 2844
rect 5328 2844 5346 2862
rect 5328 2862 5346 2880
rect 5328 2880 5346 2898
rect 5328 2898 5346 2916
rect 5328 2916 5346 2934
rect 5328 2934 5346 2952
rect 5328 2952 5346 2970
rect 5328 2970 5346 2988
rect 5328 2988 5346 3006
rect 5328 3006 5346 3024
rect 5328 3024 5346 3042
rect 5328 3042 5346 3060
rect 5328 3060 5346 3078
rect 5328 3078 5346 3096
rect 5328 3096 5346 3114
rect 5328 3114 5346 3132
rect 5328 3132 5346 3150
rect 5328 3150 5346 3168
rect 5328 3168 5346 3186
rect 5328 3186 5346 3204
rect 5328 3204 5346 3222
rect 5328 3222 5346 3240
rect 5328 3240 5346 3258
rect 5328 3258 5346 3276
rect 5328 3276 5346 3294
rect 5328 3294 5346 3312
rect 5328 3312 5346 3330
rect 5328 3330 5346 3348
rect 5328 3348 5346 3366
rect 5328 3366 5346 3384
rect 5328 3384 5346 3402
rect 5328 3402 5346 3420
rect 5328 3420 5346 3438
rect 5328 3438 5346 3456
rect 5328 3456 5346 3474
rect 5328 3474 5346 3492
rect 5328 3492 5346 3510
rect 5328 3510 5346 3528
rect 5328 3528 5346 3546
rect 5328 3546 5346 3564
rect 5328 3564 5346 3582
rect 5328 3582 5346 3600
rect 5328 3600 5346 3618
rect 5328 3618 5346 3636
rect 5328 3636 5346 3654
rect 5328 3654 5346 3672
rect 5328 3672 5346 3690
rect 5328 3690 5346 3708
rect 5328 3708 5346 3726
rect 5328 3726 5346 3744
rect 5328 3744 5346 3762
rect 5328 3762 5346 3780
rect 5328 3780 5346 3798
rect 5328 3798 5346 3816
rect 5328 3816 5346 3834
rect 5328 3834 5346 3852
rect 5328 3852 5346 3870
rect 5328 3870 5346 3888
rect 5328 3888 5346 3906
rect 5328 3906 5346 3924
rect 5328 3924 5346 3942
rect 5328 3942 5346 3960
rect 5328 3960 5346 3978
rect 5328 3978 5346 3996
rect 5328 3996 5346 4014
rect 5328 4014 5346 4032
rect 5328 4032 5346 4050
rect 5328 4050 5346 4068
rect 5328 4068 5346 4086
rect 5328 4086 5346 4104
rect 5328 4104 5346 4122
rect 5328 4122 5346 4140
rect 5328 4140 5346 4158
rect 5328 4158 5346 4176
rect 5328 4176 5346 4194
rect 5328 4194 5346 4212
rect 5328 4212 5346 4230
rect 5328 4230 5346 4248
rect 5328 4248 5346 4266
rect 5328 4266 5346 4284
rect 5328 4284 5346 4302
rect 5328 4302 5346 4320
rect 5328 4320 5346 4338
rect 5328 4338 5346 4356
rect 5328 4356 5346 4374
rect 5328 4374 5346 4392
rect 5328 4392 5346 4410
rect 5328 4410 5346 4428
rect 5328 4428 5346 4446
rect 5328 4446 5346 4464
rect 5328 4464 5346 4482
rect 5328 4482 5346 4500
rect 5328 4500 5346 4518
rect 5328 4518 5346 4536
rect 5328 4536 5346 4554
rect 5328 4554 5346 4572
rect 5328 4572 5346 4590
rect 5328 4590 5346 4608
rect 5328 4608 5346 4626
rect 5328 4626 5346 4644
rect 5328 4644 5346 4662
rect 5328 4662 5346 4680
rect 5328 4680 5346 4698
rect 5328 4698 5346 4716
rect 5328 4716 5346 4734
rect 5328 4950 5346 4968
rect 5328 4968 5346 4986
rect 5328 4986 5346 5004
rect 5328 5004 5346 5022
rect 5328 5022 5346 5040
rect 5328 5040 5346 5058
rect 5328 5058 5346 5076
rect 5328 5076 5346 5094
rect 5328 5094 5346 5112
rect 5328 5112 5346 5130
rect 5328 5130 5346 5148
rect 5328 5148 5346 5166
rect 5328 5166 5346 5184
rect 5328 5184 5346 5202
rect 5328 5202 5346 5220
rect 5328 5220 5346 5238
rect 5328 5238 5346 5256
rect 5328 5256 5346 5274
rect 5328 5274 5346 5292
rect 5328 5292 5346 5310
rect 5328 5310 5346 5328
rect 5328 5328 5346 5346
rect 5328 5346 5346 5364
rect 5328 5364 5346 5382
rect 5328 5382 5346 5400
rect 5328 5400 5346 5418
rect 5328 5418 5346 5436
rect 5328 5436 5346 5454
rect 5328 5454 5346 5472
rect 5328 5472 5346 5490
rect 5328 5490 5346 5508
rect 5328 5508 5346 5526
rect 5328 5526 5346 5544
rect 5328 5544 5346 5562
rect 5328 5562 5346 5580
rect 5328 5580 5346 5598
rect 5328 5598 5346 5616
rect 5328 5616 5346 5634
rect 5328 5634 5346 5652
rect 5328 5652 5346 5670
rect 5328 5670 5346 5688
rect 5328 5688 5346 5706
rect 5328 5706 5346 5724
rect 5328 5724 5346 5742
rect 5328 5742 5346 5760
rect 5328 5760 5346 5778
rect 5328 5778 5346 5796
rect 5328 5796 5346 5814
rect 5328 5814 5346 5832
rect 5328 5832 5346 5850
rect 5328 5850 5346 5868
rect 5328 5868 5346 5886
rect 5328 5886 5346 5904
rect 5328 5904 5346 5922
rect 5328 5922 5346 5940
rect 5328 5940 5346 5958
rect 5328 5958 5346 5976
rect 5328 5976 5346 5994
rect 5328 5994 5346 6012
rect 5328 6012 5346 6030
rect 5328 6030 5346 6048
rect 5328 6048 5346 6066
rect 5328 6066 5346 6084
rect 5328 6084 5346 6102
rect 5328 6102 5346 6120
rect 5328 6120 5346 6138
rect 5328 6138 5346 6156
rect 5328 6156 5346 6174
rect 5328 6174 5346 6192
rect 5328 6192 5346 6210
rect 5328 6210 5346 6228
rect 5328 6228 5346 6246
rect 5328 6246 5346 6264
rect 5328 6264 5346 6282
rect 5328 6282 5346 6300
rect 5328 6300 5346 6318
rect 5328 6318 5346 6336
rect 5328 6336 5346 6354
rect 5328 6354 5346 6372
rect 5328 6372 5346 6390
rect 5328 6390 5346 6408
rect 5328 6408 5346 6426
rect 5328 6426 5346 6444
rect 5328 6444 5346 6462
rect 5328 6462 5346 6480
rect 5328 6480 5346 6498
rect 5328 6498 5346 6516
rect 5328 6516 5346 6534
rect 5328 6534 5346 6552
rect 5328 6552 5346 6570
rect 5328 6570 5346 6588
rect 5328 6588 5346 6606
rect 5328 6606 5346 6624
rect 5328 6624 5346 6642
rect 5328 6642 5346 6660
rect 5328 6660 5346 6678
rect 5328 6678 5346 6696
rect 5328 6696 5346 6714
rect 5328 6714 5346 6732
rect 5328 6732 5346 6750
rect 5328 6750 5346 6768
rect 5328 6768 5346 6786
rect 5328 6786 5346 6804
rect 5328 6804 5346 6822
rect 5328 6822 5346 6840
rect 5328 6840 5346 6858
rect 5328 6858 5346 6876
rect 5328 6876 5346 6894
rect 5328 6894 5346 6912
rect 5328 6912 5346 6930
rect 5328 6930 5346 6948
rect 5328 6948 5346 6966
rect 5328 6966 5346 6984
rect 5328 6984 5346 7002
rect 5328 7002 5346 7020
rect 5328 7020 5346 7038
rect 5328 7038 5346 7056
rect 5328 7056 5346 7074
rect 5328 7074 5346 7092
rect 5328 7092 5346 7110
rect 5328 7110 5346 7128
rect 5328 7128 5346 7146
rect 5328 7146 5346 7164
rect 5328 7164 5346 7182
rect 5328 7182 5346 7200
rect 5328 7200 5346 7218
rect 5328 7218 5346 7236
rect 5328 7236 5346 7254
rect 5328 7254 5346 7272
rect 5328 7272 5346 7290
rect 5328 7290 5346 7308
rect 5328 7308 5346 7326
rect 5328 7326 5346 7344
rect 5328 7344 5346 7362
rect 5328 7362 5346 7380
rect 5328 7380 5346 7398
rect 5328 7398 5346 7416
rect 5328 7416 5346 7434
rect 5328 7434 5346 7452
rect 5328 7452 5346 7470
rect 5328 7470 5346 7488
rect 5328 7488 5346 7506
rect 5328 7506 5346 7524
rect 5328 7524 5346 7542
rect 5328 7542 5346 7560
rect 5328 7560 5346 7578
rect 5328 7578 5346 7596
rect 5328 7596 5346 7614
rect 5328 7614 5346 7632
rect 5328 7632 5346 7650
rect 5328 7650 5346 7668
rect 5328 7668 5346 7686
rect 5328 7686 5346 7704
rect 5328 7704 5346 7722
rect 5328 7722 5346 7740
rect 5328 7740 5346 7758
rect 5328 7758 5346 7776
rect 5328 7776 5346 7794
rect 5328 7794 5346 7812
rect 5328 7812 5346 7830
rect 5328 7830 5346 7848
rect 5328 7848 5346 7866
rect 5328 7866 5346 7884
rect 5328 7884 5346 7902
rect 5328 7902 5346 7920
rect 5328 7920 5346 7938
rect 5328 7938 5346 7956
rect 5328 7956 5346 7974
rect 5328 7974 5346 7992
rect 5328 7992 5346 8010
rect 5328 8010 5346 8028
rect 5328 8028 5346 8046
rect 5328 8046 5346 8064
rect 5328 8064 5346 8082
rect 5328 8082 5346 8100
rect 5328 8100 5346 8118
rect 5328 8118 5346 8136
rect 5328 8136 5346 8154
rect 5328 8154 5346 8172
rect 5328 8172 5346 8190
rect 5328 8190 5346 8208
rect 5328 8208 5346 8226
rect 5328 8226 5346 8244
rect 5328 8244 5346 8262
rect 5328 8262 5346 8280
rect 5328 8280 5346 8298
rect 5328 8298 5346 8316
rect 5346 432 5364 450
rect 5346 450 5364 468
rect 5346 468 5364 486
rect 5346 486 5364 504
rect 5346 504 5364 522
rect 5346 522 5364 540
rect 5346 540 5364 558
rect 5346 558 5364 576
rect 5346 576 5364 594
rect 5346 594 5364 612
rect 5346 612 5364 630
rect 5346 630 5364 648
rect 5346 648 5364 666
rect 5346 666 5364 684
rect 5346 684 5364 702
rect 5346 702 5364 720
rect 5346 720 5364 738
rect 5346 738 5364 756
rect 5346 756 5364 774
rect 5346 774 5364 792
rect 5346 792 5364 810
rect 5346 810 5364 828
rect 5346 828 5364 846
rect 5346 846 5364 864
rect 5346 990 5364 1008
rect 5346 1008 5364 1026
rect 5346 1026 5364 1044
rect 5346 1044 5364 1062
rect 5346 1062 5364 1080
rect 5346 1080 5364 1098
rect 5346 1098 5364 1116
rect 5346 1116 5364 1134
rect 5346 1134 5364 1152
rect 5346 1152 5364 1170
rect 5346 1170 5364 1188
rect 5346 1188 5364 1206
rect 5346 1206 5364 1224
rect 5346 1224 5364 1242
rect 5346 1242 5364 1260
rect 5346 1260 5364 1278
rect 5346 1278 5364 1296
rect 5346 1296 5364 1314
rect 5346 1314 5364 1332
rect 5346 1332 5364 1350
rect 5346 1350 5364 1368
rect 5346 1368 5364 1386
rect 5346 1386 5364 1404
rect 5346 1404 5364 1422
rect 5346 1422 5364 1440
rect 5346 1440 5364 1458
rect 5346 1458 5364 1476
rect 5346 1476 5364 1494
rect 5346 1494 5364 1512
rect 5346 1512 5364 1530
rect 5346 1530 5364 1548
rect 5346 1548 5364 1566
rect 5346 1566 5364 1584
rect 5346 1584 5364 1602
rect 5346 1602 5364 1620
rect 5346 1620 5364 1638
rect 5346 1638 5364 1656
rect 5346 1656 5364 1674
rect 5346 1674 5364 1692
rect 5346 1692 5364 1710
rect 5346 1710 5364 1728
rect 5346 1728 5364 1746
rect 5346 1746 5364 1764
rect 5346 1764 5364 1782
rect 5346 1782 5364 1800
rect 5346 1800 5364 1818
rect 5346 1818 5364 1836
rect 5346 1836 5364 1854
rect 5346 1854 5364 1872
rect 5346 1872 5364 1890
rect 5346 1890 5364 1908
rect 5346 1908 5364 1926
rect 5346 1926 5364 1944
rect 5346 1944 5364 1962
rect 5346 1962 5364 1980
rect 5346 1980 5364 1998
rect 5346 1998 5364 2016
rect 5346 2016 5364 2034
rect 5346 2034 5364 2052
rect 5346 2052 5364 2070
rect 5346 2070 5364 2088
rect 5346 2088 5364 2106
rect 5346 2106 5364 2124
rect 5346 2124 5364 2142
rect 5346 2142 5364 2160
rect 5346 2160 5364 2178
rect 5346 2178 5364 2196
rect 5346 2196 5364 2214
rect 5346 2214 5364 2232
rect 5346 2232 5364 2250
rect 5346 2250 5364 2268
rect 5346 2268 5364 2286
rect 5346 2286 5364 2304
rect 5346 2304 5364 2322
rect 5346 2322 5364 2340
rect 5346 2340 5364 2358
rect 5346 2358 5364 2376
rect 5346 2376 5364 2394
rect 5346 2394 5364 2412
rect 5346 2412 5364 2430
rect 5346 2646 5364 2664
rect 5346 2664 5364 2682
rect 5346 2682 5364 2700
rect 5346 2700 5364 2718
rect 5346 2718 5364 2736
rect 5346 2736 5364 2754
rect 5346 2754 5364 2772
rect 5346 2772 5364 2790
rect 5346 2790 5364 2808
rect 5346 2808 5364 2826
rect 5346 2826 5364 2844
rect 5346 2844 5364 2862
rect 5346 2862 5364 2880
rect 5346 2880 5364 2898
rect 5346 2898 5364 2916
rect 5346 2916 5364 2934
rect 5346 2934 5364 2952
rect 5346 2952 5364 2970
rect 5346 2970 5364 2988
rect 5346 2988 5364 3006
rect 5346 3006 5364 3024
rect 5346 3024 5364 3042
rect 5346 3042 5364 3060
rect 5346 3060 5364 3078
rect 5346 3078 5364 3096
rect 5346 3096 5364 3114
rect 5346 3114 5364 3132
rect 5346 3132 5364 3150
rect 5346 3150 5364 3168
rect 5346 3168 5364 3186
rect 5346 3186 5364 3204
rect 5346 3204 5364 3222
rect 5346 3222 5364 3240
rect 5346 3240 5364 3258
rect 5346 3258 5364 3276
rect 5346 3276 5364 3294
rect 5346 3294 5364 3312
rect 5346 3312 5364 3330
rect 5346 3330 5364 3348
rect 5346 3348 5364 3366
rect 5346 3366 5364 3384
rect 5346 3384 5364 3402
rect 5346 3402 5364 3420
rect 5346 3420 5364 3438
rect 5346 3438 5364 3456
rect 5346 3456 5364 3474
rect 5346 3474 5364 3492
rect 5346 3492 5364 3510
rect 5346 3510 5364 3528
rect 5346 3528 5364 3546
rect 5346 3546 5364 3564
rect 5346 3564 5364 3582
rect 5346 3582 5364 3600
rect 5346 3600 5364 3618
rect 5346 3618 5364 3636
rect 5346 3636 5364 3654
rect 5346 3654 5364 3672
rect 5346 3672 5364 3690
rect 5346 3690 5364 3708
rect 5346 3708 5364 3726
rect 5346 3726 5364 3744
rect 5346 3744 5364 3762
rect 5346 3762 5364 3780
rect 5346 3780 5364 3798
rect 5346 3798 5364 3816
rect 5346 3816 5364 3834
rect 5346 3834 5364 3852
rect 5346 3852 5364 3870
rect 5346 3870 5364 3888
rect 5346 3888 5364 3906
rect 5346 3906 5364 3924
rect 5346 3924 5364 3942
rect 5346 3942 5364 3960
rect 5346 3960 5364 3978
rect 5346 3978 5364 3996
rect 5346 3996 5364 4014
rect 5346 4014 5364 4032
rect 5346 4032 5364 4050
rect 5346 4050 5364 4068
rect 5346 4068 5364 4086
rect 5346 4086 5364 4104
rect 5346 4104 5364 4122
rect 5346 4122 5364 4140
rect 5346 4140 5364 4158
rect 5346 4158 5364 4176
rect 5346 4176 5364 4194
rect 5346 4194 5364 4212
rect 5346 4212 5364 4230
rect 5346 4230 5364 4248
rect 5346 4248 5364 4266
rect 5346 4266 5364 4284
rect 5346 4284 5364 4302
rect 5346 4302 5364 4320
rect 5346 4320 5364 4338
rect 5346 4338 5364 4356
rect 5346 4356 5364 4374
rect 5346 4374 5364 4392
rect 5346 4392 5364 4410
rect 5346 4410 5364 4428
rect 5346 4428 5364 4446
rect 5346 4446 5364 4464
rect 5346 4464 5364 4482
rect 5346 4482 5364 4500
rect 5346 4500 5364 4518
rect 5346 4518 5364 4536
rect 5346 4536 5364 4554
rect 5346 4554 5364 4572
rect 5346 4572 5364 4590
rect 5346 4590 5364 4608
rect 5346 4608 5364 4626
rect 5346 4626 5364 4644
rect 5346 4644 5364 4662
rect 5346 4662 5364 4680
rect 5346 4680 5364 4698
rect 5346 4698 5364 4716
rect 5346 4716 5364 4734
rect 5346 4734 5364 4752
rect 5346 4968 5364 4986
rect 5346 4986 5364 5004
rect 5346 5004 5364 5022
rect 5346 5022 5364 5040
rect 5346 5040 5364 5058
rect 5346 5058 5364 5076
rect 5346 5076 5364 5094
rect 5346 5094 5364 5112
rect 5346 5112 5364 5130
rect 5346 5130 5364 5148
rect 5346 5148 5364 5166
rect 5346 5166 5364 5184
rect 5346 5184 5364 5202
rect 5346 5202 5364 5220
rect 5346 5220 5364 5238
rect 5346 5238 5364 5256
rect 5346 5256 5364 5274
rect 5346 5274 5364 5292
rect 5346 5292 5364 5310
rect 5346 5310 5364 5328
rect 5346 5328 5364 5346
rect 5346 5346 5364 5364
rect 5346 5364 5364 5382
rect 5346 5382 5364 5400
rect 5346 5400 5364 5418
rect 5346 5418 5364 5436
rect 5346 5436 5364 5454
rect 5346 5454 5364 5472
rect 5346 5472 5364 5490
rect 5346 5490 5364 5508
rect 5346 5508 5364 5526
rect 5346 5526 5364 5544
rect 5346 5544 5364 5562
rect 5346 5562 5364 5580
rect 5346 5580 5364 5598
rect 5346 5598 5364 5616
rect 5346 5616 5364 5634
rect 5346 5634 5364 5652
rect 5346 5652 5364 5670
rect 5346 5670 5364 5688
rect 5346 5688 5364 5706
rect 5346 5706 5364 5724
rect 5346 5724 5364 5742
rect 5346 5742 5364 5760
rect 5346 5760 5364 5778
rect 5346 5778 5364 5796
rect 5346 5796 5364 5814
rect 5346 5814 5364 5832
rect 5346 5832 5364 5850
rect 5346 5850 5364 5868
rect 5346 5868 5364 5886
rect 5346 5886 5364 5904
rect 5346 5904 5364 5922
rect 5346 5922 5364 5940
rect 5346 5940 5364 5958
rect 5346 5958 5364 5976
rect 5346 5976 5364 5994
rect 5346 5994 5364 6012
rect 5346 6012 5364 6030
rect 5346 6030 5364 6048
rect 5346 6048 5364 6066
rect 5346 6066 5364 6084
rect 5346 6084 5364 6102
rect 5346 6102 5364 6120
rect 5346 6120 5364 6138
rect 5346 6138 5364 6156
rect 5346 6156 5364 6174
rect 5346 6174 5364 6192
rect 5346 6192 5364 6210
rect 5346 6210 5364 6228
rect 5346 6228 5364 6246
rect 5346 6246 5364 6264
rect 5346 6264 5364 6282
rect 5346 6282 5364 6300
rect 5346 6300 5364 6318
rect 5346 6318 5364 6336
rect 5346 6336 5364 6354
rect 5346 6354 5364 6372
rect 5346 6372 5364 6390
rect 5346 6390 5364 6408
rect 5346 6408 5364 6426
rect 5346 6426 5364 6444
rect 5346 6444 5364 6462
rect 5346 6462 5364 6480
rect 5346 6480 5364 6498
rect 5346 6498 5364 6516
rect 5346 6516 5364 6534
rect 5346 6534 5364 6552
rect 5346 6552 5364 6570
rect 5346 6570 5364 6588
rect 5346 6588 5364 6606
rect 5346 6606 5364 6624
rect 5346 6624 5364 6642
rect 5346 6642 5364 6660
rect 5346 6660 5364 6678
rect 5346 6678 5364 6696
rect 5346 6696 5364 6714
rect 5346 6714 5364 6732
rect 5346 6732 5364 6750
rect 5346 6750 5364 6768
rect 5346 6768 5364 6786
rect 5346 6786 5364 6804
rect 5346 6804 5364 6822
rect 5346 6822 5364 6840
rect 5346 6840 5364 6858
rect 5346 6858 5364 6876
rect 5346 6876 5364 6894
rect 5346 6894 5364 6912
rect 5346 6912 5364 6930
rect 5346 6930 5364 6948
rect 5346 6948 5364 6966
rect 5346 6966 5364 6984
rect 5346 6984 5364 7002
rect 5346 7002 5364 7020
rect 5346 7020 5364 7038
rect 5346 7038 5364 7056
rect 5346 7056 5364 7074
rect 5346 7074 5364 7092
rect 5346 7092 5364 7110
rect 5346 7110 5364 7128
rect 5346 7128 5364 7146
rect 5346 7146 5364 7164
rect 5346 7164 5364 7182
rect 5346 7182 5364 7200
rect 5346 7200 5364 7218
rect 5346 7218 5364 7236
rect 5346 7236 5364 7254
rect 5346 7254 5364 7272
rect 5346 7272 5364 7290
rect 5346 7290 5364 7308
rect 5346 7308 5364 7326
rect 5346 7326 5364 7344
rect 5346 7344 5364 7362
rect 5346 7362 5364 7380
rect 5346 7380 5364 7398
rect 5346 7398 5364 7416
rect 5346 7416 5364 7434
rect 5346 7434 5364 7452
rect 5346 7452 5364 7470
rect 5346 7470 5364 7488
rect 5346 7488 5364 7506
rect 5346 7506 5364 7524
rect 5346 7524 5364 7542
rect 5346 7542 5364 7560
rect 5346 7560 5364 7578
rect 5346 7578 5364 7596
rect 5346 7596 5364 7614
rect 5346 7614 5364 7632
rect 5346 7632 5364 7650
rect 5346 7650 5364 7668
rect 5346 7668 5364 7686
rect 5346 7686 5364 7704
rect 5346 7704 5364 7722
rect 5346 7722 5364 7740
rect 5346 7740 5364 7758
rect 5346 7758 5364 7776
rect 5346 7776 5364 7794
rect 5346 7794 5364 7812
rect 5346 7812 5364 7830
rect 5346 7830 5364 7848
rect 5346 7848 5364 7866
rect 5346 7866 5364 7884
rect 5346 7884 5364 7902
rect 5346 7902 5364 7920
rect 5346 7920 5364 7938
rect 5346 7938 5364 7956
rect 5346 7956 5364 7974
rect 5346 7974 5364 7992
rect 5346 7992 5364 8010
rect 5346 8010 5364 8028
rect 5346 8028 5364 8046
rect 5346 8046 5364 8064
rect 5346 8064 5364 8082
rect 5346 8082 5364 8100
rect 5346 8100 5364 8118
rect 5346 8118 5364 8136
rect 5346 8136 5364 8154
rect 5346 8154 5364 8172
rect 5346 8172 5364 8190
rect 5346 8190 5364 8208
rect 5346 8208 5364 8226
rect 5346 8226 5364 8244
rect 5346 8244 5364 8262
rect 5346 8262 5364 8280
rect 5346 8280 5364 8298
rect 5346 8298 5364 8316
rect 5346 8316 5364 8334
rect 5346 8334 5364 8352
rect 5364 432 5382 450
rect 5364 450 5382 468
rect 5364 468 5382 486
rect 5364 486 5382 504
rect 5364 504 5382 522
rect 5364 522 5382 540
rect 5364 540 5382 558
rect 5364 558 5382 576
rect 5364 576 5382 594
rect 5364 594 5382 612
rect 5364 612 5382 630
rect 5364 630 5382 648
rect 5364 648 5382 666
rect 5364 666 5382 684
rect 5364 684 5382 702
rect 5364 702 5382 720
rect 5364 720 5382 738
rect 5364 738 5382 756
rect 5364 756 5382 774
rect 5364 774 5382 792
rect 5364 792 5382 810
rect 5364 810 5382 828
rect 5364 828 5382 846
rect 5364 846 5382 864
rect 5364 1008 5382 1026
rect 5364 1026 5382 1044
rect 5364 1044 5382 1062
rect 5364 1062 5382 1080
rect 5364 1080 5382 1098
rect 5364 1098 5382 1116
rect 5364 1116 5382 1134
rect 5364 1134 5382 1152
rect 5364 1152 5382 1170
rect 5364 1170 5382 1188
rect 5364 1188 5382 1206
rect 5364 1206 5382 1224
rect 5364 1224 5382 1242
rect 5364 1242 5382 1260
rect 5364 1260 5382 1278
rect 5364 1278 5382 1296
rect 5364 1296 5382 1314
rect 5364 1314 5382 1332
rect 5364 1332 5382 1350
rect 5364 1350 5382 1368
rect 5364 1368 5382 1386
rect 5364 1386 5382 1404
rect 5364 1404 5382 1422
rect 5364 1422 5382 1440
rect 5364 1440 5382 1458
rect 5364 1458 5382 1476
rect 5364 1476 5382 1494
rect 5364 1494 5382 1512
rect 5364 1512 5382 1530
rect 5364 1530 5382 1548
rect 5364 1548 5382 1566
rect 5364 1566 5382 1584
rect 5364 1584 5382 1602
rect 5364 1602 5382 1620
rect 5364 1620 5382 1638
rect 5364 1638 5382 1656
rect 5364 1656 5382 1674
rect 5364 1674 5382 1692
rect 5364 1692 5382 1710
rect 5364 1710 5382 1728
rect 5364 1728 5382 1746
rect 5364 1746 5382 1764
rect 5364 1764 5382 1782
rect 5364 1782 5382 1800
rect 5364 1800 5382 1818
rect 5364 1818 5382 1836
rect 5364 1836 5382 1854
rect 5364 1854 5382 1872
rect 5364 1872 5382 1890
rect 5364 1890 5382 1908
rect 5364 1908 5382 1926
rect 5364 1926 5382 1944
rect 5364 1944 5382 1962
rect 5364 1962 5382 1980
rect 5364 1980 5382 1998
rect 5364 1998 5382 2016
rect 5364 2016 5382 2034
rect 5364 2034 5382 2052
rect 5364 2052 5382 2070
rect 5364 2070 5382 2088
rect 5364 2088 5382 2106
rect 5364 2106 5382 2124
rect 5364 2124 5382 2142
rect 5364 2142 5382 2160
rect 5364 2160 5382 2178
rect 5364 2178 5382 2196
rect 5364 2196 5382 2214
rect 5364 2214 5382 2232
rect 5364 2232 5382 2250
rect 5364 2250 5382 2268
rect 5364 2268 5382 2286
rect 5364 2286 5382 2304
rect 5364 2304 5382 2322
rect 5364 2322 5382 2340
rect 5364 2340 5382 2358
rect 5364 2358 5382 2376
rect 5364 2376 5382 2394
rect 5364 2394 5382 2412
rect 5364 2412 5382 2430
rect 5364 2430 5382 2448
rect 5364 2646 5382 2664
rect 5364 2664 5382 2682
rect 5364 2682 5382 2700
rect 5364 2700 5382 2718
rect 5364 2718 5382 2736
rect 5364 2736 5382 2754
rect 5364 2754 5382 2772
rect 5364 2772 5382 2790
rect 5364 2790 5382 2808
rect 5364 2808 5382 2826
rect 5364 2826 5382 2844
rect 5364 2844 5382 2862
rect 5364 2862 5382 2880
rect 5364 2880 5382 2898
rect 5364 2898 5382 2916
rect 5364 2916 5382 2934
rect 5364 2934 5382 2952
rect 5364 2952 5382 2970
rect 5364 2970 5382 2988
rect 5364 2988 5382 3006
rect 5364 3006 5382 3024
rect 5364 3024 5382 3042
rect 5364 3042 5382 3060
rect 5364 3060 5382 3078
rect 5364 3078 5382 3096
rect 5364 3096 5382 3114
rect 5364 3114 5382 3132
rect 5364 3132 5382 3150
rect 5364 3150 5382 3168
rect 5364 3168 5382 3186
rect 5364 3186 5382 3204
rect 5364 3204 5382 3222
rect 5364 3222 5382 3240
rect 5364 3240 5382 3258
rect 5364 3258 5382 3276
rect 5364 3276 5382 3294
rect 5364 3294 5382 3312
rect 5364 3312 5382 3330
rect 5364 3330 5382 3348
rect 5364 3348 5382 3366
rect 5364 3366 5382 3384
rect 5364 3384 5382 3402
rect 5364 3402 5382 3420
rect 5364 3420 5382 3438
rect 5364 3438 5382 3456
rect 5364 3456 5382 3474
rect 5364 3474 5382 3492
rect 5364 3492 5382 3510
rect 5364 3510 5382 3528
rect 5364 3528 5382 3546
rect 5364 3546 5382 3564
rect 5364 3564 5382 3582
rect 5364 3582 5382 3600
rect 5364 3600 5382 3618
rect 5364 3618 5382 3636
rect 5364 3636 5382 3654
rect 5364 3654 5382 3672
rect 5364 3672 5382 3690
rect 5364 3690 5382 3708
rect 5364 3708 5382 3726
rect 5364 3726 5382 3744
rect 5364 3744 5382 3762
rect 5364 3762 5382 3780
rect 5364 3780 5382 3798
rect 5364 3798 5382 3816
rect 5364 3816 5382 3834
rect 5364 3834 5382 3852
rect 5364 3852 5382 3870
rect 5364 3870 5382 3888
rect 5364 3888 5382 3906
rect 5364 3906 5382 3924
rect 5364 3924 5382 3942
rect 5364 3942 5382 3960
rect 5364 3960 5382 3978
rect 5364 3978 5382 3996
rect 5364 3996 5382 4014
rect 5364 4014 5382 4032
rect 5364 4032 5382 4050
rect 5364 4050 5382 4068
rect 5364 4068 5382 4086
rect 5364 4086 5382 4104
rect 5364 4104 5382 4122
rect 5364 4122 5382 4140
rect 5364 4140 5382 4158
rect 5364 4158 5382 4176
rect 5364 4176 5382 4194
rect 5364 4194 5382 4212
rect 5364 4212 5382 4230
rect 5364 4230 5382 4248
rect 5364 4248 5382 4266
rect 5364 4266 5382 4284
rect 5364 4284 5382 4302
rect 5364 4302 5382 4320
rect 5364 4320 5382 4338
rect 5364 4338 5382 4356
rect 5364 4356 5382 4374
rect 5364 4374 5382 4392
rect 5364 4392 5382 4410
rect 5364 4410 5382 4428
rect 5364 4428 5382 4446
rect 5364 4446 5382 4464
rect 5364 4464 5382 4482
rect 5364 4482 5382 4500
rect 5364 4500 5382 4518
rect 5364 4518 5382 4536
rect 5364 4536 5382 4554
rect 5364 4554 5382 4572
rect 5364 4572 5382 4590
rect 5364 4590 5382 4608
rect 5364 4608 5382 4626
rect 5364 4626 5382 4644
rect 5364 4644 5382 4662
rect 5364 4662 5382 4680
rect 5364 4680 5382 4698
rect 5364 4698 5382 4716
rect 5364 4716 5382 4734
rect 5364 4734 5382 4752
rect 5364 4752 5382 4770
rect 5364 4986 5382 5004
rect 5364 5004 5382 5022
rect 5364 5022 5382 5040
rect 5364 5040 5382 5058
rect 5364 5058 5382 5076
rect 5364 5076 5382 5094
rect 5364 5094 5382 5112
rect 5364 5112 5382 5130
rect 5364 5130 5382 5148
rect 5364 5148 5382 5166
rect 5364 5166 5382 5184
rect 5364 5184 5382 5202
rect 5364 5202 5382 5220
rect 5364 5220 5382 5238
rect 5364 5238 5382 5256
rect 5364 5256 5382 5274
rect 5364 5274 5382 5292
rect 5364 5292 5382 5310
rect 5364 5310 5382 5328
rect 5364 5328 5382 5346
rect 5364 5346 5382 5364
rect 5364 5364 5382 5382
rect 5364 5382 5382 5400
rect 5364 5400 5382 5418
rect 5364 5418 5382 5436
rect 5364 5436 5382 5454
rect 5364 5454 5382 5472
rect 5364 5472 5382 5490
rect 5364 5490 5382 5508
rect 5364 5508 5382 5526
rect 5364 5526 5382 5544
rect 5364 5544 5382 5562
rect 5364 5562 5382 5580
rect 5364 5580 5382 5598
rect 5364 5598 5382 5616
rect 5364 5616 5382 5634
rect 5364 5634 5382 5652
rect 5364 5652 5382 5670
rect 5364 5670 5382 5688
rect 5364 5688 5382 5706
rect 5364 5706 5382 5724
rect 5364 5724 5382 5742
rect 5364 5742 5382 5760
rect 5364 5760 5382 5778
rect 5364 5778 5382 5796
rect 5364 5796 5382 5814
rect 5364 5814 5382 5832
rect 5364 5832 5382 5850
rect 5364 5850 5382 5868
rect 5364 5868 5382 5886
rect 5364 5886 5382 5904
rect 5364 5904 5382 5922
rect 5364 5922 5382 5940
rect 5364 5940 5382 5958
rect 5364 5958 5382 5976
rect 5364 5976 5382 5994
rect 5364 5994 5382 6012
rect 5364 6012 5382 6030
rect 5364 6030 5382 6048
rect 5364 6048 5382 6066
rect 5364 6066 5382 6084
rect 5364 6084 5382 6102
rect 5364 6102 5382 6120
rect 5364 6120 5382 6138
rect 5364 6138 5382 6156
rect 5364 6156 5382 6174
rect 5364 6174 5382 6192
rect 5364 6192 5382 6210
rect 5364 6210 5382 6228
rect 5364 6228 5382 6246
rect 5364 6246 5382 6264
rect 5364 6264 5382 6282
rect 5364 6282 5382 6300
rect 5364 6300 5382 6318
rect 5364 6318 5382 6336
rect 5364 6336 5382 6354
rect 5364 6354 5382 6372
rect 5364 6372 5382 6390
rect 5364 6390 5382 6408
rect 5364 6408 5382 6426
rect 5364 6426 5382 6444
rect 5364 6444 5382 6462
rect 5364 6462 5382 6480
rect 5364 6480 5382 6498
rect 5364 6498 5382 6516
rect 5364 6516 5382 6534
rect 5364 6534 5382 6552
rect 5364 6552 5382 6570
rect 5364 6570 5382 6588
rect 5364 6588 5382 6606
rect 5364 6606 5382 6624
rect 5364 6624 5382 6642
rect 5364 6642 5382 6660
rect 5364 6660 5382 6678
rect 5364 6678 5382 6696
rect 5364 6696 5382 6714
rect 5364 6714 5382 6732
rect 5364 6732 5382 6750
rect 5364 6750 5382 6768
rect 5364 6768 5382 6786
rect 5364 6786 5382 6804
rect 5364 6804 5382 6822
rect 5364 6822 5382 6840
rect 5364 6840 5382 6858
rect 5364 6858 5382 6876
rect 5364 6876 5382 6894
rect 5364 6894 5382 6912
rect 5364 6912 5382 6930
rect 5364 6930 5382 6948
rect 5364 6948 5382 6966
rect 5364 6966 5382 6984
rect 5364 6984 5382 7002
rect 5364 7002 5382 7020
rect 5364 7020 5382 7038
rect 5364 7038 5382 7056
rect 5364 7056 5382 7074
rect 5364 7074 5382 7092
rect 5364 7092 5382 7110
rect 5364 7110 5382 7128
rect 5364 7128 5382 7146
rect 5364 7146 5382 7164
rect 5364 7164 5382 7182
rect 5364 7182 5382 7200
rect 5364 7200 5382 7218
rect 5364 7218 5382 7236
rect 5364 7236 5382 7254
rect 5364 7254 5382 7272
rect 5364 7272 5382 7290
rect 5364 7290 5382 7308
rect 5364 7308 5382 7326
rect 5364 7326 5382 7344
rect 5364 7344 5382 7362
rect 5364 7362 5382 7380
rect 5364 7380 5382 7398
rect 5364 7398 5382 7416
rect 5364 7416 5382 7434
rect 5364 7434 5382 7452
rect 5364 7452 5382 7470
rect 5364 7470 5382 7488
rect 5364 7488 5382 7506
rect 5364 7506 5382 7524
rect 5364 7524 5382 7542
rect 5364 7542 5382 7560
rect 5364 7560 5382 7578
rect 5364 7578 5382 7596
rect 5364 7596 5382 7614
rect 5364 7614 5382 7632
rect 5364 7632 5382 7650
rect 5364 7650 5382 7668
rect 5364 7668 5382 7686
rect 5364 7686 5382 7704
rect 5364 7704 5382 7722
rect 5364 7722 5382 7740
rect 5364 7740 5382 7758
rect 5364 7758 5382 7776
rect 5364 7776 5382 7794
rect 5364 7794 5382 7812
rect 5364 7812 5382 7830
rect 5364 7830 5382 7848
rect 5364 7848 5382 7866
rect 5364 7866 5382 7884
rect 5364 7884 5382 7902
rect 5364 7902 5382 7920
rect 5364 7920 5382 7938
rect 5364 7938 5382 7956
rect 5364 7956 5382 7974
rect 5364 7974 5382 7992
rect 5364 7992 5382 8010
rect 5364 8010 5382 8028
rect 5364 8028 5382 8046
rect 5364 8046 5382 8064
rect 5364 8064 5382 8082
rect 5364 8082 5382 8100
rect 5364 8100 5382 8118
rect 5364 8118 5382 8136
rect 5364 8136 5382 8154
rect 5364 8154 5382 8172
rect 5364 8172 5382 8190
rect 5364 8190 5382 8208
rect 5364 8208 5382 8226
rect 5364 8226 5382 8244
rect 5364 8244 5382 8262
rect 5364 8262 5382 8280
rect 5364 8280 5382 8298
rect 5364 8298 5382 8316
rect 5364 8316 5382 8334
rect 5364 8334 5382 8352
rect 5364 8352 5382 8370
rect 5382 450 5400 468
rect 5382 468 5400 486
rect 5382 486 5400 504
rect 5382 504 5400 522
rect 5382 522 5400 540
rect 5382 540 5400 558
rect 5382 558 5400 576
rect 5382 576 5400 594
rect 5382 594 5400 612
rect 5382 612 5400 630
rect 5382 630 5400 648
rect 5382 648 5400 666
rect 5382 666 5400 684
rect 5382 684 5400 702
rect 5382 702 5400 720
rect 5382 720 5400 738
rect 5382 738 5400 756
rect 5382 756 5400 774
rect 5382 774 5400 792
rect 5382 792 5400 810
rect 5382 810 5400 828
rect 5382 828 5400 846
rect 5382 846 5400 864
rect 5382 864 5400 882
rect 5382 1008 5400 1026
rect 5382 1026 5400 1044
rect 5382 1044 5400 1062
rect 5382 1062 5400 1080
rect 5382 1080 5400 1098
rect 5382 1098 5400 1116
rect 5382 1116 5400 1134
rect 5382 1134 5400 1152
rect 5382 1152 5400 1170
rect 5382 1170 5400 1188
rect 5382 1188 5400 1206
rect 5382 1206 5400 1224
rect 5382 1224 5400 1242
rect 5382 1242 5400 1260
rect 5382 1260 5400 1278
rect 5382 1278 5400 1296
rect 5382 1296 5400 1314
rect 5382 1314 5400 1332
rect 5382 1332 5400 1350
rect 5382 1350 5400 1368
rect 5382 1368 5400 1386
rect 5382 1386 5400 1404
rect 5382 1404 5400 1422
rect 5382 1422 5400 1440
rect 5382 1440 5400 1458
rect 5382 1458 5400 1476
rect 5382 1476 5400 1494
rect 5382 1494 5400 1512
rect 5382 1512 5400 1530
rect 5382 1530 5400 1548
rect 5382 1548 5400 1566
rect 5382 1566 5400 1584
rect 5382 1584 5400 1602
rect 5382 1602 5400 1620
rect 5382 1620 5400 1638
rect 5382 1638 5400 1656
rect 5382 1656 5400 1674
rect 5382 1674 5400 1692
rect 5382 1692 5400 1710
rect 5382 1710 5400 1728
rect 5382 1728 5400 1746
rect 5382 1746 5400 1764
rect 5382 1764 5400 1782
rect 5382 1782 5400 1800
rect 5382 1800 5400 1818
rect 5382 1818 5400 1836
rect 5382 1836 5400 1854
rect 5382 1854 5400 1872
rect 5382 1872 5400 1890
rect 5382 1890 5400 1908
rect 5382 1908 5400 1926
rect 5382 1926 5400 1944
rect 5382 1944 5400 1962
rect 5382 1962 5400 1980
rect 5382 1980 5400 1998
rect 5382 1998 5400 2016
rect 5382 2016 5400 2034
rect 5382 2034 5400 2052
rect 5382 2052 5400 2070
rect 5382 2070 5400 2088
rect 5382 2088 5400 2106
rect 5382 2106 5400 2124
rect 5382 2124 5400 2142
rect 5382 2142 5400 2160
rect 5382 2160 5400 2178
rect 5382 2178 5400 2196
rect 5382 2196 5400 2214
rect 5382 2214 5400 2232
rect 5382 2232 5400 2250
rect 5382 2250 5400 2268
rect 5382 2268 5400 2286
rect 5382 2286 5400 2304
rect 5382 2304 5400 2322
rect 5382 2322 5400 2340
rect 5382 2340 5400 2358
rect 5382 2358 5400 2376
rect 5382 2376 5400 2394
rect 5382 2394 5400 2412
rect 5382 2412 5400 2430
rect 5382 2430 5400 2448
rect 5382 2664 5400 2682
rect 5382 2682 5400 2700
rect 5382 2700 5400 2718
rect 5382 2718 5400 2736
rect 5382 2736 5400 2754
rect 5382 2754 5400 2772
rect 5382 2772 5400 2790
rect 5382 2790 5400 2808
rect 5382 2808 5400 2826
rect 5382 2826 5400 2844
rect 5382 2844 5400 2862
rect 5382 2862 5400 2880
rect 5382 2880 5400 2898
rect 5382 2898 5400 2916
rect 5382 2916 5400 2934
rect 5382 2934 5400 2952
rect 5382 2952 5400 2970
rect 5382 2970 5400 2988
rect 5382 2988 5400 3006
rect 5382 3006 5400 3024
rect 5382 3024 5400 3042
rect 5382 3042 5400 3060
rect 5382 3060 5400 3078
rect 5382 3078 5400 3096
rect 5382 3096 5400 3114
rect 5382 3114 5400 3132
rect 5382 3132 5400 3150
rect 5382 3150 5400 3168
rect 5382 3168 5400 3186
rect 5382 3186 5400 3204
rect 5382 3204 5400 3222
rect 5382 3222 5400 3240
rect 5382 3240 5400 3258
rect 5382 3258 5400 3276
rect 5382 3276 5400 3294
rect 5382 3294 5400 3312
rect 5382 3312 5400 3330
rect 5382 3330 5400 3348
rect 5382 3348 5400 3366
rect 5382 3366 5400 3384
rect 5382 3384 5400 3402
rect 5382 3402 5400 3420
rect 5382 3420 5400 3438
rect 5382 3438 5400 3456
rect 5382 3456 5400 3474
rect 5382 3474 5400 3492
rect 5382 3492 5400 3510
rect 5382 3510 5400 3528
rect 5382 3528 5400 3546
rect 5382 3546 5400 3564
rect 5382 3564 5400 3582
rect 5382 3582 5400 3600
rect 5382 3600 5400 3618
rect 5382 3618 5400 3636
rect 5382 3636 5400 3654
rect 5382 3654 5400 3672
rect 5382 3672 5400 3690
rect 5382 3690 5400 3708
rect 5382 3708 5400 3726
rect 5382 3726 5400 3744
rect 5382 3744 5400 3762
rect 5382 3762 5400 3780
rect 5382 3780 5400 3798
rect 5382 3798 5400 3816
rect 5382 3816 5400 3834
rect 5382 3834 5400 3852
rect 5382 3852 5400 3870
rect 5382 3870 5400 3888
rect 5382 3888 5400 3906
rect 5382 3906 5400 3924
rect 5382 3924 5400 3942
rect 5382 3942 5400 3960
rect 5382 3960 5400 3978
rect 5382 3978 5400 3996
rect 5382 3996 5400 4014
rect 5382 4014 5400 4032
rect 5382 4032 5400 4050
rect 5382 4050 5400 4068
rect 5382 4068 5400 4086
rect 5382 4086 5400 4104
rect 5382 4104 5400 4122
rect 5382 4122 5400 4140
rect 5382 4140 5400 4158
rect 5382 4158 5400 4176
rect 5382 4176 5400 4194
rect 5382 4194 5400 4212
rect 5382 4212 5400 4230
rect 5382 4230 5400 4248
rect 5382 4248 5400 4266
rect 5382 4266 5400 4284
rect 5382 4284 5400 4302
rect 5382 4302 5400 4320
rect 5382 4320 5400 4338
rect 5382 4338 5400 4356
rect 5382 4356 5400 4374
rect 5382 4374 5400 4392
rect 5382 4392 5400 4410
rect 5382 4410 5400 4428
rect 5382 4428 5400 4446
rect 5382 4446 5400 4464
rect 5382 4464 5400 4482
rect 5382 4482 5400 4500
rect 5382 4500 5400 4518
rect 5382 4518 5400 4536
rect 5382 4536 5400 4554
rect 5382 4554 5400 4572
rect 5382 4572 5400 4590
rect 5382 4590 5400 4608
rect 5382 4608 5400 4626
rect 5382 4626 5400 4644
rect 5382 4644 5400 4662
rect 5382 4662 5400 4680
rect 5382 4680 5400 4698
rect 5382 4698 5400 4716
rect 5382 4716 5400 4734
rect 5382 4734 5400 4752
rect 5382 4752 5400 4770
rect 5382 4770 5400 4788
rect 5382 5004 5400 5022
rect 5382 5022 5400 5040
rect 5382 5040 5400 5058
rect 5382 5058 5400 5076
rect 5382 5076 5400 5094
rect 5382 5094 5400 5112
rect 5382 5112 5400 5130
rect 5382 5130 5400 5148
rect 5382 5148 5400 5166
rect 5382 5166 5400 5184
rect 5382 5184 5400 5202
rect 5382 5202 5400 5220
rect 5382 5220 5400 5238
rect 5382 5238 5400 5256
rect 5382 5256 5400 5274
rect 5382 5274 5400 5292
rect 5382 5292 5400 5310
rect 5382 5310 5400 5328
rect 5382 5328 5400 5346
rect 5382 5346 5400 5364
rect 5382 5364 5400 5382
rect 5382 5382 5400 5400
rect 5382 5400 5400 5418
rect 5382 5418 5400 5436
rect 5382 5436 5400 5454
rect 5382 5454 5400 5472
rect 5382 5472 5400 5490
rect 5382 5490 5400 5508
rect 5382 5508 5400 5526
rect 5382 5526 5400 5544
rect 5382 5544 5400 5562
rect 5382 5562 5400 5580
rect 5382 5580 5400 5598
rect 5382 5598 5400 5616
rect 5382 5616 5400 5634
rect 5382 5634 5400 5652
rect 5382 5652 5400 5670
rect 5382 5670 5400 5688
rect 5382 5688 5400 5706
rect 5382 5706 5400 5724
rect 5382 5724 5400 5742
rect 5382 5742 5400 5760
rect 5382 5760 5400 5778
rect 5382 5778 5400 5796
rect 5382 5796 5400 5814
rect 5382 5814 5400 5832
rect 5382 5832 5400 5850
rect 5382 5850 5400 5868
rect 5382 5868 5400 5886
rect 5382 5886 5400 5904
rect 5382 5904 5400 5922
rect 5382 5922 5400 5940
rect 5382 5940 5400 5958
rect 5382 5958 5400 5976
rect 5382 5976 5400 5994
rect 5382 5994 5400 6012
rect 5382 6012 5400 6030
rect 5382 6030 5400 6048
rect 5382 6048 5400 6066
rect 5382 6066 5400 6084
rect 5382 6084 5400 6102
rect 5382 6102 5400 6120
rect 5382 6120 5400 6138
rect 5382 6138 5400 6156
rect 5382 6156 5400 6174
rect 5382 6174 5400 6192
rect 5382 6192 5400 6210
rect 5382 6210 5400 6228
rect 5382 6228 5400 6246
rect 5382 6246 5400 6264
rect 5382 6264 5400 6282
rect 5382 6282 5400 6300
rect 5382 6300 5400 6318
rect 5382 6318 5400 6336
rect 5382 6336 5400 6354
rect 5382 6354 5400 6372
rect 5382 6372 5400 6390
rect 5382 6390 5400 6408
rect 5382 6408 5400 6426
rect 5382 6426 5400 6444
rect 5382 6444 5400 6462
rect 5382 6462 5400 6480
rect 5382 6480 5400 6498
rect 5382 6498 5400 6516
rect 5382 6516 5400 6534
rect 5382 6534 5400 6552
rect 5382 6552 5400 6570
rect 5382 6570 5400 6588
rect 5382 6588 5400 6606
rect 5382 6606 5400 6624
rect 5382 6624 5400 6642
rect 5382 6642 5400 6660
rect 5382 6660 5400 6678
rect 5382 6678 5400 6696
rect 5382 6696 5400 6714
rect 5382 6714 5400 6732
rect 5382 6732 5400 6750
rect 5382 6750 5400 6768
rect 5382 6768 5400 6786
rect 5382 6786 5400 6804
rect 5382 6804 5400 6822
rect 5382 6822 5400 6840
rect 5382 6840 5400 6858
rect 5382 6858 5400 6876
rect 5382 6876 5400 6894
rect 5382 6894 5400 6912
rect 5382 6912 5400 6930
rect 5382 6930 5400 6948
rect 5382 6948 5400 6966
rect 5382 6966 5400 6984
rect 5382 6984 5400 7002
rect 5382 7002 5400 7020
rect 5382 7020 5400 7038
rect 5382 7038 5400 7056
rect 5382 7056 5400 7074
rect 5382 7074 5400 7092
rect 5382 7092 5400 7110
rect 5382 7110 5400 7128
rect 5382 7128 5400 7146
rect 5382 7146 5400 7164
rect 5382 7164 5400 7182
rect 5382 7182 5400 7200
rect 5382 7200 5400 7218
rect 5382 7218 5400 7236
rect 5382 7236 5400 7254
rect 5382 7254 5400 7272
rect 5382 7272 5400 7290
rect 5382 7290 5400 7308
rect 5382 7308 5400 7326
rect 5382 7326 5400 7344
rect 5382 7344 5400 7362
rect 5382 7362 5400 7380
rect 5382 7380 5400 7398
rect 5382 7398 5400 7416
rect 5382 7416 5400 7434
rect 5382 7434 5400 7452
rect 5382 7452 5400 7470
rect 5382 7470 5400 7488
rect 5382 7488 5400 7506
rect 5382 7506 5400 7524
rect 5382 7524 5400 7542
rect 5382 7542 5400 7560
rect 5382 7560 5400 7578
rect 5382 7578 5400 7596
rect 5382 7596 5400 7614
rect 5382 7614 5400 7632
rect 5382 7632 5400 7650
rect 5382 7650 5400 7668
rect 5382 7668 5400 7686
rect 5382 7686 5400 7704
rect 5382 7704 5400 7722
rect 5382 7722 5400 7740
rect 5382 7740 5400 7758
rect 5382 7758 5400 7776
rect 5382 7776 5400 7794
rect 5382 7794 5400 7812
rect 5382 7812 5400 7830
rect 5382 7830 5400 7848
rect 5382 7848 5400 7866
rect 5382 7866 5400 7884
rect 5382 7884 5400 7902
rect 5382 7902 5400 7920
rect 5382 7920 5400 7938
rect 5382 7938 5400 7956
rect 5382 7956 5400 7974
rect 5382 7974 5400 7992
rect 5382 7992 5400 8010
rect 5382 8010 5400 8028
rect 5382 8028 5400 8046
rect 5382 8046 5400 8064
rect 5382 8064 5400 8082
rect 5382 8082 5400 8100
rect 5382 8100 5400 8118
rect 5382 8118 5400 8136
rect 5382 8136 5400 8154
rect 5382 8154 5400 8172
rect 5382 8172 5400 8190
rect 5382 8190 5400 8208
rect 5382 8208 5400 8226
rect 5382 8226 5400 8244
rect 5382 8244 5400 8262
rect 5382 8262 5400 8280
rect 5382 8280 5400 8298
rect 5382 8298 5400 8316
rect 5382 8316 5400 8334
rect 5382 8334 5400 8352
rect 5382 8352 5400 8370
rect 5382 8370 5400 8388
rect 5382 8388 5400 8406
rect 5400 468 5418 486
rect 5400 486 5418 504
rect 5400 504 5418 522
rect 5400 522 5418 540
rect 5400 540 5418 558
rect 5400 558 5418 576
rect 5400 576 5418 594
rect 5400 594 5418 612
rect 5400 612 5418 630
rect 5400 630 5418 648
rect 5400 648 5418 666
rect 5400 666 5418 684
rect 5400 684 5418 702
rect 5400 702 5418 720
rect 5400 720 5418 738
rect 5400 738 5418 756
rect 5400 756 5418 774
rect 5400 774 5418 792
rect 5400 792 5418 810
rect 5400 810 5418 828
rect 5400 828 5418 846
rect 5400 846 5418 864
rect 5400 864 5418 882
rect 5400 1026 5418 1044
rect 5400 1044 5418 1062
rect 5400 1062 5418 1080
rect 5400 1080 5418 1098
rect 5400 1098 5418 1116
rect 5400 1116 5418 1134
rect 5400 1134 5418 1152
rect 5400 1152 5418 1170
rect 5400 1170 5418 1188
rect 5400 1188 5418 1206
rect 5400 1206 5418 1224
rect 5400 1224 5418 1242
rect 5400 1242 5418 1260
rect 5400 1260 5418 1278
rect 5400 1278 5418 1296
rect 5400 1296 5418 1314
rect 5400 1314 5418 1332
rect 5400 1332 5418 1350
rect 5400 1350 5418 1368
rect 5400 1368 5418 1386
rect 5400 1386 5418 1404
rect 5400 1404 5418 1422
rect 5400 1422 5418 1440
rect 5400 1440 5418 1458
rect 5400 1458 5418 1476
rect 5400 1476 5418 1494
rect 5400 1494 5418 1512
rect 5400 1512 5418 1530
rect 5400 1530 5418 1548
rect 5400 1548 5418 1566
rect 5400 1566 5418 1584
rect 5400 1584 5418 1602
rect 5400 1602 5418 1620
rect 5400 1620 5418 1638
rect 5400 1638 5418 1656
rect 5400 1656 5418 1674
rect 5400 1674 5418 1692
rect 5400 1692 5418 1710
rect 5400 1710 5418 1728
rect 5400 1728 5418 1746
rect 5400 1746 5418 1764
rect 5400 1764 5418 1782
rect 5400 1782 5418 1800
rect 5400 1800 5418 1818
rect 5400 1818 5418 1836
rect 5400 1836 5418 1854
rect 5400 1854 5418 1872
rect 5400 1872 5418 1890
rect 5400 1890 5418 1908
rect 5400 1908 5418 1926
rect 5400 1926 5418 1944
rect 5400 1944 5418 1962
rect 5400 1962 5418 1980
rect 5400 1980 5418 1998
rect 5400 1998 5418 2016
rect 5400 2016 5418 2034
rect 5400 2034 5418 2052
rect 5400 2052 5418 2070
rect 5400 2070 5418 2088
rect 5400 2088 5418 2106
rect 5400 2106 5418 2124
rect 5400 2124 5418 2142
rect 5400 2142 5418 2160
rect 5400 2160 5418 2178
rect 5400 2178 5418 2196
rect 5400 2196 5418 2214
rect 5400 2214 5418 2232
rect 5400 2232 5418 2250
rect 5400 2250 5418 2268
rect 5400 2268 5418 2286
rect 5400 2286 5418 2304
rect 5400 2304 5418 2322
rect 5400 2322 5418 2340
rect 5400 2340 5418 2358
rect 5400 2358 5418 2376
rect 5400 2376 5418 2394
rect 5400 2394 5418 2412
rect 5400 2412 5418 2430
rect 5400 2430 5418 2448
rect 5400 2448 5418 2466
rect 5400 2664 5418 2682
rect 5400 2682 5418 2700
rect 5400 2700 5418 2718
rect 5400 2718 5418 2736
rect 5400 2736 5418 2754
rect 5400 2754 5418 2772
rect 5400 2772 5418 2790
rect 5400 2790 5418 2808
rect 5400 2808 5418 2826
rect 5400 2826 5418 2844
rect 5400 2844 5418 2862
rect 5400 2862 5418 2880
rect 5400 2880 5418 2898
rect 5400 2898 5418 2916
rect 5400 2916 5418 2934
rect 5400 2934 5418 2952
rect 5400 2952 5418 2970
rect 5400 2970 5418 2988
rect 5400 2988 5418 3006
rect 5400 3006 5418 3024
rect 5400 3024 5418 3042
rect 5400 3042 5418 3060
rect 5400 3060 5418 3078
rect 5400 3078 5418 3096
rect 5400 3096 5418 3114
rect 5400 3114 5418 3132
rect 5400 3132 5418 3150
rect 5400 3150 5418 3168
rect 5400 3168 5418 3186
rect 5400 3186 5418 3204
rect 5400 3204 5418 3222
rect 5400 3222 5418 3240
rect 5400 3240 5418 3258
rect 5400 3258 5418 3276
rect 5400 3276 5418 3294
rect 5400 3294 5418 3312
rect 5400 3312 5418 3330
rect 5400 3330 5418 3348
rect 5400 3348 5418 3366
rect 5400 3366 5418 3384
rect 5400 3384 5418 3402
rect 5400 3402 5418 3420
rect 5400 3420 5418 3438
rect 5400 3438 5418 3456
rect 5400 3456 5418 3474
rect 5400 3474 5418 3492
rect 5400 3492 5418 3510
rect 5400 3510 5418 3528
rect 5400 3528 5418 3546
rect 5400 3546 5418 3564
rect 5400 3564 5418 3582
rect 5400 3582 5418 3600
rect 5400 3600 5418 3618
rect 5400 3618 5418 3636
rect 5400 3636 5418 3654
rect 5400 3654 5418 3672
rect 5400 3672 5418 3690
rect 5400 3690 5418 3708
rect 5400 3708 5418 3726
rect 5400 3726 5418 3744
rect 5400 3744 5418 3762
rect 5400 3762 5418 3780
rect 5400 3780 5418 3798
rect 5400 3798 5418 3816
rect 5400 3816 5418 3834
rect 5400 3834 5418 3852
rect 5400 3852 5418 3870
rect 5400 3870 5418 3888
rect 5400 3888 5418 3906
rect 5400 3906 5418 3924
rect 5400 3924 5418 3942
rect 5400 3942 5418 3960
rect 5400 3960 5418 3978
rect 5400 3978 5418 3996
rect 5400 3996 5418 4014
rect 5400 4014 5418 4032
rect 5400 4032 5418 4050
rect 5400 4050 5418 4068
rect 5400 4068 5418 4086
rect 5400 4086 5418 4104
rect 5400 4104 5418 4122
rect 5400 4122 5418 4140
rect 5400 4140 5418 4158
rect 5400 4158 5418 4176
rect 5400 4176 5418 4194
rect 5400 4194 5418 4212
rect 5400 4212 5418 4230
rect 5400 4230 5418 4248
rect 5400 4248 5418 4266
rect 5400 4266 5418 4284
rect 5400 4284 5418 4302
rect 5400 4302 5418 4320
rect 5400 4320 5418 4338
rect 5400 4338 5418 4356
rect 5400 4356 5418 4374
rect 5400 4374 5418 4392
rect 5400 4392 5418 4410
rect 5400 4410 5418 4428
rect 5400 4428 5418 4446
rect 5400 4446 5418 4464
rect 5400 4464 5418 4482
rect 5400 4482 5418 4500
rect 5400 4500 5418 4518
rect 5400 4518 5418 4536
rect 5400 4536 5418 4554
rect 5400 4554 5418 4572
rect 5400 4572 5418 4590
rect 5400 4590 5418 4608
rect 5400 4608 5418 4626
rect 5400 4626 5418 4644
rect 5400 4644 5418 4662
rect 5400 4662 5418 4680
rect 5400 4680 5418 4698
rect 5400 4698 5418 4716
rect 5400 4716 5418 4734
rect 5400 4734 5418 4752
rect 5400 4752 5418 4770
rect 5400 4770 5418 4788
rect 5400 4788 5418 4806
rect 5400 5022 5418 5040
rect 5400 5040 5418 5058
rect 5400 5058 5418 5076
rect 5400 5076 5418 5094
rect 5400 5094 5418 5112
rect 5400 5112 5418 5130
rect 5400 5130 5418 5148
rect 5400 5148 5418 5166
rect 5400 5166 5418 5184
rect 5400 5184 5418 5202
rect 5400 5202 5418 5220
rect 5400 5220 5418 5238
rect 5400 5238 5418 5256
rect 5400 5256 5418 5274
rect 5400 5274 5418 5292
rect 5400 5292 5418 5310
rect 5400 5310 5418 5328
rect 5400 5328 5418 5346
rect 5400 5346 5418 5364
rect 5400 5364 5418 5382
rect 5400 5382 5418 5400
rect 5400 5400 5418 5418
rect 5400 5418 5418 5436
rect 5400 5436 5418 5454
rect 5400 5454 5418 5472
rect 5400 5472 5418 5490
rect 5400 5490 5418 5508
rect 5400 5508 5418 5526
rect 5400 5526 5418 5544
rect 5400 5544 5418 5562
rect 5400 5562 5418 5580
rect 5400 5580 5418 5598
rect 5400 5598 5418 5616
rect 5400 5616 5418 5634
rect 5400 5634 5418 5652
rect 5400 5652 5418 5670
rect 5400 5670 5418 5688
rect 5400 5688 5418 5706
rect 5400 5706 5418 5724
rect 5400 5724 5418 5742
rect 5400 5742 5418 5760
rect 5400 5760 5418 5778
rect 5400 5778 5418 5796
rect 5400 5796 5418 5814
rect 5400 5814 5418 5832
rect 5400 5832 5418 5850
rect 5400 5850 5418 5868
rect 5400 5868 5418 5886
rect 5400 5886 5418 5904
rect 5400 5904 5418 5922
rect 5400 5922 5418 5940
rect 5400 5940 5418 5958
rect 5400 5958 5418 5976
rect 5400 5976 5418 5994
rect 5400 5994 5418 6012
rect 5400 6012 5418 6030
rect 5400 6030 5418 6048
rect 5400 6048 5418 6066
rect 5400 6066 5418 6084
rect 5400 6084 5418 6102
rect 5400 6102 5418 6120
rect 5400 6120 5418 6138
rect 5400 6138 5418 6156
rect 5400 6156 5418 6174
rect 5400 6174 5418 6192
rect 5400 6192 5418 6210
rect 5400 6210 5418 6228
rect 5400 6228 5418 6246
rect 5400 6246 5418 6264
rect 5400 6264 5418 6282
rect 5400 6282 5418 6300
rect 5400 6300 5418 6318
rect 5400 6318 5418 6336
rect 5400 6336 5418 6354
rect 5400 6354 5418 6372
rect 5400 6372 5418 6390
rect 5400 6390 5418 6408
rect 5400 6408 5418 6426
rect 5400 6426 5418 6444
rect 5400 6444 5418 6462
rect 5400 6462 5418 6480
rect 5400 6480 5418 6498
rect 5400 6498 5418 6516
rect 5400 6516 5418 6534
rect 5400 6534 5418 6552
rect 5400 6552 5418 6570
rect 5400 6570 5418 6588
rect 5400 6588 5418 6606
rect 5400 6606 5418 6624
rect 5400 6624 5418 6642
rect 5400 6642 5418 6660
rect 5400 6660 5418 6678
rect 5400 6678 5418 6696
rect 5400 6696 5418 6714
rect 5400 6714 5418 6732
rect 5400 6732 5418 6750
rect 5400 6750 5418 6768
rect 5400 6768 5418 6786
rect 5400 6786 5418 6804
rect 5400 6804 5418 6822
rect 5400 6822 5418 6840
rect 5400 6840 5418 6858
rect 5400 6858 5418 6876
rect 5400 6876 5418 6894
rect 5400 6894 5418 6912
rect 5400 6912 5418 6930
rect 5400 6930 5418 6948
rect 5400 6948 5418 6966
rect 5400 6966 5418 6984
rect 5400 6984 5418 7002
rect 5400 7002 5418 7020
rect 5400 7020 5418 7038
rect 5400 7038 5418 7056
rect 5400 7056 5418 7074
rect 5400 7074 5418 7092
rect 5400 7092 5418 7110
rect 5400 7110 5418 7128
rect 5400 7128 5418 7146
rect 5400 7146 5418 7164
rect 5400 7164 5418 7182
rect 5400 7182 5418 7200
rect 5400 7200 5418 7218
rect 5400 7218 5418 7236
rect 5400 7236 5418 7254
rect 5400 7254 5418 7272
rect 5400 7272 5418 7290
rect 5400 7290 5418 7308
rect 5400 7308 5418 7326
rect 5400 7326 5418 7344
rect 5400 7344 5418 7362
rect 5400 7362 5418 7380
rect 5400 7380 5418 7398
rect 5400 7398 5418 7416
rect 5400 7416 5418 7434
rect 5400 7434 5418 7452
rect 5400 7452 5418 7470
rect 5400 7470 5418 7488
rect 5400 7488 5418 7506
rect 5400 7506 5418 7524
rect 5400 7524 5418 7542
rect 5400 7542 5418 7560
rect 5400 7560 5418 7578
rect 5400 7578 5418 7596
rect 5400 7596 5418 7614
rect 5400 7614 5418 7632
rect 5400 7632 5418 7650
rect 5400 7650 5418 7668
rect 5400 7668 5418 7686
rect 5400 7686 5418 7704
rect 5400 7704 5418 7722
rect 5400 7722 5418 7740
rect 5400 7740 5418 7758
rect 5400 7758 5418 7776
rect 5400 7776 5418 7794
rect 5400 7794 5418 7812
rect 5400 7812 5418 7830
rect 5400 7830 5418 7848
rect 5400 7848 5418 7866
rect 5400 7866 5418 7884
rect 5400 7884 5418 7902
rect 5400 7902 5418 7920
rect 5400 7920 5418 7938
rect 5400 7938 5418 7956
rect 5400 7956 5418 7974
rect 5400 7974 5418 7992
rect 5400 7992 5418 8010
rect 5400 8010 5418 8028
rect 5400 8028 5418 8046
rect 5400 8046 5418 8064
rect 5400 8064 5418 8082
rect 5400 8082 5418 8100
rect 5400 8100 5418 8118
rect 5400 8118 5418 8136
rect 5400 8136 5418 8154
rect 5400 8154 5418 8172
rect 5400 8172 5418 8190
rect 5400 8190 5418 8208
rect 5400 8208 5418 8226
rect 5400 8226 5418 8244
rect 5400 8244 5418 8262
rect 5400 8262 5418 8280
rect 5400 8280 5418 8298
rect 5400 8298 5418 8316
rect 5400 8316 5418 8334
rect 5400 8334 5418 8352
rect 5400 8352 5418 8370
rect 5400 8370 5418 8388
rect 5400 8388 5418 8406
rect 5400 8406 5418 8424
rect 5418 468 5436 486
rect 5418 486 5436 504
rect 5418 504 5436 522
rect 5418 522 5436 540
rect 5418 540 5436 558
rect 5418 558 5436 576
rect 5418 576 5436 594
rect 5418 594 5436 612
rect 5418 612 5436 630
rect 5418 630 5436 648
rect 5418 648 5436 666
rect 5418 666 5436 684
rect 5418 684 5436 702
rect 5418 702 5436 720
rect 5418 720 5436 738
rect 5418 738 5436 756
rect 5418 756 5436 774
rect 5418 774 5436 792
rect 5418 792 5436 810
rect 5418 810 5436 828
rect 5418 828 5436 846
rect 5418 846 5436 864
rect 5418 864 5436 882
rect 5418 1026 5436 1044
rect 5418 1044 5436 1062
rect 5418 1062 5436 1080
rect 5418 1080 5436 1098
rect 5418 1098 5436 1116
rect 5418 1116 5436 1134
rect 5418 1134 5436 1152
rect 5418 1152 5436 1170
rect 5418 1170 5436 1188
rect 5418 1188 5436 1206
rect 5418 1206 5436 1224
rect 5418 1224 5436 1242
rect 5418 1242 5436 1260
rect 5418 1260 5436 1278
rect 5418 1278 5436 1296
rect 5418 1296 5436 1314
rect 5418 1314 5436 1332
rect 5418 1332 5436 1350
rect 5418 1350 5436 1368
rect 5418 1368 5436 1386
rect 5418 1386 5436 1404
rect 5418 1404 5436 1422
rect 5418 1422 5436 1440
rect 5418 1440 5436 1458
rect 5418 1458 5436 1476
rect 5418 1476 5436 1494
rect 5418 1494 5436 1512
rect 5418 1512 5436 1530
rect 5418 1530 5436 1548
rect 5418 1548 5436 1566
rect 5418 1566 5436 1584
rect 5418 1584 5436 1602
rect 5418 1602 5436 1620
rect 5418 1620 5436 1638
rect 5418 1638 5436 1656
rect 5418 1656 5436 1674
rect 5418 1674 5436 1692
rect 5418 1692 5436 1710
rect 5418 1710 5436 1728
rect 5418 1728 5436 1746
rect 5418 1746 5436 1764
rect 5418 1764 5436 1782
rect 5418 1782 5436 1800
rect 5418 1800 5436 1818
rect 5418 1818 5436 1836
rect 5418 1836 5436 1854
rect 5418 1854 5436 1872
rect 5418 1872 5436 1890
rect 5418 1890 5436 1908
rect 5418 1908 5436 1926
rect 5418 1926 5436 1944
rect 5418 1944 5436 1962
rect 5418 1962 5436 1980
rect 5418 1980 5436 1998
rect 5418 1998 5436 2016
rect 5418 2016 5436 2034
rect 5418 2034 5436 2052
rect 5418 2052 5436 2070
rect 5418 2070 5436 2088
rect 5418 2088 5436 2106
rect 5418 2106 5436 2124
rect 5418 2124 5436 2142
rect 5418 2142 5436 2160
rect 5418 2160 5436 2178
rect 5418 2178 5436 2196
rect 5418 2196 5436 2214
rect 5418 2214 5436 2232
rect 5418 2232 5436 2250
rect 5418 2250 5436 2268
rect 5418 2268 5436 2286
rect 5418 2286 5436 2304
rect 5418 2304 5436 2322
rect 5418 2322 5436 2340
rect 5418 2340 5436 2358
rect 5418 2358 5436 2376
rect 5418 2376 5436 2394
rect 5418 2394 5436 2412
rect 5418 2412 5436 2430
rect 5418 2430 5436 2448
rect 5418 2448 5436 2466
rect 5418 2466 5436 2484
rect 5418 2682 5436 2700
rect 5418 2700 5436 2718
rect 5418 2718 5436 2736
rect 5418 2736 5436 2754
rect 5418 2754 5436 2772
rect 5418 2772 5436 2790
rect 5418 2790 5436 2808
rect 5418 2808 5436 2826
rect 5418 2826 5436 2844
rect 5418 2844 5436 2862
rect 5418 2862 5436 2880
rect 5418 2880 5436 2898
rect 5418 2898 5436 2916
rect 5418 2916 5436 2934
rect 5418 2934 5436 2952
rect 5418 2952 5436 2970
rect 5418 2970 5436 2988
rect 5418 2988 5436 3006
rect 5418 3006 5436 3024
rect 5418 3024 5436 3042
rect 5418 3042 5436 3060
rect 5418 3060 5436 3078
rect 5418 3078 5436 3096
rect 5418 3096 5436 3114
rect 5418 3114 5436 3132
rect 5418 3132 5436 3150
rect 5418 3150 5436 3168
rect 5418 3168 5436 3186
rect 5418 3186 5436 3204
rect 5418 3204 5436 3222
rect 5418 3222 5436 3240
rect 5418 3240 5436 3258
rect 5418 3258 5436 3276
rect 5418 3276 5436 3294
rect 5418 3294 5436 3312
rect 5418 3312 5436 3330
rect 5418 3330 5436 3348
rect 5418 3348 5436 3366
rect 5418 3366 5436 3384
rect 5418 3384 5436 3402
rect 5418 3402 5436 3420
rect 5418 3420 5436 3438
rect 5418 3438 5436 3456
rect 5418 3456 5436 3474
rect 5418 3474 5436 3492
rect 5418 3492 5436 3510
rect 5418 3510 5436 3528
rect 5418 3528 5436 3546
rect 5418 3546 5436 3564
rect 5418 3564 5436 3582
rect 5418 3582 5436 3600
rect 5418 3600 5436 3618
rect 5418 3618 5436 3636
rect 5418 3636 5436 3654
rect 5418 3654 5436 3672
rect 5418 3672 5436 3690
rect 5418 3690 5436 3708
rect 5418 3708 5436 3726
rect 5418 3726 5436 3744
rect 5418 3744 5436 3762
rect 5418 3762 5436 3780
rect 5418 3780 5436 3798
rect 5418 3798 5436 3816
rect 5418 3816 5436 3834
rect 5418 3834 5436 3852
rect 5418 3852 5436 3870
rect 5418 3870 5436 3888
rect 5418 3888 5436 3906
rect 5418 3906 5436 3924
rect 5418 3924 5436 3942
rect 5418 3942 5436 3960
rect 5418 3960 5436 3978
rect 5418 3978 5436 3996
rect 5418 3996 5436 4014
rect 5418 4014 5436 4032
rect 5418 4032 5436 4050
rect 5418 4050 5436 4068
rect 5418 4068 5436 4086
rect 5418 4086 5436 4104
rect 5418 4104 5436 4122
rect 5418 4122 5436 4140
rect 5418 4140 5436 4158
rect 5418 4158 5436 4176
rect 5418 4176 5436 4194
rect 5418 4194 5436 4212
rect 5418 4212 5436 4230
rect 5418 4230 5436 4248
rect 5418 4248 5436 4266
rect 5418 4266 5436 4284
rect 5418 4284 5436 4302
rect 5418 4302 5436 4320
rect 5418 4320 5436 4338
rect 5418 4338 5436 4356
rect 5418 4356 5436 4374
rect 5418 4374 5436 4392
rect 5418 4392 5436 4410
rect 5418 4410 5436 4428
rect 5418 4428 5436 4446
rect 5418 4446 5436 4464
rect 5418 4464 5436 4482
rect 5418 4482 5436 4500
rect 5418 4500 5436 4518
rect 5418 4518 5436 4536
rect 5418 4536 5436 4554
rect 5418 4554 5436 4572
rect 5418 4572 5436 4590
rect 5418 4590 5436 4608
rect 5418 4608 5436 4626
rect 5418 4626 5436 4644
rect 5418 4644 5436 4662
rect 5418 4662 5436 4680
rect 5418 4680 5436 4698
rect 5418 4698 5436 4716
rect 5418 4716 5436 4734
rect 5418 4734 5436 4752
rect 5418 4752 5436 4770
rect 5418 4770 5436 4788
rect 5418 4788 5436 4806
rect 5418 4806 5436 4824
rect 5418 5040 5436 5058
rect 5418 5058 5436 5076
rect 5418 5076 5436 5094
rect 5418 5094 5436 5112
rect 5418 5112 5436 5130
rect 5418 5130 5436 5148
rect 5418 5148 5436 5166
rect 5418 5166 5436 5184
rect 5418 5184 5436 5202
rect 5418 5202 5436 5220
rect 5418 5220 5436 5238
rect 5418 5238 5436 5256
rect 5418 5256 5436 5274
rect 5418 5274 5436 5292
rect 5418 5292 5436 5310
rect 5418 5310 5436 5328
rect 5418 5328 5436 5346
rect 5418 5346 5436 5364
rect 5418 5364 5436 5382
rect 5418 5382 5436 5400
rect 5418 5400 5436 5418
rect 5418 5418 5436 5436
rect 5418 5436 5436 5454
rect 5418 5454 5436 5472
rect 5418 5472 5436 5490
rect 5418 5490 5436 5508
rect 5418 5508 5436 5526
rect 5418 5526 5436 5544
rect 5418 5544 5436 5562
rect 5418 5562 5436 5580
rect 5418 5580 5436 5598
rect 5418 5598 5436 5616
rect 5418 5616 5436 5634
rect 5418 5634 5436 5652
rect 5418 5652 5436 5670
rect 5418 5670 5436 5688
rect 5418 5688 5436 5706
rect 5418 5706 5436 5724
rect 5418 5724 5436 5742
rect 5418 5742 5436 5760
rect 5418 5760 5436 5778
rect 5418 5778 5436 5796
rect 5418 5796 5436 5814
rect 5418 5814 5436 5832
rect 5418 5832 5436 5850
rect 5418 5850 5436 5868
rect 5418 5868 5436 5886
rect 5418 5886 5436 5904
rect 5418 5904 5436 5922
rect 5418 5922 5436 5940
rect 5418 5940 5436 5958
rect 5418 5958 5436 5976
rect 5418 5976 5436 5994
rect 5418 5994 5436 6012
rect 5418 6012 5436 6030
rect 5418 6030 5436 6048
rect 5418 6048 5436 6066
rect 5418 6066 5436 6084
rect 5418 6084 5436 6102
rect 5418 6102 5436 6120
rect 5418 6120 5436 6138
rect 5418 6138 5436 6156
rect 5418 6156 5436 6174
rect 5418 6174 5436 6192
rect 5418 6192 5436 6210
rect 5418 6210 5436 6228
rect 5418 6228 5436 6246
rect 5418 6246 5436 6264
rect 5418 6264 5436 6282
rect 5418 6282 5436 6300
rect 5418 6300 5436 6318
rect 5418 6318 5436 6336
rect 5418 6336 5436 6354
rect 5418 6354 5436 6372
rect 5418 6372 5436 6390
rect 5418 6390 5436 6408
rect 5418 6408 5436 6426
rect 5418 6426 5436 6444
rect 5418 6444 5436 6462
rect 5418 6462 5436 6480
rect 5418 6480 5436 6498
rect 5418 6498 5436 6516
rect 5418 6516 5436 6534
rect 5418 6534 5436 6552
rect 5418 6552 5436 6570
rect 5418 6570 5436 6588
rect 5418 6588 5436 6606
rect 5418 6606 5436 6624
rect 5418 6624 5436 6642
rect 5418 6642 5436 6660
rect 5418 6660 5436 6678
rect 5418 6678 5436 6696
rect 5418 6696 5436 6714
rect 5418 6714 5436 6732
rect 5418 6732 5436 6750
rect 5418 6750 5436 6768
rect 5418 6768 5436 6786
rect 5418 6786 5436 6804
rect 5418 6804 5436 6822
rect 5418 6822 5436 6840
rect 5418 6840 5436 6858
rect 5418 6858 5436 6876
rect 5418 6876 5436 6894
rect 5418 6894 5436 6912
rect 5418 6912 5436 6930
rect 5418 6930 5436 6948
rect 5418 6948 5436 6966
rect 5418 6966 5436 6984
rect 5418 6984 5436 7002
rect 5418 7002 5436 7020
rect 5418 7020 5436 7038
rect 5418 7038 5436 7056
rect 5418 7056 5436 7074
rect 5418 7074 5436 7092
rect 5418 7092 5436 7110
rect 5418 7110 5436 7128
rect 5418 7128 5436 7146
rect 5418 7146 5436 7164
rect 5418 7164 5436 7182
rect 5418 7182 5436 7200
rect 5418 7200 5436 7218
rect 5418 7218 5436 7236
rect 5418 7236 5436 7254
rect 5418 7254 5436 7272
rect 5418 7272 5436 7290
rect 5418 7290 5436 7308
rect 5418 7308 5436 7326
rect 5418 7326 5436 7344
rect 5418 7344 5436 7362
rect 5418 7362 5436 7380
rect 5418 7380 5436 7398
rect 5418 7398 5436 7416
rect 5418 7416 5436 7434
rect 5418 7434 5436 7452
rect 5418 7452 5436 7470
rect 5418 7470 5436 7488
rect 5418 7488 5436 7506
rect 5418 7506 5436 7524
rect 5418 7524 5436 7542
rect 5418 7542 5436 7560
rect 5418 7560 5436 7578
rect 5418 7578 5436 7596
rect 5418 7596 5436 7614
rect 5418 7614 5436 7632
rect 5418 7632 5436 7650
rect 5418 7650 5436 7668
rect 5418 7668 5436 7686
rect 5418 7686 5436 7704
rect 5418 7704 5436 7722
rect 5418 7722 5436 7740
rect 5418 7740 5436 7758
rect 5418 7758 5436 7776
rect 5418 7776 5436 7794
rect 5418 7794 5436 7812
rect 5418 7812 5436 7830
rect 5418 7830 5436 7848
rect 5418 7848 5436 7866
rect 5418 7866 5436 7884
rect 5418 7884 5436 7902
rect 5418 7902 5436 7920
rect 5418 7920 5436 7938
rect 5418 7938 5436 7956
rect 5418 7956 5436 7974
rect 5418 7974 5436 7992
rect 5418 7992 5436 8010
rect 5418 8010 5436 8028
rect 5418 8028 5436 8046
rect 5418 8046 5436 8064
rect 5418 8064 5436 8082
rect 5418 8082 5436 8100
rect 5418 8100 5436 8118
rect 5418 8118 5436 8136
rect 5418 8136 5436 8154
rect 5418 8154 5436 8172
rect 5418 8172 5436 8190
rect 5418 8190 5436 8208
rect 5418 8208 5436 8226
rect 5418 8226 5436 8244
rect 5418 8244 5436 8262
rect 5418 8262 5436 8280
rect 5418 8280 5436 8298
rect 5418 8298 5436 8316
rect 5418 8316 5436 8334
rect 5418 8334 5436 8352
rect 5418 8352 5436 8370
rect 5418 8370 5436 8388
rect 5418 8388 5436 8406
rect 5418 8406 5436 8424
rect 5418 8424 5436 8442
rect 5436 486 5454 504
rect 5436 504 5454 522
rect 5436 522 5454 540
rect 5436 540 5454 558
rect 5436 558 5454 576
rect 5436 576 5454 594
rect 5436 594 5454 612
rect 5436 612 5454 630
rect 5436 630 5454 648
rect 5436 648 5454 666
rect 5436 666 5454 684
rect 5436 684 5454 702
rect 5436 702 5454 720
rect 5436 720 5454 738
rect 5436 738 5454 756
rect 5436 756 5454 774
rect 5436 774 5454 792
rect 5436 792 5454 810
rect 5436 810 5454 828
rect 5436 828 5454 846
rect 5436 846 5454 864
rect 5436 864 5454 882
rect 5436 882 5454 900
rect 5436 1026 5454 1044
rect 5436 1044 5454 1062
rect 5436 1062 5454 1080
rect 5436 1080 5454 1098
rect 5436 1098 5454 1116
rect 5436 1116 5454 1134
rect 5436 1134 5454 1152
rect 5436 1152 5454 1170
rect 5436 1170 5454 1188
rect 5436 1188 5454 1206
rect 5436 1206 5454 1224
rect 5436 1224 5454 1242
rect 5436 1242 5454 1260
rect 5436 1260 5454 1278
rect 5436 1278 5454 1296
rect 5436 1296 5454 1314
rect 5436 1314 5454 1332
rect 5436 1332 5454 1350
rect 5436 1350 5454 1368
rect 5436 1368 5454 1386
rect 5436 1386 5454 1404
rect 5436 1404 5454 1422
rect 5436 1422 5454 1440
rect 5436 1440 5454 1458
rect 5436 1458 5454 1476
rect 5436 1476 5454 1494
rect 5436 1494 5454 1512
rect 5436 1512 5454 1530
rect 5436 1530 5454 1548
rect 5436 1548 5454 1566
rect 5436 1566 5454 1584
rect 5436 1584 5454 1602
rect 5436 1602 5454 1620
rect 5436 1620 5454 1638
rect 5436 1638 5454 1656
rect 5436 1656 5454 1674
rect 5436 1674 5454 1692
rect 5436 1692 5454 1710
rect 5436 1710 5454 1728
rect 5436 1728 5454 1746
rect 5436 1746 5454 1764
rect 5436 1764 5454 1782
rect 5436 1782 5454 1800
rect 5436 1800 5454 1818
rect 5436 1818 5454 1836
rect 5436 1836 5454 1854
rect 5436 1854 5454 1872
rect 5436 1872 5454 1890
rect 5436 1890 5454 1908
rect 5436 1908 5454 1926
rect 5436 1926 5454 1944
rect 5436 1944 5454 1962
rect 5436 1962 5454 1980
rect 5436 1980 5454 1998
rect 5436 1998 5454 2016
rect 5436 2016 5454 2034
rect 5436 2034 5454 2052
rect 5436 2052 5454 2070
rect 5436 2070 5454 2088
rect 5436 2088 5454 2106
rect 5436 2106 5454 2124
rect 5436 2124 5454 2142
rect 5436 2142 5454 2160
rect 5436 2160 5454 2178
rect 5436 2178 5454 2196
rect 5436 2196 5454 2214
rect 5436 2214 5454 2232
rect 5436 2232 5454 2250
rect 5436 2250 5454 2268
rect 5436 2268 5454 2286
rect 5436 2286 5454 2304
rect 5436 2304 5454 2322
rect 5436 2322 5454 2340
rect 5436 2340 5454 2358
rect 5436 2358 5454 2376
rect 5436 2376 5454 2394
rect 5436 2394 5454 2412
rect 5436 2412 5454 2430
rect 5436 2430 5454 2448
rect 5436 2448 5454 2466
rect 5436 2466 5454 2484
rect 5436 2682 5454 2700
rect 5436 2700 5454 2718
rect 5436 2718 5454 2736
rect 5436 2736 5454 2754
rect 5436 2754 5454 2772
rect 5436 2772 5454 2790
rect 5436 2790 5454 2808
rect 5436 2808 5454 2826
rect 5436 2826 5454 2844
rect 5436 2844 5454 2862
rect 5436 2862 5454 2880
rect 5436 2880 5454 2898
rect 5436 2898 5454 2916
rect 5436 2916 5454 2934
rect 5436 2934 5454 2952
rect 5436 2952 5454 2970
rect 5436 2970 5454 2988
rect 5436 2988 5454 3006
rect 5436 3006 5454 3024
rect 5436 3024 5454 3042
rect 5436 3042 5454 3060
rect 5436 3060 5454 3078
rect 5436 3078 5454 3096
rect 5436 3096 5454 3114
rect 5436 3114 5454 3132
rect 5436 3132 5454 3150
rect 5436 3150 5454 3168
rect 5436 3168 5454 3186
rect 5436 3186 5454 3204
rect 5436 3204 5454 3222
rect 5436 3222 5454 3240
rect 5436 3240 5454 3258
rect 5436 3258 5454 3276
rect 5436 3276 5454 3294
rect 5436 3294 5454 3312
rect 5436 3312 5454 3330
rect 5436 3330 5454 3348
rect 5436 3348 5454 3366
rect 5436 3366 5454 3384
rect 5436 3384 5454 3402
rect 5436 3402 5454 3420
rect 5436 3420 5454 3438
rect 5436 3438 5454 3456
rect 5436 3456 5454 3474
rect 5436 3474 5454 3492
rect 5436 3492 5454 3510
rect 5436 3510 5454 3528
rect 5436 3528 5454 3546
rect 5436 3546 5454 3564
rect 5436 3564 5454 3582
rect 5436 3582 5454 3600
rect 5436 3600 5454 3618
rect 5436 3618 5454 3636
rect 5436 3636 5454 3654
rect 5436 3654 5454 3672
rect 5436 3672 5454 3690
rect 5436 3690 5454 3708
rect 5436 3708 5454 3726
rect 5436 3726 5454 3744
rect 5436 3744 5454 3762
rect 5436 3762 5454 3780
rect 5436 3780 5454 3798
rect 5436 3798 5454 3816
rect 5436 3816 5454 3834
rect 5436 3834 5454 3852
rect 5436 3852 5454 3870
rect 5436 3870 5454 3888
rect 5436 3888 5454 3906
rect 5436 3906 5454 3924
rect 5436 3924 5454 3942
rect 5436 3942 5454 3960
rect 5436 3960 5454 3978
rect 5436 3978 5454 3996
rect 5436 3996 5454 4014
rect 5436 4014 5454 4032
rect 5436 4032 5454 4050
rect 5436 4050 5454 4068
rect 5436 4068 5454 4086
rect 5436 4086 5454 4104
rect 5436 4104 5454 4122
rect 5436 4122 5454 4140
rect 5436 4140 5454 4158
rect 5436 4158 5454 4176
rect 5436 4176 5454 4194
rect 5436 4194 5454 4212
rect 5436 4212 5454 4230
rect 5436 4230 5454 4248
rect 5436 4248 5454 4266
rect 5436 4266 5454 4284
rect 5436 4284 5454 4302
rect 5436 4302 5454 4320
rect 5436 4320 5454 4338
rect 5436 4338 5454 4356
rect 5436 4356 5454 4374
rect 5436 4374 5454 4392
rect 5436 4392 5454 4410
rect 5436 4410 5454 4428
rect 5436 4428 5454 4446
rect 5436 4446 5454 4464
rect 5436 4464 5454 4482
rect 5436 4482 5454 4500
rect 5436 4500 5454 4518
rect 5436 4518 5454 4536
rect 5436 4536 5454 4554
rect 5436 4554 5454 4572
rect 5436 4572 5454 4590
rect 5436 4590 5454 4608
rect 5436 4608 5454 4626
rect 5436 4626 5454 4644
rect 5436 4644 5454 4662
rect 5436 4662 5454 4680
rect 5436 4680 5454 4698
rect 5436 4698 5454 4716
rect 5436 4716 5454 4734
rect 5436 4734 5454 4752
rect 5436 4752 5454 4770
rect 5436 4770 5454 4788
rect 5436 4788 5454 4806
rect 5436 4806 5454 4824
rect 5436 4824 5454 4842
rect 5436 5058 5454 5076
rect 5436 5076 5454 5094
rect 5436 5094 5454 5112
rect 5436 5112 5454 5130
rect 5436 5130 5454 5148
rect 5436 5148 5454 5166
rect 5436 5166 5454 5184
rect 5436 5184 5454 5202
rect 5436 5202 5454 5220
rect 5436 5220 5454 5238
rect 5436 5238 5454 5256
rect 5436 5256 5454 5274
rect 5436 5274 5454 5292
rect 5436 5292 5454 5310
rect 5436 5310 5454 5328
rect 5436 5328 5454 5346
rect 5436 5346 5454 5364
rect 5436 5364 5454 5382
rect 5436 5382 5454 5400
rect 5436 5400 5454 5418
rect 5436 5418 5454 5436
rect 5436 5436 5454 5454
rect 5436 5454 5454 5472
rect 5436 5472 5454 5490
rect 5436 5490 5454 5508
rect 5436 5508 5454 5526
rect 5436 5526 5454 5544
rect 5436 5544 5454 5562
rect 5436 5562 5454 5580
rect 5436 5580 5454 5598
rect 5436 5598 5454 5616
rect 5436 5616 5454 5634
rect 5436 5634 5454 5652
rect 5436 5652 5454 5670
rect 5436 5670 5454 5688
rect 5436 5688 5454 5706
rect 5436 5706 5454 5724
rect 5436 5724 5454 5742
rect 5436 5742 5454 5760
rect 5436 5760 5454 5778
rect 5436 5778 5454 5796
rect 5436 5796 5454 5814
rect 5436 5814 5454 5832
rect 5436 5832 5454 5850
rect 5436 5850 5454 5868
rect 5436 5868 5454 5886
rect 5436 5886 5454 5904
rect 5436 5904 5454 5922
rect 5436 5922 5454 5940
rect 5436 5940 5454 5958
rect 5436 5958 5454 5976
rect 5436 5976 5454 5994
rect 5436 5994 5454 6012
rect 5436 6012 5454 6030
rect 5436 6030 5454 6048
rect 5436 6048 5454 6066
rect 5436 6066 5454 6084
rect 5436 6084 5454 6102
rect 5436 6102 5454 6120
rect 5436 6120 5454 6138
rect 5436 6138 5454 6156
rect 5436 6156 5454 6174
rect 5436 6174 5454 6192
rect 5436 6192 5454 6210
rect 5436 6210 5454 6228
rect 5436 6228 5454 6246
rect 5436 6246 5454 6264
rect 5436 6264 5454 6282
rect 5436 6282 5454 6300
rect 5436 6300 5454 6318
rect 5436 6318 5454 6336
rect 5436 6336 5454 6354
rect 5436 6354 5454 6372
rect 5436 6372 5454 6390
rect 5436 6390 5454 6408
rect 5436 6408 5454 6426
rect 5436 6426 5454 6444
rect 5436 6444 5454 6462
rect 5436 6462 5454 6480
rect 5436 6480 5454 6498
rect 5436 6498 5454 6516
rect 5436 6516 5454 6534
rect 5436 6534 5454 6552
rect 5436 6552 5454 6570
rect 5436 6570 5454 6588
rect 5436 6588 5454 6606
rect 5436 6606 5454 6624
rect 5436 6624 5454 6642
rect 5436 6642 5454 6660
rect 5436 6660 5454 6678
rect 5436 6678 5454 6696
rect 5436 6696 5454 6714
rect 5436 6714 5454 6732
rect 5436 6732 5454 6750
rect 5436 6750 5454 6768
rect 5436 6768 5454 6786
rect 5436 6786 5454 6804
rect 5436 6804 5454 6822
rect 5436 6822 5454 6840
rect 5436 6840 5454 6858
rect 5436 6858 5454 6876
rect 5436 6876 5454 6894
rect 5436 6894 5454 6912
rect 5436 6912 5454 6930
rect 5436 6930 5454 6948
rect 5436 6948 5454 6966
rect 5436 6966 5454 6984
rect 5436 6984 5454 7002
rect 5436 7002 5454 7020
rect 5436 7020 5454 7038
rect 5436 7038 5454 7056
rect 5436 7056 5454 7074
rect 5436 7074 5454 7092
rect 5436 7092 5454 7110
rect 5436 7110 5454 7128
rect 5436 7128 5454 7146
rect 5436 7146 5454 7164
rect 5436 7164 5454 7182
rect 5436 7182 5454 7200
rect 5436 7200 5454 7218
rect 5436 7218 5454 7236
rect 5436 7236 5454 7254
rect 5436 7254 5454 7272
rect 5436 7272 5454 7290
rect 5436 7290 5454 7308
rect 5436 7308 5454 7326
rect 5436 7326 5454 7344
rect 5436 7344 5454 7362
rect 5436 7362 5454 7380
rect 5436 7380 5454 7398
rect 5436 7398 5454 7416
rect 5436 7416 5454 7434
rect 5436 7434 5454 7452
rect 5436 7452 5454 7470
rect 5436 7470 5454 7488
rect 5436 7488 5454 7506
rect 5436 7506 5454 7524
rect 5436 7524 5454 7542
rect 5436 7542 5454 7560
rect 5436 7560 5454 7578
rect 5436 7578 5454 7596
rect 5436 7596 5454 7614
rect 5436 7614 5454 7632
rect 5436 7632 5454 7650
rect 5436 7650 5454 7668
rect 5436 7668 5454 7686
rect 5436 7686 5454 7704
rect 5436 7704 5454 7722
rect 5436 7722 5454 7740
rect 5436 7740 5454 7758
rect 5436 7758 5454 7776
rect 5436 7776 5454 7794
rect 5436 7794 5454 7812
rect 5436 7812 5454 7830
rect 5436 7830 5454 7848
rect 5436 7848 5454 7866
rect 5436 7866 5454 7884
rect 5436 7884 5454 7902
rect 5436 7902 5454 7920
rect 5436 7920 5454 7938
rect 5436 7938 5454 7956
rect 5436 7956 5454 7974
rect 5436 7974 5454 7992
rect 5436 7992 5454 8010
rect 5436 8010 5454 8028
rect 5436 8028 5454 8046
rect 5436 8046 5454 8064
rect 5436 8064 5454 8082
rect 5436 8082 5454 8100
rect 5436 8100 5454 8118
rect 5436 8118 5454 8136
rect 5436 8136 5454 8154
rect 5436 8154 5454 8172
rect 5436 8172 5454 8190
rect 5436 8190 5454 8208
rect 5436 8208 5454 8226
rect 5436 8226 5454 8244
rect 5436 8244 5454 8262
rect 5436 8262 5454 8280
rect 5436 8280 5454 8298
rect 5436 8298 5454 8316
rect 5436 8316 5454 8334
rect 5436 8334 5454 8352
rect 5436 8352 5454 8370
rect 5436 8370 5454 8388
rect 5436 8388 5454 8406
rect 5436 8406 5454 8424
rect 5436 8424 5454 8442
rect 5436 8442 5454 8460
rect 5436 8460 5454 8478
rect 5454 486 5472 504
rect 5454 504 5472 522
rect 5454 522 5472 540
rect 5454 540 5472 558
rect 5454 558 5472 576
rect 5454 576 5472 594
rect 5454 594 5472 612
rect 5454 612 5472 630
rect 5454 630 5472 648
rect 5454 648 5472 666
rect 5454 666 5472 684
rect 5454 684 5472 702
rect 5454 702 5472 720
rect 5454 720 5472 738
rect 5454 738 5472 756
rect 5454 756 5472 774
rect 5454 774 5472 792
rect 5454 792 5472 810
rect 5454 810 5472 828
rect 5454 828 5472 846
rect 5454 846 5472 864
rect 5454 864 5472 882
rect 5454 882 5472 900
rect 5454 1044 5472 1062
rect 5454 1062 5472 1080
rect 5454 1080 5472 1098
rect 5454 1098 5472 1116
rect 5454 1116 5472 1134
rect 5454 1134 5472 1152
rect 5454 1152 5472 1170
rect 5454 1170 5472 1188
rect 5454 1188 5472 1206
rect 5454 1206 5472 1224
rect 5454 1224 5472 1242
rect 5454 1242 5472 1260
rect 5454 1260 5472 1278
rect 5454 1278 5472 1296
rect 5454 1296 5472 1314
rect 5454 1314 5472 1332
rect 5454 1332 5472 1350
rect 5454 1350 5472 1368
rect 5454 1368 5472 1386
rect 5454 1386 5472 1404
rect 5454 1404 5472 1422
rect 5454 1422 5472 1440
rect 5454 1440 5472 1458
rect 5454 1458 5472 1476
rect 5454 1476 5472 1494
rect 5454 1494 5472 1512
rect 5454 1512 5472 1530
rect 5454 1530 5472 1548
rect 5454 1548 5472 1566
rect 5454 1566 5472 1584
rect 5454 1584 5472 1602
rect 5454 1602 5472 1620
rect 5454 1620 5472 1638
rect 5454 1638 5472 1656
rect 5454 1656 5472 1674
rect 5454 1674 5472 1692
rect 5454 1692 5472 1710
rect 5454 1710 5472 1728
rect 5454 1728 5472 1746
rect 5454 1746 5472 1764
rect 5454 1764 5472 1782
rect 5454 1782 5472 1800
rect 5454 1800 5472 1818
rect 5454 1818 5472 1836
rect 5454 1836 5472 1854
rect 5454 1854 5472 1872
rect 5454 1872 5472 1890
rect 5454 1890 5472 1908
rect 5454 1908 5472 1926
rect 5454 1926 5472 1944
rect 5454 1944 5472 1962
rect 5454 1962 5472 1980
rect 5454 1980 5472 1998
rect 5454 1998 5472 2016
rect 5454 2016 5472 2034
rect 5454 2034 5472 2052
rect 5454 2052 5472 2070
rect 5454 2070 5472 2088
rect 5454 2088 5472 2106
rect 5454 2106 5472 2124
rect 5454 2124 5472 2142
rect 5454 2142 5472 2160
rect 5454 2160 5472 2178
rect 5454 2178 5472 2196
rect 5454 2196 5472 2214
rect 5454 2214 5472 2232
rect 5454 2232 5472 2250
rect 5454 2250 5472 2268
rect 5454 2268 5472 2286
rect 5454 2286 5472 2304
rect 5454 2304 5472 2322
rect 5454 2322 5472 2340
rect 5454 2340 5472 2358
rect 5454 2358 5472 2376
rect 5454 2376 5472 2394
rect 5454 2394 5472 2412
rect 5454 2412 5472 2430
rect 5454 2430 5472 2448
rect 5454 2448 5472 2466
rect 5454 2466 5472 2484
rect 5454 2484 5472 2502
rect 5454 2700 5472 2718
rect 5454 2718 5472 2736
rect 5454 2736 5472 2754
rect 5454 2754 5472 2772
rect 5454 2772 5472 2790
rect 5454 2790 5472 2808
rect 5454 2808 5472 2826
rect 5454 2826 5472 2844
rect 5454 2844 5472 2862
rect 5454 2862 5472 2880
rect 5454 2880 5472 2898
rect 5454 2898 5472 2916
rect 5454 2916 5472 2934
rect 5454 2934 5472 2952
rect 5454 2952 5472 2970
rect 5454 2970 5472 2988
rect 5454 2988 5472 3006
rect 5454 3006 5472 3024
rect 5454 3024 5472 3042
rect 5454 3042 5472 3060
rect 5454 3060 5472 3078
rect 5454 3078 5472 3096
rect 5454 3096 5472 3114
rect 5454 3114 5472 3132
rect 5454 3132 5472 3150
rect 5454 3150 5472 3168
rect 5454 3168 5472 3186
rect 5454 3186 5472 3204
rect 5454 3204 5472 3222
rect 5454 3222 5472 3240
rect 5454 3240 5472 3258
rect 5454 3258 5472 3276
rect 5454 3276 5472 3294
rect 5454 3294 5472 3312
rect 5454 3312 5472 3330
rect 5454 3330 5472 3348
rect 5454 3348 5472 3366
rect 5454 3366 5472 3384
rect 5454 3384 5472 3402
rect 5454 3402 5472 3420
rect 5454 3420 5472 3438
rect 5454 3438 5472 3456
rect 5454 3456 5472 3474
rect 5454 3474 5472 3492
rect 5454 3492 5472 3510
rect 5454 3510 5472 3528
rect 5454 3528 5472 3546
rect 5454 3546 5472 3564
rect 5454 3564 5472 3582
rect 5454 3582 5472 3600
rect 5454 3600 5472 3618
rect 5454 3618 5472 3636
rect 5454 3636 5472 3654
rect 5454 3654 5472 3672
rect 5454 3672 5472 3690
rect 5454 3690 5472 3708
rect 5454 3708 5472 3726
rect 5454 3726 5472 3744
rect 5454 3744 5472 3762
rect 5454 3762 5472 3780
rect 5454 3780 5472 3798
rect 5454 3798 5472 3816
rect 5454 3816 5472 3834
rect 5454 3834 5472 3852
rect 5454 3852 5472 3870
rect 5454 3870 5472 3888
rect 5454 3888 5472 3906
rect 5454 3906 5472 3924
rect 5454 3924 5472 3942
rect 5454 3942 5472 3960
rect 5454 3960 5472 3978
rect 5454 3978 5472 3996
rect 5454 3996 5472 4014
rect 5454 4014 5472 4032
rect 5454 4032 5472 4050
rect 5454 4050 5472 4068
rect 5454 4068 5472 4086
rect 5454 4086 5472 4104
rect 5454 4104 5472 4122
rect 5454 4122 5472 4140
rect 5454 4140 5472 4158
rect 5454 4158 5472 4176
rect 5454 4176 5472 4194
rect 5454 4194 5472 4212
rect 5454 4212 5472 4230
rect 5454 4230 5472 4248
rect 5454 4248 5472 4266
rect 5454 4266 5472 4284
rect 5454 4284 5472 4302
rect 5454 4302 5472 4320
rect 5454 4320 5472 4338
rect 5454 4338 5472 4356
rect 5454 4356 5472 4374
rect 5454 4374 5472 4392
rect 5454 4392 5472 4410
rect 5454 4410 5472 4428
rect 5454 4428 5472 4446
rect 5454 4446 5472 4464
rect 5454 4464 5472 4482
rect 5454 4482 5472 4500
rect 5454 4500 5472 4518
rect 5454 4518 5472 4536
rect 5454 4536 5472 4554
rect 5454 4554 5472 4572
rect 5454 4572 5472 4590
rect 5454 4590 5472 4608
rect 5454 4608 5472 4626
rect 5454 4626 5472 4644
rect 5454 4644 5472 4662
rect 5454 4662 5472 4680
rect 5454 4680 5472 4698
rect 5454 4698 5472 4716
rect 5454 4716 5472 4734
rect 5454 4734 5472 4752
rect 5454 4752 5472 4770
rect 5454 4770 5472 4788
rect 5454 4788 5472 4806
rect 5454 4806 5472 4824
rect 5454 4824 5472 4842
rect 5454 4842 5472 4860
rect 5454 5076 5472 5094
rect 5454 5094 5472 5112
rect 5454 5112 5472 5130
rect 5454 5130 5472 5148
rect 5454 5148 5472 5166
rect 5454 5166 5472 5184
rect 5454 5184 5472 5202
rect 5454 5202 5472 5220
rect 5454 5220 5472 5238
rect 5454 5238 5472 5256
rect 5454 5256 5472 5274
rect 5454 5274 5472 5292
rect 5454 5292 5472 5310
rect 5454 5310 5472 5328
rect 5454 5328 5472 5346
rect 5454 5346 5472 5364
rect 5454 5364 5472 5382
rect 5454 5382 5472 5400
rect 5454 5400 5472 5418
rect 5454 5418 5472 5436
rect 5454 5436 5472 5454
rect 5454 5454 5472 5472
rect 5454 5472 5472 5490
rect 5454 5490 5472 5508
rect 5454 5508 5472 5526
rect 5454 5526 5472 5544
rect 5454 5544 5472 5562
rect 5454 5562 5472 5580
rect 5454 5580 5472 5598
rect 5454 5598 5472 5616
rect 5454 5616 5472 5634
rect 5454 5634 5472 5652
rect 5454 5652 5472 5670
rect 5454 5670 5472 5688
rect 5454 5688 5472 5706
rect 5454 5706 5472 5724
rect 5454 5724 5472 5742
rect 5454 5742 5472 5760
rect 5454 5760 5472 5778
rect 5454 5778 5472 5796
rect 5454 5796 5472 5814
rect 5454 5814 5472 5832
rect 5454 5832 5472 5850
rect 5454 5850 5472 5868
rect 5454 5868 5472 5886
rect 5454 5886 5472 5904
rect 5454 5904 5472 5922
rect 5454 5922 5472 5940
rect 5454 5940 5472 5958
rect 5454 5958 5472 5976
rect 5454 5976 5472 5994
rect 5454 5994 5472 6012
rect 5454 6012 5472 6030
rect 5454 6030 5472 6048
rect 5454 6048 5472 6066
rect 5454 6066 5472 6084
rect 5454 6084 5472 6102
rect 5454 6102 5472 6120
rect 5454 6120 5472 6138
rect 5454 6138 5472 6156
rect 5454 6156 5472 6174
rect 5454 6174 5472 6192
rect 5454 6192 5472 6210
rect 5454 6210 5472 6228
rect 5454 6228 5472 6246
rect 5454 6246 5472 6264
rect 5454 6264 5472 6282
rect 5454 6282 5472 6300
rect 5454 6300 5472 6318
rect 5454 6318 5472 6336
rect 5454 6336 5472 6354
rect 5454 6354 5472 6372
rect 5454 6372 5472 6390
rect 5454 6390 5472 6408
rect 5454 6408 5472 6426
rect 5454 6426 5472 6444
rect 5454 6444 5472 6462
rect 5454 6462 5472 6480
rect 5454 6480 5472 6498
rect 5454 6498 5472 6516
rect 5454 6516 5472 6534
rect 5454 6534 5472 6552
rect 5454 6552 5472 6570
rect 5454 6570 5472 6588
rect 5454 6588 5472 6606
rect 5454 6606 5472 6624
rect 5454 6624 5472 6642
rect 5454 6642 5472 6660
rect 5454 6660 5472 6678
rect 5454 6678 5472 6696
rect 5454 6696 5472 6714
rect 5454 6714 5472 6732
rect 5454 6732 5472 6750
rect 5454 6750 5472 6768
rect 5454 6768 5472 6786
rect 5454 6786 5472 6804
rect 5454 6804 5472 6822
rect 5454 6822 5472 6840
rect 5454 6840 5472 6858
rect 5454 6858 5472 6876
rect 5454 6876 5472 6894
rect 5454 6894 5472 6912
rect 5454 6912 5472 6930
rect 5454 6930 5472 6948
rect 5454 6948 5472 6966
rect 5454 6966 5472 6984
rect 5454 6984 5472 7002
rect 5454 7002 5472 7020
rect 5454 7020 5472 7038
rect 5454 7038 5472 7056
rect 5454 7056 5472 7074
rect 5454 7074 5472 7092
rect 5454 7092 5472 7110
rect 5454 7110 5472 7128
rect 5454 7128 5472 7146
rect 5454 7146 5472 7164
rect 5454 7164 5472 7182
rect 5454 7182 5472 7200
rect 5454 7200 5472 7218
rect 5454 7218 5472 7236
rect 5454 7236 5472 7254
rect 5454 7254 5472 7272
rect 5454 7272 5472 7290
rect 5454 7290 5472 7308
rect 5454 7308 5472 7326
rect 5454 7326 5472 7344
rect 5454 7344 5472 7362
rect 5454 7362 5472 7380
rect 5454 7380 5472 7398
rect 5454 7398 5472 7416
rect 5454 7416 5472 7434
rect 5454 7434 5472 7452
rect 5454 7452 5472 7470
rect 5454 7470 5472 7488
rect 5454 7488 5472 7506
rect 5454 7506 5472 7524
rect 5454 7524 5472 7542
rect 5454 7542 5472 7560
rect 5454 7560 5472 7578
rect 5454 7578 5472 7596
rect 5454 7596 5472 7614
rect 5454 7614 5472 7632
rect 5454 7632 5472 7650
rect 5454 7650 5472 7668
rect 5454 7668 5472 7686
rect 5454 7686 5472 7704
rect 5454 7704 5472 7722
rect 5454 7722 5472 7740
rect 5454 7740 5472 7758
rect 5454 7758 5472 7776
rect 5454 7776 5472 7794
rect 5454 7794 5472 7812
rect 5454 7812 5472 7830
rect 5454 7830 5472 7848
rect 5454 7848 5472 7866
rect 5454 7866 5472 7884
rect 5454 7884 5472 7902
rect 5454 7902 5472 7920
rect 5454 7920 5472 7938
rect 5454 7938 5472 7956
rect 5454 7956 5472 7974
rect 5454 7974 5472 7992
rect 5454 7992 5472 8010
rect 5454 8010 5472 8028
rect 5454 8028 5472 8046
rect 5454 8046 5472 8064
rect 5454 8064 5472 8082
rect 5454 8082 5472 8100
rect 5454 8100 5472 8118
rect 5454 8118 5472 8136
rect 5454 8136 5472 8154
rect 5454 8154 5472 8172
rect 5454 8172 5472 8190
rect 5454 8190 5472 8208
rect 5454 8208 5472 8226
rect 5454 8226 5472 8244
rect 5454 8244 5472 8262
rect 5454 8262 5472 8280
rect 5454 8280 5472 8298
rect 5454 8298 5472 8316
rect 5454 8316 5472 8334
rect 5454 8334 5472 8352
rect 5454 8352 5472 8370
rect 5454 8370 5472 8388
rect 5454 8388 5472 8406
rect 5454 8406 5472 8424
rect 5454 8424 5472 8442
rect 5454 8442 5472 8460
rect 5454 8460 5472 8478
rect 5454 8478 5472 8496
rect 5472 504 5490 522
rect 5472 522 5490 540
rect 5472 540 5490 558
rect 5472 558 5490 576
rect 5472 576 5490 594
rect 5472 594 5490 612
rect 5472 612 5490 630
rect 5472 630 5490 648
rect 5472 648 5490 666
rect 5472 666 5490 684
rect 5472 684 5490 702
rect 5472 702 5490 720
rect 5472 720 5490 738
rect 5472 738 5490 756
rect 5472 756 5490 774
rect 5472 774 5490 792
rect 5472 792 5490 810
rect 5472 810 5490 828
rect 5472 828 5490 846
rect 5472 846 5490 864
rect 5472 864 5490 882
rect 5472 882 5490 900
rect 5472 900 5490 918
rect 5472 1044 5490 1062
rect 5472 1062 5490 1080
rect 5472 1080 5490 1098
rect 5472 1098 5490 1116
rect 5472 1116 5490 1134
rect 5472 1134 5490 1152
rect 5472 1152 5490 1170
rect 5472 1170 5490 1188
rect 5472 1188 5490 1206
rect 5472 1206 5490 1224
rect 5472 1224 5490 1242
rect 5472 1242 5490 1260
rect 5472 1260 5490 1278
rect 5472 1278 5490 1296
rect 5472 1296 5490 1314
rect 5472 1314 5490 1332
rect 5472 1332 5490 1350
rect 5472 1350 5490 1368
rect 5472 1368 5490 1386
rect 5472 1386 5490 1404
rect 5472 1404 5490 1422
rect 5472 1422 5490 1440
rect 5472 1440 5490 1458
rect 5472 1458 5490 1476
rect 5472 1476 5490 1494
rect 5472 1494 5490 1512
rect 5472 1512 5490 1530
rect 5472 1530 5490 1548
rect 5472 1548 5490 1566
rect 5472 1566 5490 1584
rect 5472 1584 5490 1602
rect 5472 1602 5490 1620
rect 5472 1620 5490 1638
rect 5472 1638 5490 1656
rect 5472 1656 5490 1674
rect 5472 1674 5490 1692
rect 5472 1692 5490 1710
rect 5472 1710 5490 1728
rect 5472 1728 5490 1746
rect 5472 1746 5490 1764
rect 5472 1764 5490 1782
rect 5472 1782 5490 1800
rect 5472 1800 5490 1818
rect 5472 1818 5490 1836
rect 5472 1836 5490 1854
rect 5472 1854 5490 1872
rect 5472 1872 5490 1890
rect 5472 1890 5490 1908
rect 5472 1908 5490 1926
rect 5472 1926 5490 1944
rect 5472 1944 5490 1962
rect 5472 1962 5490 1980
rect 5472 1980 5490 1998
rect 5472 1998 5490 2016
rect 5472 2016 5490 2034
rect 5472 2034 5490 2052
rect 5472 2052 5490 2070
rect 5472 2070 5490 2088
rect 5472 2088 5490 2106
rect 5472 2106 5490 2124
rect 5472 2124 5490 2142
rect 5472 2142 5490 2160
rect 5472 2160 5490 2178
rect 5472 2178 5490 2196
rect 5472 2196 5490 2214
rect 5472 2214 5490 2232
rect 5472 2232 5490 2250
rect 5472 2250 5490 2268
rect 5472 2268 5490 2286
rect 5472 2286 5490 2304
rect 5472 2304 5490 2322
rect 5472 2322 5490 2340
rect 5472 2340 5490 2358
rect 5472 2358 5490 2376
rect 5472 2376 5490 2394
rect 5472 2394 5490 2412
rect 5472 2412 5490 2430
rect 5472 2430 5490 2448
rect 5472 2448 5490 2466
rect 5472 2466 5490 2484
rect 5472 2484 5490 2502
rect 5472 2700 5490 2718
rect 5472 2718 5490 2736
rect 5472 2736 5490 2754
rect 5472 2754 5490 2772
rect 5472 2772 5490 2790
rect 5472 2790 5490 2808
rect 5472 2808 5490 2826
rect 5472 2826 5490 2844
rect 5472 2844 5490 2862
rect 5472 2862 5490 2880
rect 5472 2880 5490 2898
rect 5472 2898 5490 2916
rect 5472 2916 5490 2934
rect 5472 2934 5490 2952
rect 5472 2952 5490 2970
rect 5472 2970 5490 2988
rect 5472 2988 5490 3006
rect 5472 3006 5490 3024
rect 5472 3024 5490 3042
rect 5472 3042 5490 3060
rect 5472 3060 5490 3078
rect 5472 3078 5490 3096
rect 5472 3096 5490 3114
rect 5472 3114 5490 3132
rect 5472 3132 5490 3150
rect 5472 3150 5490 3168
rect 5472 3168 5490 3186
rect 5472 3186 5490 3204
rect 5472 3204 5490 3222
rect 5472 3222 5490 3240
rect 5472 3240 5490 3258
rect 5472 3258 5490 3276
rect 5472 3276 5490 3294
rect 5472 3294 5490 3312
rect 5472 3312 5490 3330
rect 5472 3330 5490 3348
rect 5472 3348 5490 3366
rect 5472 3366 5490 3384
rect 5472 3384 5490 3402
rect 5472 3402 5490 3420
rect 5472 3420 5490 3438
rect 5472 3438 5490 3456
rect 5472 3456 5490 3474
rect 5472 3474 5490 3492
rect 5472 3492 5490 3510
rect 5472 3510 5490 3528
rect 5472 3528 5490 3546
rect 5472 3546 5490 3564
rect 5472 3564 5490 3582
rect 5472 3582 5490 3600
rect 5472 3600 5490 3618
rect 5472 3618 5490 3636
rect 5472 3636 5490 3654
rect 5472 3654 5490 3672
rect 5472 3672 5490 3690
rect 5472 3690 5490 3708
rect 5472 3708 5490 3726
rect 5472 3726 5490 3744
rect 5472 3744 5490 3762
rect 5472 3762 5490 3780
rect 5472 3780 5490 3798
rect 5472 3798 5490 3816
rect 5472 3816 5490 3834
rect 5472 3834 5490 3852
rect 5472 3852 5490 3870
rect 5472 3870 5490 3888
rect 5472 3888 5490 3906
rect 5472 3906 5490 3924
rect 5472 3924 5490 3942
rect 5472 3942 5490 3960
rect 5472 3960 5490 3978
rect 5472 3978 5490 3996
rect 5472 3996 5490 4014
rect 5472 4014 5490 4032
rect 5472 4032 5490 4050
rect 5472 4050 5490 4068
rect 5472 4068 5490 4086
rect 5472 4086 5490 4104
rect 5472 4104 5490 4122
rect 5472 4122 5490 4140
rect 5472 4140 5490 4158
rect 5472 4158 5490 4176
rect 5472 4176 5490 4194
rect 5472 4194 5490 4212
rect 5472 4212 5490 4230
rect 5472 4230 5490 4248
rect 5472 4248 5490 4266
rect 5472 4266 5490 4284
rect 5472 4284 5490 4302
rect 5472 4302 5490 4320
rect 5472 4320 5490 4338
rect 5472 4338 5490 4356
rect 5472 4356 5490 4374
rect 5472 4374 5490 4392
rect 5472 4392 5490 4410
rect 5472 4410 5490 4428
rect 5472 4428 5490 4446
rect 5472 4446 5490 4464
rect 5472 4464 5490 4482
rect 5472 4482 5490 4500
rect 5472 4500 5490 4518
rect 5472 4518 5490 4536
rect 5472 4536 5490 4554
rect 5472 4554 5490 4572
rect 5472 4572 5490 4590
rect 5472 4590 5490 4608
rect 5472 4608 5490 4626
rect 5472 4626 5490 4644
rect 5472 4644 5490 4662
rect 5472 4662 5490 4680
rect 5472 4680 5490 4698
rect 5472 4698 5490 4716
rect 5472 4716 5490 4734
rect 5472 4734 5490 4752
rect 5472 4752 5490 4770
rect 5472 4770 5490 4788
rect 5472 4788 5490 4806
rect 5472 4806 5490 4824
rect 5472 4824 5490 4842
rect 5472 4842 5490 4860
rect 5472 4860 5490 4878
rect 5472 5094 5490 5112
rect 5472 5112 5490 5130
rect 5472 5130 5490 5148
rect 5472 5148 5490 5166
rect 5472 5166 5490 5184
rect 5472 5184 5490 5202
rect 5472 5202 5490 5220
rect 5472 5220 5490 5238
rect 5472 5238 5490 5256
rect 5472 5256 5490 5274
rect 5472 5274 5490 5292
rect 5472 5292 5490 5310
rect 5472 5310 5490 5328
rect 5472 5328 5490 5346
rect 5472 5346 5490 5364
rect 5472 5364 5490 5382
rect 5472 5382 5490 5400
rect 5472 5400 5490 5418
rect 5472 5418 5490 5436
rect 5472 5436 5490 5454
rect 5472 5454 5490 5472
rect 5472 5472 5490 5490
rect 5472 5490 5490 5508
rect 5472 5508 5490 5526
rect 5472 5526 5490 5544
rect 5472 5544 5490 5562
rect 5472 5562 5490 5580
rect 5472 5580 5490 5598
rect 5472 5598 5490 5616
rect 5472 5616 5490 5634
rect 5472 5634 5490 5652
rect 5472 5652 5490 5670
rect 5472 5670 5490 5688
rect 5472 5688 5490 5706
rect 5472 5706 5490 5724
rect 5472 5724 5490 5742
rect 5472 5742 5490 5760
rect 5472 5760 5490 5778
rect 5472 5778 5490 5796
rect 5472 5796 5490 5814
rect 5472 5814 5490 5832
rect 5472 5832 5490 5850
rect 5472 5850 5490 5868
rect 5472 5868 5490 5886
rect 5472 5886 5490 5904
rect 5472 5904 5490 5922
rect 5472 5922 5490 5940
rect 5472 5940 5490 5958
rect 5472 5958 5490 5976
rect 5472 5976 5490 5994
rect 5472 5994 5490 6012
rect 5472 6012 5490 6030
rect 5472 6030 5490 6048
rect 5472 6048 5490 6066
rect 5472 6066 5490 6084
rect 5472 6084 5490 6102
rect 5472 6102 5490 6120
rect 5472 6120 5490 6138
rect 5472 6138 5490 6156
rect 5472 6156 5490 6174
rect 5472 6174 5490 6192
rect 5472 6192 5490 6210
rect 5472 6210 5490 6228
rect 5472 6228 5490 6246
rect 5472 6246 5490 6264
rect 5472 6264 5490 6282
rect 5472 6282 5490 6300
rect 5472 6300 5490 6318
rect 5472 6318 5490 6336
rect 5472 6336 5490 6354
rect 5472 6354 5490 6372
rect 5472 6372 5490 6390
rect 5472 6390 5490 6408
rect 5472 6408 5490 6426
rect 5472 6426 5490 6444
rect 5472 6444 5490 6462
rect 5472 6462 5490 6480
rect 5472 6480 5490 6498
rect 5472 6498 5490 6516
rect 5472 6516 5490 6534
rect 5472 6534 5490 6552
rect 5472 6552 5490 6570
rect 5472 6570 5490 6588
rect 5472 6588 5490 6606
rect 5472 6606 5490 6624
rect 5472 6624 5490 6642
rect 5472 6642 5490 6660
rect 5472 6660 5490 6678
rect 5472 6678 5490 6696
rect 5472 6696 5490 6714
rect 5472 6714 5490 6732
rect 5472 6732 5490 6750
rect 5472 6750 5490 6768
rect 5472 6768 5490 6786
rect 5472 6786 5490 6804
rect 5472 6804 5490 6822
rect 5472 6822 5490 6840
rect 5472 6840 5490 6858
rect 5472 6858 5490 6876
rect 5472 6876 5490 6894
rect 5472 6894 5490 6912
rect 5472 6912 5490 6930
rect 5472 6930 5490 6948
rect 5472 6948 5490 6966
rect 5472 6966 5490 6984
rect 5472 6984 5490 7002
rect 5472 7002 5490 7020
rect 5472 7020 5490 7038
rect 5472 7038 5490 7056
rect 5472 7056 5490 7074
rect 5472 7074 5490 7092
rect 5472 7092 5490 7110
rect 5472 7110 5490 7128
rect 5472 7128 5490 7146
rect 5472 7146 5490 7164
rect 5472 7164 5490 7182
rect 5472 7182 5490 7200
rect 5472 7200 5490 7218
rect 5472 7218 5490 7236
rect 5472 7236 5490 7254
rect 5472 7254 5490 7272
rect 5472 7272 5490 7290
rect 5472 7290 5490 7308
rect 5472 7308 5490 7326
rect 5472 7326 5490 7344
rect 5472 7344 5490 7362
rect 5472 7362 5490 7380
rect 5472 7380 5490 7398
rect 5472 7398 5490 7416
rect 5472 7416 5490 7434
rect 5472 7434 5490 7452
rect 5472 7452 5490 7470
rect 5472 7470 5490 7488
rect 5472 7488 5490 7506
rect 5472 7506 5490 7524
rect 5472 7524 5490 7542
rect 5472 7542 5490 7560
rect 5472 7560 5490 7578
rect 5472 7578 5490 7596
rect 5472 7596 5490 7614
rect 5472 7614 5490 7632
rect 5472 7632 5490 7650
rect 5472 7650 5490 7668
rect 5472 7668 5490 7686
rect 5472 7686 5490 7704
rect 5472 7704 5490 7722
rect 5472 7722 5490 7740
rect 5472 7740 5490 7758
rect 5472 7758 5490 7776
rect 5472 7776 5490 7794
rect 5472 7794 5490 7812
rect 5472 7812 5490 7830
rect 5472 7830 5490 7848
rect 5472 7848 5490 7866
rect 5472 7866 5490 7884
rect 5472 7884 5490 7902
rect 5472 7902 5490 7920
rect 5472 7920 5490 7938
rect 5472 7938 5490 7956
rect 5472 7956 5490 7974
rect 5472 7974 5490 7992
rect 5472 7992 5490 8010
rect 5472 8010 5490 8028
rect 5472 8028 5490 8046
rect 5472 8046 5490 8064
rect 5472 8064 5490 8082
rect 5472 8082 5490 8100
rect 5472 8100 5490 8118
rect 5472 8118 5490 8136
rect 5472 8136 5490 8154
rect 5472 8154 5490 8172
rect 5472 8172 5490 8190
rect 5472 8190 5490 8208
rect 5472 8208 5490 8226
rect 5472 8226 5490 8244
rect 5472 8244 5490 8262
rect 5472 8262 5490 8280
rect 5472 8280 5490 8298
rect 5472 8298 5490 8316
rect 5472 8316 5490 8334
rect 5472 8334 5490 8352
rect 5472 8352 5490 8370
rect 5472 8370 5490 8388
rect 5472 8388 5490 8406
rect 5472 8406 5490 8424
rect 5472 8424 5490 8442
rect 5472 8442 5490 8460
rect 5472 8460 5490 8478
rect 5472 8478 5490 8496
rect 5472 8496 5490 8514
rect 5472 8514 5490 8532
rect 5490 522 5508 540
rect 5490 540 5508 558
rect 5490 558 5508 576
rect 5490 576 5508 594
rect 5490 594 5508 612
rect 5490 612 5508 630
rect 5490 630 5508 648
rect 5490 648 5508 666
rect 5490 666 5508 684
rect 5490 684 5508 702
rect 5490 702 5508 720
rect 5490 720 5508 738
rect 5490 738 5508 756
rect 5490 756 5508 774
rect 5490 774 5508 792
rect 5490 792 5508 810
rect 5490 810 5508 828
rect 5490 828 5508 846
rect 5490 846 5508 864
rect 5490 864 5508 882
rect 5490 882 5508 900
rect 5490 900 5508 918
rect 5490 1044 5508 1062
rect 5490 1062 5508 1080
rect 5490 1080 5508 1098
rect 5490 1098 5508 1116
rect 5490 1116 5508 1134
rect 5490 1134 5508 1152
rect 5490 1152 5508 1170
rect 5490 1170 5508 1188
rect 5490 1188 5508 1206
rect 5490 1206 5508 1224
rect 5490 1224 5508 1242
rect 5490 1242 5508 1260
rect 5490 1260 5508 1278
rect 5490 1278 5508 1296
rect 5490 1296 5508 1314
rect 5490 1314 5508 1332
rect 5490 1332 5508 1350
rect 5490 1350 5508 1368
rect 5490 1368 5508 1386
rect 5490 1386 5508 1404
rect 5490 1404 5508 1422
rect 5490 1422 5508 1440
rect 5490 1440 5508 1458
rect 5490 1458 5508 1476
rect 5490 1476 5508 1494
rect 5490 1494 5508 1512
rect 5490 1512 5508 1530
rect 5490 1530 5508 1548
rect 5490 1548 5508 1566
rect 5490 1566 5508 1584
rect 5490 1584 5508 1602
rect 5490 1602 5508 1620
rect 5490 1620 5508 1638
rect 5490 1638 5508 1656
rect 5490 1656 5508 1674
rect 5490 1674 5508 1692
rect 5490 1692 5508 1710
rect 5490 1710 5508 1728
rect 5490 1728 5508 1746
rect 5490 1746 5508 1764
rect 5490 1764 5508 1782
rect 5490 1782 5508 1800
rect 5490 1800 5508 1818
rect 5490 1818 5508 1836
rect 5490 1836 5508 1854
rect 5490 1854 5508 1872
rect 5490 1872 5508 1890
rect 5490 1890 5508 1908
rect 5490 1908 5508 1926
rect 5490 1926 5508 1944
rect 5490 1944 5508 1962
rect 5490 1962 5508 1980
rect 5490 1980 5508 1998
rect 5490 1998 5508 2016
rect 5490 2016 5508 2034
rect 5490 2034 5508 2052
rect 5490 2052 5508 2070
rect 5490 2070 5508 2088
rect 5490 2088 5508 2106
rect 5490 2106 5508 2124
rect 5490 2124 5508 2142
rect 5490 2142 5508 2160
rect 5490 2160 5508 2178
rect 5490 2178 5508 2196
rect 5490 2196 5508 2214
rect 5490 2214 5508 2232
rect 5490 2232 5508 2250
rect 5490 2250 5508 2268
rect 5490 2268 5508 2286
rect 5490 2286 5508 2304
rect 5490 2304 5508 2322
rect 5490 2322 5508 2340
rect 5490 2340 5508 2358
rect 5490 2358 5508 2376
rect 5490 2376 5508 2394
rect 5490 2394 5508 2412
rect 5490 2412 5508 2430
rect 5490 2430 5508 2448
rect 5490 2448 5508 2466
rect 5490 2466 5508 2484
rect 5490 2484 5508 2502
rect 5490 2502 5508 2520
rect 5490 2718 5508 2736
rect 5490 2736 5508 2754
rect 5490 2754 5508 2772
rect 5490 2772 5508 2790
rect 5490 2790 5508 2808
rect 5490 2808 5508 2826
rect 5490 2826 5508 2844
rect 5490 2844 5508 2862
rect 5490 2862 5508 2880
rect 5490 2880 5508 2898
rect 5490 2898 5508 2916
rect 5490 2916 5508 2934
rect 5490 2934 5508 2952
rect 5490 2952 5508 2970
rect 5490 2970 5508 2988
rect 5490 2988 5508 3006
rect 5490 3006 5508 3024
rect 5490 3024 5508 3042
rect 5490 3042 5508 3060
rect 5490 3060 5508 3078
rect 5490 3078 5508 3096
rect 5490 3096 5508 3114
rect 5490 3114 5508 3132
rect 5490 3132 5508 3150
rect 5490 3150 5508 3168
rect 5490 3168 5508 3186
rect 5490 3186 5508 3204
rect 5490 3204 5508 3222
rect 5490 3222 5508 3240
rect 5490 3240 5508 3258
rect 5490 3258 5508 3276
rect 5490 3276 5508 3294
rect 5490 3294 5508 3312
rect 5490 3312 5508 3330
rect 5490 3330 5508 3348
rect 5490 3348 5508 3366
rect 5490 3366 5508 3384
rect 5490 3384 5508 3402
rect 5490 3402 5508 3420
rect 5490 3420 5508 3438
rect 5490 3438 5508 3456
rect 5490 3456 5508 3474
rect 5490 3474 5508 3492
rect 5490 3492 5508 3510
rect 5490 3510 5508 3528
rect 5490 3528 5508 3546
rect 5490 3546 5508 3564
rect 5490 3564 5508 3582
rect 5490 3582 5508 3600
rect 5490 3600 5508 3618
rect 5490 3618 5508 3636
rect 5490 3636 5508 3654
rect 5490 3654 5508 3672
rect 5490 3672 5508 3690
rect 5490 3690 5508 3708
rect 5490 3708 5508 3726
rect 5490 3726 5508 3744
rect 5490 3744 5508 3762
rect 5490 3762 5508 3780
rect 5490 3780 5508 3798
rect 5490 3798 5508 3816
rect 5490 3816 5508 3834
rect 5490 3834 5508 3852
rect 5490 3852 5508 3870
rect 5490 3870 5508 3888
rect 5490 3888 5508 3906
rect 5490 3906 5508 3924
rect 5490 3924 5508 3942
rect 5490 3942 5508 3960
rect 5490 3960 5508 3978
rect 5490 3978 5508 3996
rect 5490 3996 5508 4014
rect 5490 4014 5508 4032
rect 5490 4032 5508 4050
rect 5490 4050 5508 4068
rect 5490 4068 5508 4086
rect 5490 4086 5508 4104
rect 5490 4104 5508 4122
rect 5490 4122 5508 4140
rect 5490 4140 5508 4158
rect 5490 4158 5508 4176
rect 5490 4176 5508 4194
rect 5490 4194 5508 4212
rect 5490 4212 5508 4230
rect 5490 4230 5508 4248
rect 5490 4248 5508 4266
rect 5490 4266 5508 4284
rect 5490 4284 5508 4302
rect 5490 4302 5508 4320
rect 5490 4320 5508 4338
rect 5490 4338 5508 4356
rect 5490 4356 5508 4374
rect 5490 4374 5508 4392
rect 5490 4392 5508 4410
rect 5490 4410 5508 4428
rect 5490 4428 5508 4446
rect 5490 4446 5508 4464
rect 5490 4464 5508 4482
rect 5490 4482 5508 4500
rect 5490 4500 5508 4518
rect 5490 4518 5508 4536
rect 5490 4536 5508 4554
rect 5490 4554 5508 4572
rect 5490 4572 5508 4590
rect 5490 4590 5508 4608
rect 5490 4608 5508 4626
rect 5490 4626 5508 4644
rect 5490 4644 5508 4662
rect 5490 4662 5508 4680
rect 5490 4680 5508 4698
rect 5490 4698 5508 4716
rect 5490 4716 5508 4734
rect 5490 4734 5508 4752
rect 5490 4752 5508 4770
rect 5490 4770 5508 4788
rect 5490 4788 5508 4806
rect 5490 4806 5508 4824
rect 5490 4824 5508 4842
rect 5490 4842 5508 4860
rect 5490 4860 5508 4878
rect 5490 4878 5508 4896
rect 5490 5112 5508 5130
rect 5490 5130 5508 5148
rect 5490 5148 5508 5166
rect 5490 5166 5508 5184
rect 5490 5184 5508 5202
rect 5490 5202 5508 5220
rect 5490 5220 5508 5238
rect 5490 5238 5508 5256
rect 5490 5256 5508 5274
rect 5490 5274 5508 5292
rect 5490 5292 5508 5310
rect 5490 5310 5508 5328
rect 5490 5328 5508 5346
rect 5490 5346 5508 5364
rect 5490 5364 5508 5382
rect 5490 5382 5508 5400
rect 5490 5400 5508 5418
rect 5490 5418 5508 5436
rect 5490 5436 5508 5454
rect 5490 5454 5508 5472
rect 5490 5472 5508 5490
rect 5490 5490 5508 5508
rect 5490 5508 5508 5526
rect 5490 5526 5508 5544
rect 5490 5544 5508 5562
rect 5490 5562 5508 5580
rect 5490 5580 5508 5598
rect 5490 5598 5508 5616
rect 5490 5616 5508 5634
rect 5490 5634 5508 5652
rect 5490 5652 5508 5670
rect 5490 5670 5508 5688
rect 5490 5688 5508 5706
rect 5490 5706 5508 5724
rect 5490 5724 5508 5742
rect 5490 5742 5508 5760
rect 5490 5760 5508 5778
rect 5490 5778 5508 5796
rect 5490 5796 5508 5814
rect 5490 5814 5508 5832
rect 5490 5832 5508 5850
rect 5490 5850 5508 5868
rect 5490 5868 5508 5886
rect 5490 5886 5508 5904
rect 5490 5904 5508 5922
rect 5490 5922 5508 5940
rect 5490 5940 5508 5958
rect 5490 5958 5508 5976
rect 5490 5976 5508 5994
rect 5490 5994 5508 6012
rect 5490 6012 5508 6030
rect 5490 6030 5508 6048
rect 5490 6048 5508 6066
rect 5490 6066 5508 6084
rect 5490 6084 5508 6102
rect 5490 6102 5508 6120
rect 5490 6120 5508 6138
rect 5490 6138 5508 6156
rect 5490 6156 5508 6174
rect 5490 6174 5508 6192
rect 5490 6192 5508 6210
rect 5490 6210 5508 6228
rect 5490 6228 5508 6246
rect 5490 6246 5508 6264
rect 5490 6264 5508 6282
rect 5490 6282 5508 6300
rect 5490 6300 5508 6318
rect 5490 6318 5508 6336
rect 5490 6336 5508 6354
rect 5490 6354 5508 6372
rect 5490 6372 5508 6390
rect 5490 6390 5508 6408
rect 5490 6408 5508 6426
rect 5490 6426 5508 6444
rect 5490 6444 5508 6462
rect 5490 6462 5508 6480
rect 5490 6480 5508 6498
rect 5490 6498 5508 6516
rect 5490 6516 5508 6534
rect 5490 6534 5508 6552
rect 5490 6552 5508 6570
rect 5490 6570 5508 6588
rect 5490 6588 5508 6606
rect 5490 6606 5508 6624
rect 5490 6624 5508 6642
rect 5490 6642 5508 6660
rect 5490 6660 5508 6678
rect 5490 6678 5508 6696
rect 5490 6696 5508 6714
rect 5490 6714 5508 6732
rect 5490 6732 5508 6750
rect 5490 6750 5508 6768
rect 5490 6768 5508 6786
rect 5490 6786 5508 6804
rect 5490 6804 5508 6822
rect 5490 6822 5508 6840
rect 5490 6840 5508 6858
rect 5490 6858 5508 6876
rect 5490 6876 5508 6894
rect 5490 6894 5508 6912
rect 5490 6912 5508 6930
rect 5490 6930 5508 6948
rect 5490 6948 5508 6966
rect 5490 6966 5508 6984
rect 5490 6984 5508 7002
rect 5490 7002 5508 7020
rect 5490 7020 5508 7038
rect 5490 7038 5508 7056
rect 5490 7056 5508 7074
rect 5490 7074 5508 7092
rect 5490 7092 5508 7110
rect 5490 7110 5508 7128
rect 5490 7128 5508 7146
rect 5490 7146 5508 7164
rect 5490 7164 5508 7182
rect 5490 7182 5508 7200
rect 5490 7200 5508 7218
rect 5490 7218 5508 7236
rect 5490 7236 5508 7254
rect 5490 7254 5508 7272
rect 5490 7272 5508 7290
rect 5490 7290 5508 7308
rect 5490 7308 5508 7326
rect 5490 7326 5508 7344
rect 5490 7344 5508 7362
rect 5490 7362 5508 7380
rect 5490 7380 5508 7398
rect 5490 7398 5508 7416
rect 5490 7416 5508 7434
rect 5490 7434 5508 7452
rect 5490 7452 5508 7470
rect 5490 7470 5508 7488
rect 5490 7488 5508 7506
rect 5490 7506 5508 7524
rect 5490 7524 5508 7542
rect 5490 7542 5508 7560
rect 5490 7560 5508 7578
rect 5490 7578 5508 7596
rect 5490 7596 5508 7614
rect 5490 7614 5508 7632
rect 5490 7632 5508 7650
rect 5490 7650 5508 7668
rect 5490 7668 5508 7686
rect 5490 7686 5508 7704
rect 5490 7704 5508 7722
rect 5490 7722 5508 7740
rect 5490 7740 5508 7758
rect 5490 7758 5508 7776
rect 5490 7776 5508 7794
rect 5490 7794 5508 7812
rect 5490 7812 5508 7830
rect 5490 7830 5508 7848
rect 5490 7848 5508 7866
rect 5490 7866 5508 7884
rect 5490 7884 5508 7902
rect 5490 7902 5508 7920
rect 5490 7920 5508 7938
rect 5490 7938 5508 7956
rect 5490 7956 5508 7974
rect 5490 7974 5508 7992
rect 5490 7992 5508 8010
rect 5490 8010 5508 8028
rect 5490 8028 5508 8046
rect 5490 8046 5508 8064
rect 5490 8064 5508 8082
rect 5490 8082 5508 8100
rect 5490 8100 5508 8118
rect 5490 8118 5508 8136
rect 5490 8136 5508 8154
rect 5490 8154 5508 8172
rect 5490 8172 5508 8190
rect 5490 8190 5508 8208
rect 5490 8208 5508 8226
rect 5490 8226 5508 8244
rect 5490 8244 5508 8262
rect 5490 8262 5508 8280
rect 5490 8280 5508 8298
rect 5490 8298 5508 8316
rect 5490 8316 5508 8334
rect 5490 8334 5508 8352
rect 5490 8352 5508 8370
rect 5490 8370 5508 8388
rect 5490 8388 5508 8406
rect 5490 8406 5508 8424
rect 5490 8424 5508 8442
rect 5490 8442 5508 8460
rect 5490 8460 5508 8478
rect 5490 8478 5508 8496
rect 5490 8496 5508 8514
rect 5490 8514 5508 8532
rect 5490 8532 5508 8550
rect 5508 522 5526 540
rect 5508 540 5526 558
rect 5508 558 5526 576
rect 5508 576 5526 594
rect 5508 594 5526 612
rect 5508 612 5526 630
rect 5508 630 5526 648
rect 5508 648 5526 666
rect 5508 666 5526 684
rect 5508 684 5526 702
rect 5508 702 5526 720
rect 5508 720 5526 738
rect 5508 738 5526 756
rect 5508 756 5526 774
rect 5508 774 5526 792
rect 5508 792 5526 810
rect 5508 810 5526 828
rect 5508 828 5526 846
rect 5508 846 5526 864
rect 5508 864 5526 882
rect 5508 882 5526 900
rect 5508 900 5526 918
rect 5508 1062 5526 1080
rect 5508 1080 5526 1098
rect 5508 1098 5526 1116
rect 5508 1116 5526 1134
rect 5508 1134 5526 1152
rect 5508 1152 5526 1170
rect 5508 1170 5526 1188
rect 5508 1188 5526 1206
rect 5508 1206 5526 1224
rect 5508 1224 5526 1242
rect 5508 1242 5526 1260
rect 5508 1260 5526 1278
rect 5508 1278 5526 1296
rect 5508 1296 5526 1314
rect 5508 1314 5526 1332
rect 5508 1332 5526 1350
rect 5508 1350 5526 1368
rect 5508 1368 5526 1386
rect 5508 1386 5526 1404
rect 5508 1404 5526 1422
rect 5508 1422 5526 1440
rect 5508 1440 5526 1458
rect 5508 1458 5526 1476
rect 5508 1476 5526 1494
rect 5508 1494 5526 1512
rect 5508 1512 5526 1530
rect 5508 1530 5526 1548
rect 5508 1548 5526 1566
rect 5508 1566 5526 1584
rect 5508 1584 5526 1602
rect 5508 1602 5526 1620
rect 5508 1620 5526 1638
rect 5508 1638 5526 1656
rect 5508 1656 5526 1674
rect 5508 1674 5526 1692
rect 5508 1692 5526 1710
rect 5508 1710 5526 1728
rect 5508 1728 5526 1746
rect 5508 1746 5526 1764
rect 5508 1764 5526 1782
rect 5508 1782 5526 1800
rect 5508 1800 5526 1818
rect 5508 1818 5526 1836
rect 5508 1836 5526 1854
rect 5508 1854 5526 1872
rect 5508 1872 5526 1890
rect 5508 1890 5526 1908
rect 5508 1908 5526 1926
rect 5508 1926 5526 1944
rect 5508 1944 5526 1962
rect 5508 1962 5526 1980
rect 5508 1980 5526 1998
rect 5508 1998 5526 2016
rect 5508 2016 5526 2034
rect 5508 2034 5526 2052
rect 5508 2052 5526 2070
rect 5508 2070 5526 2088
rect 5508 2088 5526 2106
rect 5508 2106 5526 2124
rect 5508 2124 5526 2142
rect 5508 2142 5526 2160
rect 5508 2160 5526 2178
rect 5508 2178 5526 2196
rect 5508 2196 5526 2214
rect 5508 2214 5526 2232
rect 5508 2232 5526 2250
rect 5508 2250 5526 2268
rect 5508 2268 5526 2286
rect 5508 2286 5526 2304
rect 5508 2304 5526 2322
rect 5508 2322 5526 2340
rect 5508 2340 5526 2358
rect 5508 2358 5526 2376
rect 5508 2376 5526 2394
rect 5508 2394 5526 2412
rect 5508 2412 5526 2430
rect 5508 2430 5526 2448
rect 5508 2448 5526 2466
rect 5508 2466 5526 2484
rect 5508 2484 5526 2502
rect 5508 2502 5526 2520
rect 5508 2736 5526 2754
rect 5508 2754 5526 2772
rect 5508 2772 5526 2790
rect 5508 2790 5526 2808
rect 5508 2808 5526 2826
rect 5508 2826 5526 2844
rect 5508 2844 5526 2862
rect 5508 2862 5526 2880
rect 5508 2880 5526 2898
rect 5508 2898 5526 2916
rect 5508 2916 5526 2934
rect 5508 2934 5526 2952
rect 5508 2952 5526 2970
rect 5508 2970 5526 2988
rect 5508 2988 5526 3006
rect 5508 3006 5526 3024
rect 5508 3024 5526 3042
rect 5508 3042 5526 3060
rect 5508 3060 5526 3078
rect 5508 3078 5526 3096
rect 5508 3096 5526 3114
rect 5508 3114 5526 3132
rect 5508 3132 5526 3150
rect 5508 3150 5526 3168
rect 5508 3168 5526 3186
rect 5508 3186 5526 3204
rect 5508 3204 5526 3222
rect 5508 3222 5526 3240
rect 5508 3240 5526 3258
rect 5508 3258 5526 3276
rect 5508 3276 5526 3294
rect 5508 3294 5526 3312
rect 5508 3312 5526 3330
rect 5508 3330 5526 3348
rect 5508 3348 5526 3366
rect 5508 3366 5526 3384
rect 5508 3384 5526 3402
rect 5508 3402 5526 3420
rect 5508 3420 5526 3438
rect 5508 3438 5526 3456
rect 5508 3456 5526 3474
rect 5508 3474 5526 3492
rect 5508 3492 5526 3510
rect 5508 3510 5526 3528
rect 5508 3528 5526 3546
rect 5508 3546 5526 3564
rect 5508 3564 5526 3582
rect 5508 3582 5526 3600
rect 5508 3600 5526 3618
rect 5508 3618 5526 3636
rect 5508 3636 5526 3654
rect 5508 3654 5526 3672
rect 5508 3672 5526 3690
rect 5508 3690 5526 3708
rect 5508 3708 5526 3726
rect 5508 3726 5526 3744
rect 5508 3744 5526 3762
rect 5508 3762 5526 3780
rect 5508 3780 5526 3798
rect 5508 3798 5526 3816
rect 5508 3816 5526 3834
rect 5508 3834 5526 3852
rect 5508 3852 5526 3870
rect 5508 3870 5526 3888
rect 5508 3888 5526 3906
rect 5508 3906 5526 3924
rect 5508 3924 5526 3942
rect 5508 3942 5526 3960
rect 5508 3960 5526 3978
rect 5508 3978 5526 3996
rect 5508 3996 5526 4014
rect 5508 4014 5526 4032
rect 5508 4032 5526 4050
rect 5508 4050 5526 4068
rect 5508 4068 5526 4086
rect 5508 4086 5526 4104
rect 5508 4104 5526 4122
rect 5508 4122 5526 4140
rect 5508 4140 5526 4158
rect 5508 4158 5526 4176
rect 5508 4176 5526 4194
rect 5508 4194 5526 4212
rect 5508 4212 5526 4230
rect 5508 4230 5526 4248
rect 5508 4248 5526 4266
rect 5508 4266 5526 4284
rect 5508 4284 5526 4302
rect 5508 4302 5526 4320
rect 5508 4320 5526 4338
rect 5508 4338 5526 4356
rect 5508 4356 5526 4374
rect 5508 4374 5526 4392
rect 5508 4392 5526 4410
rect 5508 4410 5526 4428
rect 5508 4428 5526 4446
rect 5508 4446 5526 4464
rect 5508 4464 5526 4482
rect 5508 4482 5526 4500
rect 5508 4500 5526 4518
rect 5508 4518 5526 4536
rect 5508 4536 5526 4554
rect 5508 4554 5526 4572
rect 5508 4572 5526 4590
rect 5508 4590 5526 4608
rect 5508 4608 5526 4626
rect 5508 4626 5526 4644
rect 5508 4644 5526 4662
rect 5508 4662 5526 4680
rect 5508 4680 5526 4698
rect 5508 4698 5526 4716
rect 5508 4716 5526 4734
rect 5508 4734 5526 4752
rect 5508 4752 5526 4770
rect 5508 4770 5526 4788
rect 5508 4788 5526 4806
rect 5508 4806 5526 4824
rect 5508 4824 5526 4842
rect 5508 4842 5526 4860
rect 5508 4860 5526 4878
rect 5508 4878 5526 4896
rect 5508 4896 5526 4914
rect 5508 5130 5526 5148
rect 5508 5148 5526 5166
rect 5508 5166 5526 5184
rect 5508 5184 5526 5202
rect 5508 5202 5526 5220
rect 5508 5220 5526 5238
rect 5508 5238 5526 5256
rect 5508 5256 5526 5274
rect 5508 5274 5526 5292
rect 5508 5292 5526 5310
rect 5508 5310 5526 5328
rect 5508 5328 5526 5346
rect 5508 5346 5526 5364
rect 5508 5364 5526 5382
rect 5508 5382 5526 5400
rect 5508 5400 5526 5418
rect 5508 5418 5526 5436
rect 5508 5436 5526 5454
rect 5508 5454 5526 5472
rect 5508 5472 5526 5490
rect 5508 5490 5526 5508
rect 5508 5508 5526 5526
rect 5508 5526 5526 5544
rect 5508 5544 5526 5562
rect 5508 5562 5526 5580
rect 5508 5580 5526 5598
rect 5508 5598 5526 5616
rect 5508 5616 5526 5634
rect 5508 5634 5526 5652
rect 5508 5652 5526 5670
rect 5508 5670 5526 5688
rect 5508 5688 5526 5706
rect 5508 5706 5526 5724
rect 5508 5724 5526 5742
rect 5508 5742 5526 5760
rect 5508 5760 5526 5778
rect 5508 5778 5526 5796
rect 5508 5796 5526 5814
rect 5508 5814 5526 5832
rect 5508 5832 5526 5850
rect 5508 5850 5526 5868
rect 5508 5868 5526 5886
rect 5508 5886 5526 5904
rect 5508 5904 5526 5922
rect 5508 5922 5526 5940
rect 5508 5940 5526 5958
rect 5508 5958 5526 5976
rect 5508 5976 5526 5994
rect 5508 5994 5526 6012
rect 5508 6012 5526 6030
rect 5508 6030 5526 6048
rect 5508 6048 5526 6066
rect 5508 6066 5526 6084
rect 5508 6084 5526 6102
rect 5508 6102 5526 6120
rect 5508 6120 5526 6138
rect 5508 6138 5526 6156
rect 5508 6156 5526 6174
rect 5508 6174 5526 6192
rect 5508 6192 5526 6210
rect 5508 6210 5526 6228
rect 5508 6228 5526 6246
rect 5508 6246 5526 6264
rect 5508 6264 5526 6282
rect 5508 6282 5526 6300
rect 5508 6300 5526 6318
rect 5508 6318 5526 6336
rect 5508 6336 5526 6354
rect 5508 6354 5526 6372
rect 5508 6372 5526 6390
rect 5508 6390 5526 6408
rect 5508 6408 5526 6426
rect 5508 6426 5526 6444
rect 5508 6444 5526 6462
rect 5508 6462 5526 6480
rect 5508 6480 5526 6498
rect 5508 6498 5526 6516
rect 5508 6516 5526 6534
rect 5508 6534 5526 6552
rect 5508 6552 5526 6570
rect 5508 6570 5526 6588
rect 5508 6588 5526 6606
rect 5508 6606 5526 6624
rect 5508 6624 5526 6642
rect 5508 6642 5526 6660
rect 5508 6660 5526 6678
rect 5508 6678 5526 6696
rect 5508 6696 5526 6714
rect 5508 6714 5526 6732
rect 5508 6732 5526 6750
rect 5508 6750 5526 6768
rect 5508 6768 5526 6786
rect 5508 6786 5526 6804
rect 5508 6804 5526 6822
rect 5508 6822 5526 6840
rect 5508 6840 5526 6858
rect 5508 6858 5526 6876
rect 5508 6876 5526 6894
rect 5508 6894 5526 6912
rect 5508 6912 5526 6930
rect 5508 6930 5526 6948
rect 5508 6948 5526 6966
rect 5508 6966 5526 6984
rect 5508 6984 5526 7002
rect 5508 7002 5526 7020
rect 5508 7020 5526 7038
rect 5508 7038 5526 7056
rect 5508 7056 5526 7074
rect 5508 7074 5526 7092
rect 5508 7092 5526 7110
rect 5508 7110 5526 7128
rect 5508 7128 5526 7146
rect 5508 7146 5526 7164
rect 5508 7164 5526 7182
rect 5508 7182 5526 7200
rect 5508 7200 5526 7218
rect 5508 7218 5526 7236
rect 5508 7236 5526 7254
rect 5508 7254 5526 7272
rect 5508 7272 5526 7290
rect 5508 7290 5526 7308
rect 5508 7308 5526 7326
rect 5508 7326 5526 7344
rect 5508 7344 5526 7362
rect 5508 7362 5526 7380
rect 5508 7380 5526 7398
rect 5508 7398 5526 7416
rect 5508 7416 5526 7434
rect 5508 7434 5526 7452
rect 5508 7452 5526 7470
rect 5508 7470 5526 7488
rect 5508 7488 5526 7506
rect 5508 7506 5526 7524
rect 5508 7524 5526 7542
rect 5508 7542 5526 7560
rect 5508 7560 5526 7578
rect 5508 7578 5526 7596
rect 5508 7596 5526 7614
rect 5508 7614 5526 7632
rect 5508 7632 5526 7650
rect 5508 7650 5526 7668
rect 5508 7668 5526 7686
rect 5508 7686 5526 7704
rect 5508 7704 5526 7722
rect 5508 7722 5526 7740
rect 5508 7740 5526 7758
rect 5508 7758 5526 7776
rect 5508 7776 5526 7794
rect 5508 7794 5526 7812
rect 5508 7812 5526 7830
rect 5508 7830 5526 7848
rect 5508 7848 5526 7866
rect 5508 7866 5526 7884
rect 5508 7884 5526 7902
rect 5508 7902 5526 7920
rect 5508 7920 5526 7938
rect 5508 7938 5526 7956
rect 5508 7956 5526 7974
rect 5508 7974 5526 7992
rect 5508 7992 5526 8010
rect 5508 8010 5526 8028
rect 5508 8028 5526 8046
rect 5508 8046 5526 8064
rect 5508 8064 5526 8082
rect 5508 8082 5526 8100
rect 5508 8100 5526 8118
rect 5508 8118 5526 8136
rect 5508 8136 5526 8154
rect 5508 8154 5526 8172
rect 5508 8172 5526 8190
rect 5508 8190 5526 8208
rect 5508 8208 5526 8226
rect 5508 8226 5526 8244
rect 5508 8244 5526 8262
rect 5508 8262 5526 8280
rect 5508 8280 5526 8298
rect 5508 8298 5526 8316
rect 5508 8316 5526 8334
rect 5508 8334 5526 8352
rect 5508 8352 5526 8370
rect 5508 8370 5526 8388
rect 5508 8388 5526 8406
rect 5508 8406 5526 8424
rect 5508 8424 5526 8442
rect 5508 8442 5526 8460
rect 5508 8460 5526 8478
rect 5508 8478 5526 8496
rect 5508 8496 5526 8514
rect 5508 8514 5526 8532
rect 5508 8532 5526 8550
rect 5508 8550 5526 8568
rect 5526 540 5544 558
rect 5526 558 5544 576
rect 5526 576 5544 594
rect 5526 594 5544 612
rect 5526 612 5544 630
rect 5526 630 5544 648
rect 5526 648 5544 666
rect 5526 666 5544 684
rect 5526 684 5544 702
rect 5526 702 5544 720
rect 5526 720 5544 738
rect 5526 738 5544 756
rect 5526 756 5544 774
rect 5526 774 5544 792
rect 5526 792 5544 810
rect 5526 810 5544 828
rect 5526 828 5544 846
rect 5526 846 5544 864
rect 5526 864 5544 882
rect 5526 882 5544 900
rect 5526 900 5544 918
rect 5526 918 5544 936
rect 5526 1062 5544 1080
rect 5526 1080 5544 1098
rect 5526 1098 5544 1116
rect 5526 1116 5544 1134
rect 5526 1134 5544 1152
rect 5526 1152 5544 1170
rect 5526 1170 5544 1188
rect 5526 1188 5544 1206
rect 5526 1206 5544 1224
rect 5526 1224 5544 1242
rect 5526 1242 5544 1260
rect 5526 1260 5544 1278
rect 5526 1278 5544 1296
rect 5526 1296 5544 1314
rect 5526 1314 5544 1332
rect 5526 1332 5544 1350
rect 5526 1350 5544 1368
rect 5526 1368 5544 1386
rect 5526 1386 5544 1404
rect 5526 1404 5544 1422
rect 5526 1422 5544 1440
rect 5526 1440 5544 1458
rect 5526 1458 5544 1476
rect 5526 1476 5544 1494
rect 5526 1494 5544 1512
rect 5526 1512 5544 1530
rect 5526 1530 5544 1548
rect 5526 1548 5544 1566
rect 5526 1566 5544 1584
rect 5526 1584 5544 1602
rect 5526 1602 5544 1620
rect 5526 1620 5544 1638
rect 5526 1638 5544 1656
rect 5526 1656 5544 1674
rect 5526 1674 5544 1692
rect 5526 1692 5544 1710
rect 5526 1710 5544 1728
rect 5526 1728 5544 1746
rect 5526 1746 5544 1764
rect 5526 1764 5544 1782
rect 5526 1782 5544 1800
rect 5526 1800 5544 1818
rect 5526 1818 5544 1836
rect 5526 1836 5544 1854
rect 5526 1854 5544 1872
rect 5526 1872 5544 1890
rect 5526 1890 5544 1908
rect 5526 1908 5544 1926
rect 5526 1926 5544 1944
rect 5526 1944 5544 1962
rect 5526 1962 5544 1980
rect 5526 1980 5544 1998
rect 5526 1998 5544 2016
rect 5526 2016 5544 2034
rect 5526 2034 5544 2052
rect 5526 2052 5544 2070
rect 5526 2070 5544 2088
rect 5526 2088 5544 2106
rect 5526 2106 5544 2124
rect 5526 2124 5544 2142
rect 5526 2142 5544 2160
rect 5526 2160 5544 2178
rect 5526 2178 5544 2196
rect 5526 2196 5544 2214
rect 5526 2214 5544 2232
rect 5526 2232 5544 2250
rect 5526 2250 5544 2268
rect 5526 2268 5544 2286
rect 5526 2286 5544 2304
rect 5526 2304 5544 2322
rect 5526 2322 5544 2340
rect 5526 2340 5544 2358
rect 5526 2358 5544 2376
rect 5526 2376 5544 2394
rect 5526 2394 5544 2412
rect 5526 2412 5544 2430
rect 5526 2430 5544 2448
rect 5526 2448 5544 2466
rect 5526 2466 5544 2484
rect 5526 2484 5544 2502
rect 5526 2502 5544 2520
rect 5526 2520 5544 2538
rect 5526 2736 5544 2754
rect 5526 2754 5544 2772
rect 5526 2772 5544 2790
rect 5526 2790 5544 2808
rect 5526 2808 5544 2826
rect 5526 2826 5544 2844
rect 5526 2844 5544 2862
rect 5526 2862 5544 2880
rect 5526 2880 5544 2898
rect 5526 2898 5544 2916
rect 5526 2916 5544 2934
rect 5526 2934 5544 2952
rect 5526 2952 5544 2970
rect 5526 2970 5544 2988
rect 5526 2988 5544 3006
rect 5526 3006 5544 3024
rect 5526 3024 5544 3042
rect 5526 3042 5544 3060
rect 5526 3060 5544 3078
rect 5526 3078 5544 3096
rect 5526 3096 5544 3114
rect 5526 3114 5544 3132
rect 5526 3132 5544 3150
rect 5526 3150 5544 3168
rect 5526 3168 5544 3186
rect 5526 3186 5544 3204
rect 5526 3204 5544 3222
rect 5526 3222 5544 3240
rect 5526 3240 5544 3258
rect 5526 3258 5544 3276
rect 5526 3276 5544 3294
rect 5526 3294 5544 3312
rect 5526 3312 5544 3330
rect 5526 3330 5544 3348
rect 5526 3348 5544 3366
rect 5526 3366 5544 3384
rect 5526 3384 5544 3402
rect 5526 3402 5544 3420
rect 5526 3420 5544 3438
rect 5526 3438 5544 3456
rect 5526 3456 5544 3474
rect 5526 3474 5544 3492
rect 5526 3492 5544 3510
rect 5526 3510 5544 3528
rect 5526 3528 5544 3546
rect 5526 3546 5544 3564
rect 5526 3564 5544 3582
rect 5526 3582 5544 3600
rect 5526 3600 5544 3618
rect 5526 3618 5544 3636
rect 5526 3636 5544 3654
rect 5526 3654 5544 3672
rect 5526 3672 5544 3690
rect 5526 3690 5544 3708
rect 5526 3708 5544 3726
rect 5526 3726 5544 3744
rect 5526 3744 5544 3762
rect 5526 3762 5544 3780
rect 5526 3780 5544 3798
rect 5526 3798 5544 3816
rect 5526 3816 5544 3834
rect 5526 3834 5544 3852
rect 5526 3852 5544 3870
rect 5526 3870 5544 3888
rect 5526 3888 5544 3906
rect 5526 3906 5544 3924
rect 5526 3924 5544 3942
rect 5526 3942 5544 3960
rect 5526 3960 5544 3978
rect 5526 3978 5544 3996
rect 5526 3996 5544 4014
rect 5526 4014 5544 4032
rect 5526 4032 5544 4050
rect 5526 4050 5544 4068
rect 5526 4068 5544 4086
rect 5526 4086 5544 4104
rect 5526 4104 5544 4122
rect 5526 4122 5544 4140
rect 5526 4140 5544 4158
rect 5526 4158 5544 4176
rect 5526 4176 5544 4194
rect 5526 4194 5544 4212
rect 5526 4212 5544 4230
rect 5526 4230 5544 4248
rect 5526 4248 5544 4266
rect 5526 4266 5544 4284
rect 5526 4284 5544 4302
rect 5526 4302 5544 4320
rect 5526 4320 5544 4338
rect 5526 4338 5544 4356
rect 5526 4356 5544 4374
rect 5526 4374 5544 4392
rect 5526 4392 5544 4410
rect 5526 4410 5544 4428
rect 5526 4428 5544 4446
rect 5526 4446 5544 4464
rect 5526 4464 5544 4482
rect 5526 4482 5544 4500
rect 5526 4500 5544 4518
rect 5526 4518 5544 4536
rect 5526 4536 5544 4554
rect 5526 4554 5544 4572
rect 5526 4572 5544 4590
rect 5526 4590 5544 4608
rect 5526 4608 5544 4626
rect 5526 4626 5544 4644
rect 5526 4644 5544 4662
rect 5526 4662 5544 4680
rect 5526 4680 5544 4698
rect 5526 4698 5544 4716
rect 5526 4716 5544 4734
rect 5526 4734 5544 4752
rect 5526 4752 5544 4770
rect 5526 4770 5544 4788
rect 5526 4788 5544 4806
rect 5526 4806 5544 4824
rect 5526 4824 5544 4842
rect 5526 4842 5544 4860
rect 5526 4860 5544 4878
rect 5526 4878 5544 4896
rect 5526 4896 5544 4914
rect 5526 4914 5544 4932
rect 5526 5148 5544 5166
rect 5526 5166 5544 5184
rect 5526 5184 5544 5202
rect 5526 5202 5544 5220
rect 5526 5220 5544 5238
rect 5526 5238 5544 5256
rect 5526 5256 5544 5274
rect 5526 5274 5544 5292
rect 5526 5292 5544 5310
rect 5526 5310 5544 5328
rect 5526 5328 5544 5346
rect 5526 5346 5544 5364
rect 5526 5364 5544 5382
rect 5526 5382 5544 5400
rect 5526 5400 5544 5418
rect 5526 5418 5544 5436
rect 5526 5436 5544 5454
rect 5526 5454 5544 5472
rect 5526 5472 5544 5490
rect 5526 5490 5544 5508
rect 5526 5508 5544 5526
rect 5526 5526 5544 5544
rect 5526 5544 5544 5562
rect 5526 5562 5544 5580
rect 5526 5580 5544 5598
rect 5526 5598 5544 5616
rect 5526 5616 5544 5634
rect 5526 5634 5544 5652
rect 5526 5652 5544 5670
rect 5526 5670 5544 5688
rect 5526 5688 5544 5706
rect 5526 5706 5544 5724
rect 5526 5724 5544 5742
rect 5526 5742 5544 5760
rect 5526 5760 5544 5778
rect 5526 5778 5544 5796
rect 5526 5796 5544 5814
rect 5526 5814 5544 5832
rect 5526 5832 5544 5850
rect 5526 5850 5544 5868
rect 5526 5868 5544 5886
rect 5526 5886 5544 5904
rect 5526 5904 5544 5922
rect 5526 5922 5544 5940
rect 5526 5940 5544 5958
rect 5526 5958 5544 5976
rect 5526 5976 5544 5994
rect 5526 5994 5544 6012
rect 5526 6012 5544 6030
rect 5526 6030 5544 6048
rect 5526 6048 5544 6066
rect 5526 6066 5544 6084
rect 5526 6084 5544 6102
rect 5526 6102 5544 6120
rect 5526 6120 5544 6138
rect 5526 6138 5544 6156
rect 5526 6156 5544 6174
rect 5526 6174 5544 6192
rect 5526 6192 5544 6210
rect 5526 6210 5544 6228
rect 5526 6228 5544 6246
rect 5526 6246 5544 6264
rect 5526 6264 5544 6282
rect 5526 6282 5544 6300
rect 5526 6300 5544 6318
rect 5526 6318 5544 6336
rect 5526 6336 5544 6354
rect 5526 6354 5544 6372
rect 5526 6372 5544 6390
rect 5526 6390 5544 6408
rect 5526 6408 5544 6426
rect 5526 6426 5544 6444
rect 5526 6444 5544 6462
rect 5526 6462 5544 6480
rect 5526 6480 5544 6498
rect 5526 6498 5544 6516
rect 5526 6516 5544 6534
rect 5526 6534 5544 6552
rect 5526 6552 5544 6570
rect 5526 6570 5544 6588
rect 5526 6588 5544 6606
rect 5526 6606 5544 6624
rect 5526 6624 5544 6642
rect 5526 6642 5544 6660
rect 5526 6660 5544 6678
rect 5526 6678 5544 6696
rect 5526 6696 5544 6714
rect 5526 6714 5544 6732
rect 5526 6732 5544 6750
rect 5526 6750 5544 6768
rect 5526 6768 5544 6786
rect 5526 6786 5544 6804
rect 5526 6804 5544 6822
rect 5526 6822 5544 6840
rect 5526 6840 5544 6858
rect 5526 6858 5544 6876
rect 5526 6876 5544 6894
rect 5526 6894 5544 6912
rect 5526 6912 5544 6930
rect 5526 6930 5544 6948
rect 5526 6948 5544 6966
rect 5526 6966 5544 6984
rect 5526 6984 5544 7002
rect 5526 7002 5544 7020
rect 5526 7020 5544 7038
rect 5526 7038 5544 7056
rect 5526 7056 5544 7074
rect 5526 7074 5544 7092
rect 5526 7092 5544 7110
rect 5526 7110 5544 7128
rect 5526 7128 5544 7146
rect 5526 7146 5544 7164
rect 5526 7164 5544 7182
rect 5526 7182 5544 7200
rect 5526 7200 5544 7218
rect 5526 7218 5544 7236
rect 5526 7236 5544 7254
rect 5526 7254 5544 7272
rect 5526 7272 5544 7290
rect 5526 7290 5544 7308
rect 5526 7308 5544 7326
rect 5526 7326 5544 7344
rect 5526 7344 5544 7362
rect 5526 7362 5544 7380
rect 5526 7380 5544 7398
rect 5526 7398 5544 7416
rect 5526 7416 5544 7434
rect 5526 7434 5544 7452
rect 5526 7452 5544 7470
rect 5526 7470 5544 7488
rect 5526 7488 5544 7506
rect 5526 7506 5544 7524
rect 5526 7524 5544 7542
rect 5526 7542 5544 7560
rect 5526 7560 5544 7578
rect 5526 7578 5544 7596
rect 5526 7596 5544 7614
rect 5526 7614 5544 7632
rect 5526 7632 5544 7650
rect 5526 7650 5544 7668
rect 5526 7668 5544 7686
rect 5526 7686 5544 7704
rect 5526 7704 5544 7722
rect 5526 7722 5544 7740
rect 5526 7740 5544 7758
rect 5526 7758 5544 7776
rect 5526 7776 5544 7794
rect 5526 7794 5544 7812
rect 5526 7812 5544 7830
rect 5526 7830 5544 7848
rect 5526 7848 5544 7866
rect 5526 7866 5544 7884
rect 5526 7884 5544 7902
rect 5526 7902 5544 7920
rect 5526 7920 5544 7938
rect 5526 7938 5544 7956
rect 5526 7956 5544 7974
rect 5526 7974 5544 7992
rect 5526 7992 5544 8010
rect 5526 8010 5544 8028
rect 5526 8028 5544 8046
rect 5526 8046 5544 8064
rect 5526 8064 5544 8082
rect 5526 8082 5544 8100
rect 5526 8100 5544 8118
rect 5526 8118 5544 8136
rect 5526 8136 5544 8154
rect 5526 8154 5544 8172
rect 5526 8172 5544 8190
rect 5526 8190 5544 8208
rect 5526 8208 5544 8226
rect 5526 8226 5544 8244
rect 5526 8244 5544 8262
rect 5526 8262 5544 8280
rect 5526 8280 5544 8298
rect 5526 8298 5544 8316
rect 5526 8316 5544 8334
rect 5526 8334 5544 8352
rect 5526 8352 5544 8370
rect 5526 8370 5544 8388
rect 5526 8388 5544 8406
rect 5526 8406 5544 8424
rect 5526 8424 5544 8442
rect 5526 8442 5544 8460
rect 5526 8460 5544 8478
rect 5526 8478 5544 8496
rect 5526 8496 5544 8514
rect 5526 8514 5544 8532
rect 5526 8532 5544 8550
rect 5526 8550 5544 8568
rect 5526 8568 5544 8586
rect 5526 8586 5544 8604
rect 5544 558 5562 576
rect 5544 576 5562 594
rect 5544 594 5562 612
rect 5544 612 5562 630
rect 5544 630 5562 648
rect 5544 648 5562 666
rect 5544 666 5562 684
rect 5544 684 5562 702
rect 5544 702 5562 720
rect 5544 720 5562 738
rect 5544 738 5562 756
rect 5544 756 5562 774
rect 5544 774 5562 792
rect 5544 792 5562 810
rect 5544 810 5562 828
rect 5544 828 5562 846
rect 5544 846 5562 864
rect 5544 864 5562 882
rect 5544 882 5562 900
rect 5544 900 5562 918
rect 5544 918 5562 936
rect 5544 1080 5562 1098
rect 5544 1098 5562 1116
rect 5544 1116 5562 1134
rect 5544 1134 5562 1152
rect 5544 1152 5562 1170
rect 5544 1170 5562 1188
rect 5544 1188 5562 1206
rect 5544 1206 5562 1224
rect 5544 1224 5562 1242
rect 5544 1242 5562 1260
rect 5544 1260 5562 1278
rect 5544 1278 5562 1296
rect 5544 1296 5562 1314
rect 5544 1314 5562 1332
rect 5544 1332 5562 1350
rect 5544 1350 5562 1368
rect 5544 1368 5562 1386
rect 5544 1386 5562 1404
rect 5544 1404 5562 1422
rect 5544 1422 5562 1440
rect 5544 1440 5562 1458
rect 5544 1458 5562 1476
rect 5544 1476 5562 1494
rect 5544 1494 5562 1512
rect 5544 1512 5562 1530
rect 5544 1530 5562 1548
rect 5544 1548 5562 1566
rect 5544 1566 5562 1584
rect 5544 1584 5562 1602
rect 5544 1602 5562 1620
rect 5544 1620 5562 1638
rect 5544 1638 5562 1656
rect 5544 1656 5562 1674
rect 5544 1674 5562 1692
rect 5544 1692 5562 1710
rect 5544 1710 5562 1728
rect 5544 1728 5562 1746
rect 5544 1746 5562 1764
rect 5544 1764 5562 1782
rect 5544 1782 5562 1800
rect 5544 1800 5562 1818
rect 5544 1818 5562 1836
rect 5544 1836 5562 1854
rect 5544 1854 5562 1872
rect 5544 1872 5562 1890
rect 5544 1890 5562 1908
rect 5544 1908 5562 1926
rect 5544 1926 5562 1944
rect 5544 1944 5562 1962
rect 5544 1962 5562 1980
rect 5544 1980 5562 1998
rect 5544 1998 5562 2016
rect 5544 2016 5562 2034
rect 5544 2034 5562 2052
rect 5544 2052 5562 2070
rect 5544 2070 5562 2088
rect 5544 2088 5562 2106
rect 5544 2106 5562 2124
rect 5544 2124 5562 2142
rect 5544 2142 5562 2160
rect 5544 2160 5562 2178
rect 5544 2178 5562 2196
rect 5544 2196 5562 2214
rect 5544 2214 5562 2232
rect 5544 2232 5562 2250
rect 5544 2250 5562 2268
rect 5544 2268 5562 2286
rect 5544 2286 5562 2304
rect 5544 2304 5562 2322
rect 5544 2322 5562 2340
rect 5544 2340 5562 2358
rect 5544 2358 5562 2376
rect 5544 2376 5562 2394
rect 5544 2394 5562 2412
rect 5544 2412 5562 2430
rect 5544 2430 5562 2448
rect 5544 2448 5562 2466
rect 5544 2466 5562 2484
rect 5544 2484 5562 2502
rect 5544 2502 5562 2520
rect 5544 2520 5562 2538
rect 5544 2754 5562 2772
rect 5544 2772 5562 2790
rect 5544 2790 5562 2808
rect 5544 2808 5562 2826
rect 5544 2826 5562 2844
rect 5544 2844 5562 2862
rect 5544 2862 5562 2880
rect 5544 2880 5562 2898
rect 5544 2898 5562 2916
rect 5544 2916 5562 2934
rect 5544 2934 5562 2952
rect 5544 2952 5562 2970
rect 5544 2970 5562 2988
rect 5544 2988 5562 3006
rect 5544 3006 5562 3024
rect 5544 3024 5562 3042
rect 5544 3042 5562 3060
rect 5544 3060 5562 3078
rect 5544 3078 5562 3096
rect 5544 3096 5562 3114
rect 5544 3114 5562 3132
rect 5544 3132 5562 3150
rect 5544 3150 5562 3168
rect 5544 3168 5562 3186
rect 5544 3186 5562 3204
rect 5544 3204 5562 3222
rect 5544 3222 5562 3240
rect 5544 3240 5562 3258
rect 5544 3258 5562 3276
rect 5544 3276 5562 3294
rect 5544 3294 5562 3312
rect 5544 3312 5562 3330
rect 5544 3330 5562 3348
rect 5544 3348 5562 3366
rect 5544 3366 5562 3384
rect 5544 3384 5562 3402
rect 5544 3402 5562 3420
rect 5544 3420 5562 3438
rect 5544 3438 5562 3456
rect 5544 3456 5562 3474
rect 5544 3474 5562 3492
rect 5544 3492 5562 3510
rect 5544 3510 5562 3528
rect 5544 3528 5562 3546
rect 5544 3546 5562 3564
rect 5544 3564 5562 3582
rect 5544 3582 5562 3600
rect 5544 3600 5562 3618
rect 5544 3618 5562 3636
rect 5544 3636 5562 3654
rect 5544 3654 5562 3672
rect 5544 3672 5562 3690
rect 5544 3690 5562 3708
rect 5544 3708 5562 3726
rect 5544 3726 5562 3744
rect 5544 3744 5562 3762
rect 5544 3762 5562 3780
rect 5544 3780 5562 3798
rect 5544 3798 5562 3816
rect 5544 3816 5562 3834
rect 5544 3834 5562 3852
rect 5544 3852 5562 3870
rect 5544 3870 5562 3888
rect 5544 3888 5562 3906
rect 5544 3906 5562 3924
rect 5544 3924 5562 3942
rect 5544 3942 5562 3960
rect 5544 3960 5562 3978
rect 5544 3978 5562 3996
rect 5544 3996 5562 4014
rect 5544 4014 5562 4032
rect 5544 4032 5562 4050
rect 5544 4050 5562 4068
rect 5544 4068 5562 4086
rect 5544 4086 5562 4104
rect 5544 4104 5562 4122
rect 5544 4122 5562 4140
rect 5544 4140 5562 4158
rect 5544 4158 5562 4176
rect 5544 4176 5562 4194
rect 5544 4194 5562 4212
rect 5544 4212 5562 4230
rect 5544 4230 5562 4248
rect 5544 4248 5562 4266
rect 5544 4266 5562 4284
rect 5544 4284 5562 4302
rect 5544 4302 5562 4320
rect 5544 4320 5562 4338
rect 5544 4338 5562 4356
rect 5544 4356 5562 4374
rect 5544 4374 5562 4392
rect 5544 4392 5562 4410
rect 5544 4410 5562 4428
rect 5544 4428 5562 4446
rect 5544 4446 5562 4464
rect 5544 4464 5562 4482
rect 5544 4482 5562 4500
rect 5544 4500 5562 4518
rect 5544 4518 5562 4536
rect 5544 4536 5562 4554
rect 5544 4554 5562 4572
rect 5544 4572 5562 4590
rect 5544 4590 5562 4608
rect 5544 4608 5562 4626
rect 5544 4626 5562 4644
rect 5544 4644 5562 4662
rect 5544 4662 5562 4680
rect 5544 4680 5562 4698
rect 5544 4698 5562 4716
rect 5544 4716 5562 4734
rect 5544 4734 5562 4752
rect 5544 4752 5562 4770
rect 5544 4770 5562 4788
rect 5544 4788 5562 4806
rect 5544 4806 5562 4824
rect 5544 4824 5562 4842
rect 5544 4842 5562 4860
rect 5544 4860 5562 4878
rect 5544 4878 5562 4896
rect 5544 4896 5562 4914
rect 5544 4914 5562 4932
rect 5544 4932 5562 4950
rect 5544 5166 5562 5184
rect 5544 5184 5562 5202
rect 5544 5202 5562 5220
rect 5544 5220 5562 5238
rect 5544 5238 5562 5256
rect 5544 5256 5562 5274
rect 5544 5274 5562 5292
rect 5544 5292 5562 5310
rect 5544 5310 5562 5328
rect 5544 5328 5562 5346
rect 5544 5346 5562 5364
rect 5544 5364 5562 5382
rect 5544 5382 5562 5400
rect 5544 5400 5562 5418
rect 5544 5418 5562 5436
rect 5544 5436 5562 5454
rect 5544 5454 5562 5472
rect 5544 5472 5562 5490
rect 5544 5490 5562 5508
rect 5544 5508 5562 5526
rect 5544 5526 5562 5544
rect 5544 5544 5562 5562
rect 5544 5562 5562 5580
rect 5544 5580 5562 5598
rect 5544 5598 5562 5616
rect 5544 5616 5562 5634
rect 5544 5634 5562 5652
rect 5544 5652 5562 5670
rect 5544 5670 5562 5688
rect 5544 5688 5562 5706
rect 5544 5706 5562 5724
rect 5544 5724 5562 5742
rect 5544 5742 5562 5760
rect 5544 5760 5562 5778
rect 5544 5778 5562 5796
rect 5544 5796 5562 5814
rect 5544 5814 5562 5832
rect 5544 5832 5562 5850
rect 5544 5850 5562 5868
rect 5544 5868 5562 5886
rect 5544 5886 5562 5904
rect 5544 5904 5562 5922
rect 5544 5922 5562 5940
rect 5544 5940 5562 5958
rect 5544 5958 5562 5976
rect 5544 5976 5562 5994
rect 5544 5994 5562 6012
rect 5544 6012 5562 6030
rect 5544 6030 5562 6048
rect 5544 6048 5562 6066
rect 5544 6066 5562 6084
rect 5544 6084 5562 6102
rect 5544 6102 5562 6120
rect 5544 6120 5562 6138
rect 5544 6138 5562 6156
rect 5544 6156 5562 6174
rect 5544 6174 5562 6192
rect 5544 6192 5562 6210
rect 5544 6210 5562 6228
rect 5544 6228 5562 6246
rect 5544 6246 5562 6264
rect 5544 6264 5562 6282
rect 5544 6282 5562 6300
rect 5544 6300 5562 6318
rect 5544 6318 5562 6336
rect 5544 6336 5562 6354
rect 5544 6354 5562 6372
rect 5544 6372 5562 6390
rect 5544 6390 5562 6408
rect 5544 6408 5562 6426
rect 5544 6426 5562 6444
rect 5544 6444 5562 6462
rect 5544 6462 5562 6480
rect 5544 6480 5562 6498
rect 5544 6498 5562 6516
rect 5544 6516 5562 6534
rect 5544 6534 5562 6552
rect 5544 6552 5562 6570
rect 5544 6570 5562 6588
rect 5544 6588 5562 6606
rect 5544 6606 5562 6624
rect 5544 6624 5562 6642
rect 5544 6642 5562 6660
rect 5544 6660 5562 6678
rect 5544 6678 5562 6696
rect 5544 6696 5562 6714
rect 5544 6714 5562 6732
rect 5544 6732 5562 6750
rect 5544 6750 5562 6768
rect 5544 6768 5562 6786
rect 5544 6786 5562 6804
rect 5544 6804 5562 6822
rect 5544 6822 5562 6840
rect 5544 6840 5562 6858
rect 5544 6858 5562 6876
rect 5544 6876 5562 6894
rect 5544 6894 5562 6912
rect 5544 6912 5562 6930
rect 5544 6930 5562 6948
rect 5544 6948 5562 6966
rect 5544 6966 5562 6984
rect 5544 6984 5562 7002
rect 5544 7002 5562 7020
rect 5544 7020 5562 7038
rect 5544 7038 5562 7056
rect 5544 7056 5562 7074
rect 5544 7074 5562 7092
rect 5544 7092 5562 7110
rect 5544 7110 5562 7128
rect 5544 7128 5562 7146
rect 5544 7146 5562 7164
rect 5544 7164 5562 7182
rect 5544 7182 5562 7200
rect 5544 7200 5562 7218
rect 5544 7218 5562 7236
rect 5544 7236 5562 7254
rect 5544 7254 5562 7272
rect 5544 7272 5562 7290
rect 5544 7290 5562 7308
rect 5544 7308 5562 7326
rect 5544 7326 5562 7344
rect 5544 7344 5562 7362
rect 5544 7362 5562 7380
rect 5544 7380 5562 7398
rect 5544 7398 5562 7416
rect 5544 7416 5562 7434
rect 5544 7434 5562 7452
rect 5544 7452 5562 7470
rect 5544 7470 5562 7488
rect 5544 7488 5562 7506
rect 5544 7506 5562 7524
rect 5544 7524 5562 7542
rect 5544 7542 5562 7560
rect 5544 7560 5562 7578
rect 5544 7578 5562 7596
rect 5544 7596 5562 7614
rect 5544 7614 5562 7632
rect 5544 7632 5562 7650
rect 5544 7650 5562 7668
rect 5544 7668 5562 7686
rect 5544 7686 5562 7704
rect 5544 7704 5562 7722
rect 5544 7722 5562 7740
rect 5544 7740 5562 7758
rect 5544 7758 5562 7776
rect 5544 7776 5562 7794
rect 5544 7794 5562 7812
rect 5544 7812 5562 7830
rect 5544 7830 5562 7848
rect 5544 7848 5562 7866
rect 5544 7866 5562 7884
rect 5544 7884 5562 7902
rect 5544 7902 5562 7920
rect 5544 7920 5562 7938
rect 5544 7938 5562 7956
rect 5544 7956 5562 7974
rect 5544 7974 5562 7992
rect 5544 7992 5562 8010
rect 5544 8010 5562 8028
rect 5544 8028 5562 8046
rect 5544 8046 5562 8064
rect 5544 8064 5562 8082
rect 5544 8082 5562 8100
rect 5544 8100 5562 8118
rect 5544 8118 5562 8136
rect 5544 8136 5562 8154
rect 5544 8154 5562 8172
rect 5544 8172 5562 8190
rect 5544 8190 5562 8208
rect 5544 8208 5562 8226
rect 5544 8226 5562 8244
rect 5544 8244 5562 8262
rect 5544 8262 5562 8280
rect 5544 8280 5562 8298
rect 5544 8298 5562 8316
rect 5544 8316 5562 8334
rect 5544 8334 5562 8352
rect 5544 8352 5562 8370
rect 5544 8370 5562 8388
rect 5544 8388 5562 8406
rect 5544 8406 5562 8424
rect 5544 8424 5562 8442
rect 5544 8442 5562 8460
rect 5544 8460 5562 8478
rect 5544 8478 5562 8496
rect 5544 8496 5562 8514
rect 5544 8514 5562 8532
rect 5544 8532 5562 8550
rect 5544 8550 5562 8568
rect 5544 8568 5562 8586
rect 5544 8586 5562 8604
rect 5544 8604 5562 8622
rect 5562 558 5580 576
rect 5562 576 5580 594
rect 5562 594 5580 612
rect 5562 612 5580 630
rect 5562 630 5580 648
rect 5562 648 5580 666
rect 5562 666 5580 684
rect 5562 684 5580 702
rect 5562 702 5580 720
rect 5562 720 5580 738
rect 5562 738 5580 756
rect 5562 756 5580 774
rect 5562 774 5580 792
rect 5562 792 5580 810
rect 5562 810 5580 828
rect 5562 828 5580 846
rect 5562 846 5580 864
rect 5562 864 5580 882
rect 5562 882 5580 900
rect 5562 900 5580 918
rect 5562 918 5580 936
rect 5562 1080 5580 1098
rect 5562 1098 5580 1116
rect 5562 1116 5580 1134
rect 5562 1134 5580 1152
rect 5562 1152 5580 1170
rect 5562 1170 5580 1188
rect 5562 1188 5580 1206
rect 5562 1206 5580 1224
rect 5562 1224 5580 1242
rect 5562 1242 5580 1260
rect 5562 1260 5580 1278
rect 5562 1278 5580 1296
rect 5562 1296 5580 1314
rect 5562 1314 5580 1332
rect 5562 1332 5580 1350
rect 5562 1350 5580 1368
rect 5562 1368 5580 1386
rect 5562 1386 5580 1404
rect 5562 1404 5580 1422
rect 5562 1422 5580 1440
rect 5562 1440 5580 1458
rect 5562 1458 5580 1476
rect 5562 1476 5580 1494
rect 5562 1494 5580 1512
rect 5562 1512 5580 1530
rect 5562 1530 5580 1548
rect 5562 1548 5580 1566
rect 5562 1566 5580 1584
rect 5562 1584 5580 1602
rect 5562 1602 5580 1620
rect 5562 1620 5580 1638
rect 5562 1638 5580 1656
rect 5562 1656 5580 1674
rect 5562 1674 5580 1692
rect 5562 1692 5580 1710
rect 5562 1710 5580 1728
rect 5562 1728 5580 1746
rect 5562 1746 5580 1764
rect 5562 1764 5580 1782
rect 5562 1782 5580 1800
rect 5562 1800 5580 1818
rect 5562 1818 5580 1836
rect 5562 1836 5580 1854
rect 5562 1854 5580 1872
rect 5562 1872 5580 1890
rect 5562 1890 5580 1908
rect 5562 1908 5580 1926
rect 5562 1926 5580 1944
rect 5562 1944 5580 1962
rect 5562 1962 5580 1980
rect 5562 1980 5580 1998
rect 5562 1998 5580 2016
rect 5562 2016 5580 2034
rect 5562 2034 5580 2052
rect 5562 2052 5580 2070
rect 5562 2070 5580 2088
rect 5562 2088 5580 2106
rect 5562 2106 5580 2124
rect 5562 2124 5580 2142
rect 5562 2142 5580 2160
rect 5562 2160 5580 2178
rect 5562 2178 5580 2196
rect 5562 2196 5580 2214
rect 5562 2214 5580 2232
rect 5562 2232 5580 2250
rect 5562 2250 5580 2268
rect 5562 2268 5580 2286
rect 5562 2286 5580 2304
rect 5562 2304 5580 2322
rect 5562 2322 5580 2340
rect 5562 2340 5580 2358
rect 5562 2358 5580 2376
rect 5562 2376 5580 2394
rect 5562 2394 5580 2412
rect 5562 2412 5580 2430
rect 5562 2430 5580 2448
rect 5562 2448 5580 2466
rect 5562 2466 5580 2484
rect 5562 2484 5580 2502
rect 5562 2502 5580 2520
rect 5562 2520 5580 2538
rect 5562 2538 5580 2556
rect 5562 2754 5580 2772
rect 5562 2772 5580 2790
rect 5562 2790 5580 2808
rect 5562 2808 5580 2826
rect 5562 2826 5580 2844
rect 5562 2844 5580 2862
rect 5562 2862 5580 2880
rect 5562 2880 5580 2898
rect 5562 2898 5580 2916
rect 5562 2916 5580 2934
rect 5562 2934 5580 2952
rect 5562 2952 5580 2970
rect 5562 2970 5580 2988
rect 5562 2988 5580 3006
rect 5562 3006 5580 3024
rect 5562 3024 5580 3042
rect 5562 3042 5580 3060
rect 5562 3060 5580 3078
rect 5562 3078 5580 3096
rect 5562 3096 5580 3114
rect 5562 3114 5580 3132
rect 5562 3132 5580 3150
rect 5562 3150 5580 3168
rect 5562 3168 5580 3186
rect 5562 3186 5580 3204
rect 5562 3204 5580 3222
rect 5562 3222 5580 3240
rect 5562 3240 5580 3258
rect 5562 3258 5580 3276
rect 5562 3276 5580 3294
rect 5562 3294 5580 3312
rect 5562 3312 5580 3330
rect 5562 3330 5580 3348
rect 5562 3348 5580 3366
rect 5562 3366 5580 3384
rect 5562 3384 5580 3402
rect 5562 3402 5580 3420
rect 5562 3420 5580 3438
rect 5562 3438 5580 3456
rect 5562 3456 5580 3474
rect 5562 3474 5580 3492
rect 5562 3492 5580 3510
rect 5562 3510 5580 3528
rect 5562 3528 5580 3546
rect 5562 3546 5580 3564
rect 5562 3564 5580 3582
rect 5562 3582 5580 3600
rect 5562 3600 5580 3618
rect 5562 3618 5580 3636
rect 5562 3636 5580 3654
rect 5562 3654 5580 3672
rect 5562 3672 5580 3690
rect 5562 3690 5580 3708
rect 5562 3708 5580 3726
rect 5562 3726 5580 3744
rect 5562 3744 5580 3762
rect 5562 3762 5580 3780
rect 5562 3780 5580 3798
rect 5562 3798 5580 3816
rect 5562 3816 5580 3834
rect 5562 3834 5580 3852
rect 5562 3852 5580 3870
rect 5562 3870 5580 3888
rect 5562 3888 5580 3906
rect 5562 3906 5580 3924
rect 5562 3924 5580 3942
rect 5562 3942 5580 3960
rect 5562 3960 5580 3978
rect 5562 3978 5580 3996
rect 5562 3996 5580 4014
rect 5562 4014 5580 4032
rect 5562 4032 5580 4050
rect 5562 4050 5580 4068
rect 5562 4068 5580 4086
rect 5562 4086 5580 4104
rect 5562 4104 5580 4122
rect 5562 4122 5580 4140
rect 5562 4140 5580 4158
rect 5562 4158 5580 4176
rect 5562 4176 5580 4194
rect 5562 4194 5580 4212
rect 5562 4212 5580 4230
rect 5562 4230 5580 4248
rect 5562 4248 5580 4266
rect 5562 4266 5580 4284
rect 5562 4284 5580 4302
rect 5562 4302 5580 4320
rect 5562 4320 5580 4338
rect 5562 4338 5580 4356
rect 5562 4356 5580 4374
rect 5562 4374 5580 4392
rect 5562 4392 5580 4410
rect 5562 4410 5580 4428
rect 5562 4428 5580 4446
rect 5562 4446 5580 4464
rect 5562 4464 5580 4482
rect 5562 4482 5580 4500
rect 5562 4500 5580 4518
rect 5562 4518 5580 4536
rect 5562 4536 5580 4554
rect 5562 4554 5580 4572
rect 5562 4572 5580 4590
rect 5562 4590 5580 4608
rect 5562 4608 5580 4626
rect 5562 4626 5580 4644
rect 5562 4644 5580 4662
rect 5562 4662 5580 4680
rect 5562 4680 5580 4698
rect 5562 4698 5580 4716
rect 5562 4716 5580 4734
rect 5562 4734 5580 4752
rect 5562 4752 5580 4770
rect 5562 4770 5580 4788
rect 5562 4788 5580 4806
rect 5562 4806 5580 4824
rect 5562 4824 5580 4842
rect 5562 4842 5580 4860
rect 5562 4860 5580 4878
rect 5562 4878 5580 4896
rect 5562 4896 5580 4914
rect 5562 4914 5580 4932
rect 5562 4932 5580 4950
rect 5562 4950 5580 4968
rect 5562 5184 5580 5202
rect 5562 5202 5580 5220
rect 5562 5220 5580 5238
rect 5562 5238 5580 5256
rect 5562 5256 5580 5274
rect 5562 5274 5580 5292
rect 5562 5292 5580 5310
rect 5562 5310 5580 5328
rect 5562 5328 5580 5346
rect 5562 5346 5580 5364
rect 5562 5364 5580 5382
rect 5562 5382 5580 5400
rect 5562 5400 5580 5418
rect 5562 5418 5580 5436
rect 5562 5436 5580 5454
rect 5562 5454 5580 5472
rect 5562 5472 5580 5490
rect 5562 5490 5580 5508
rect 5562 5508 5580 5526
rect 5562 5526 5580 5544
rect 5562 5544 5580 5562
rect 5562 5562 5580 5580
rect 5562 5580 5580 5598
rect 5562 5598 5580 5616
rect 5562 5616 5580 5634
rect 5562 5634 5580 5652
rect 5562 5652 5580 5670
rect 5562 5670 5580 5688
rect 5562 5688 5580 5706
rect 5562 5706 5580 5724
rect 5562 5724 5580 5742
rect 5562 5742 5580 5760
rect 5562 5760 5580 5778
rect 5562 5778 5580 5796
rect 5562 5796 5580 5814
rect 5562 5814 5580 5832
rect 5562 5832 5580 5850
rect 5562 5850 5580 5868
rect 5562 5868 5580 5886
rect 5562 5886 5580 5904
rect 5562 5904 5580 5922
rect 5562 5922 5580 5940
rect 5562 5940 5580 5958
rect 5562 5958 5580 5976
rect 5562 5976 5580 5994
rect 5562 5994 5580 6012
rect 5562 6012 5580 6030
rect 5562 6030 5580 6048
rect 5562 6048 5580 6066
rect 5562 6066 5580 6084
rect 5562 6084 5580 6102
rect 5562 6102 5580 6120
rect 5562 6120 5580 6138
rect 5562 6138 5580 6156
rect 5562 6156 5580 6174
rect 5562 6174 5580 6192
rect 5562 6192 5580 6210
rect 5562 6210 5580 6228
rect 5562 6228 5580 6246
rect 5562 6246 5580 6264
rect 5562 6264 5580 6282
rect 5562 6282 5580 6300
rect 5562 6300 5580 6318
rect 5562 6318 5580 6336
rect 5562 6336 5580 6354
rect 5562 6354 5580 6372
rect 5562 6372 5580 6390
rect 5562 6390 5580 6408
rect 5562 6408 5580 6426
rect 5562 6426 5580 6444
rect 5562 6444 5580 6462
rect 5562 6462 5580 6480
rect 5562 6480 5580 6498
rect 5562 6498 5580 6516
rect 5562 6516 5580 6534
rect 5562 6534 5580 6552
rect 5562 6552 5580 6570
rect 5562 6570 5580 6588
rect 5562 6588 5580 6606
rect 5562 6606 5580 6624
rect 5562 6624 5580 6642
rect 5562 6642 5580 6660
rect 5562 6660 5580 6678
rect 5562 6678 5580 6696
rect 5562 6696 5580 6714
rect 5562 6714 5580 6732
rect 5562 6732 5580 6750
rect 5562 6750 5580 6768
rect 5562 6768 5580 6786
rect 5562 6786 5580 6804
rect 5562 6804 5580 6822
rect 5562 6822 5580 6840
rect 5562 6840 5580 6858
rect 5562 6858 5580 6876
rect 5562 6876 5580 6894
rect 5562 6894 5580 6912
rect 5562 6912 5580 6930
rect 5562 6930 5580 6948
rect 5562 6948 5580 6966
rect 5562 6966 5580 6984
rect 5562 6984 5580 7002
rect 5562 7002 5580 7020
rect 5562 7020 5580 7038
rect 5562 7038 5580 7056
rect 5562 7056 5580 7074
rect 5562 7074 5580 7092
rect 5562 7092 5580 7110
rect 5562 7110 5580 7128
rect 5562 7128 5580 7146
rect 5562 7146 5580 7164
rect 5562 7164 5580 7182
rect 5562 7182 5580 7200
rect 5562 7200 5580 7218
rect 5562 7218 5580 7236
rect 5562 7236 5580 7254
rect 5562 7254 5580 7272
rect 5562 7272 5580 7290
rect 5562 7290 5580 7308
rect 5562 7308 5580 7326
rect 5562 7326 5580 7344
rect 5562 7344 5580 7362
rect 5562 7362 5580 7380
rect 5562 7380 5580 7398
rect 5562 7398 5580 7416
rect 5562 7416 5580 7434
rect 5562 7434 5580 7452
rect 5562 7452 5580 7470
rect 5562 7470 5580 7488
rect 5562 7488 5580 7506
rect 5562 7506 5580 7524
rect 5562 7524 5580 7542
rect 5562 7542 5580 7560
rect 5562 7560 5580 7578
rect 5562 7578 5580 7596
rect 5562 7596 5580 7614
rect 5562 7614 5580 7632
rect 5562 7632 5580 7650
rect 5562 7650 5580 7668
rect 5562 7668 5580 7686
rect 5562 7686 5580 7704
rect 5562 7704 5580 7722
rect 5562 7722 5580 7740
rect 5562 7740 5580 7758
rect 5562 7758 5580 7776
rect 5562 7776 5580 7794
rect 5562 7794 5580 7812
rect 5562 7812 5580 7830
rect 5562 7830 5580 7848
rect 5562 7848 5580 7866
rect 5562 7866 5580 7884
rect 5562 7884 5580 7902
rect 5562 7902 5580 7920
rect 5562 7920 5580 7938
rect 5562 7938 5580 7956
rect 5562 7956 5580 7974
rect 5562 7974 5580 7992
rect 5562 7992 5580 8010
rect 5562 8010 5580 8028
rect 5562 8028 5580 8046
rect 5562 8046 5580 8064
rect 5562 8064 5580 8082
rect 5562 8082 5580 8100
rect 5562 8100 5580 8118
rect 5562 8118 5580 8136
rect 5562 8136 5580 8154
rect 5562 8154 5580 8172
rect 5562 8172 5580 8190
rect 5562 8190 5580 8208
rect 5562 8208 5580 8226
rect 5562 8226 5580 8244
rect 5562 8244 5580 8262
rect 5562 8262 5580 8280
rect 5562 8280 5580 8298
rect 5562 8298 5580 8316
rect 5562 8316 5580 8334
rect 5562 8334 5580 8352
rect 5562 8352 5580 8370
rect 5562 8370 5580 8388
rect 5562 8388 5580 8406
rect 5562 8406 5580 8424
rect 5562 8424 5580 8442
rect 5562 8442 5580 8460
rect 5562 8460 5580 8478
rect 5562 8478 5580 8496
rect 5562 8496 5580 8514
rect 5562 8514 5580 8532
rect 5562 8532 5580 8550
rect 5562 8550 5580 8568
rect 5562 8568 5580 8586
rect 5562 8586 5580 8604
rect 5562 8604 5580 8622
rect 5562 8622 5580 8640
rect 5580 576 5598 594
rect 5580 594 5598 612
rect 5580 612 5598 630
rect 5580 630 5598 648
rect 5580 648 5598 666
rect 5580 666 5598 684
rect 5580 684 5598 702
rect 5580 702 5598 720
rect 5580 720 5598 738
rect 5580 738 5598 756
rect 5580 756 5598 774
rect 5580 774 5598 792
rect 5580 792 5598 810
rect 5580 810 5598 828
rect 5580 828 5598 846
rect 5580 846 5598 864
rect 5580 864 5598 882
rect 5580 882 5598 900
rect 5580 900 5598 918
rect 5580 918 5598 936
rect 5580 936 5598 954
rect 5580 1080 5598 1098
rect 5580 1098 5598 1116
rect 5580 1116 5598 1134
rect 5580 1134 5598 1152
rect 5580 1152 5598 1170
rect 5580 1170 5598 1188
rect 5580 1188 5598 1206
rect 5580 1206 5598 1224
rect 5580 1224 5598 1242
rect 5580 1242 5598 1260
rect 5580 1260 5598 1278
rect 5580 1278 5598 1296
rect 5580 1296 5598 1314
rect 5580 1314 5598 1332
rect 5580 1332 5598 1350
rect 5580 1350 5598 1368
rect 5580 1368 5598 1386
rect 5580 1386 5598 1404
rect 5580 1404 5598 1422
rect 5580 1422 5598 1440
rect 5580 1440 5598 1458
rect 5580 1458 5598 1476
rect 5580 1476 5598 1494
rect 5580 1494 5598 1512
rect 5580 1512 5598 1530
rect 5580 1530 5598 1548
rect 5580 1548 5598 1566
rect 5580 1566 5598 1584
rect 5580 1584 5598 1602
rect 5580 1602 5598 1620
rect 5580 1620 5598 1638
rect 5580 1638 5598 1656
rect 5580 1656 5598 1674
rect 5580 1674 5598 1692
rect 5580 1692 5598 1710
rect 5580 1710 5598 1728
rect 5580 1728 5598 1746
rect 5580 1746 5598 1764
rect 5580 1764 5598 1782
rect 5580 1782 5598 1800
rect 5580 1800 5598 1818
rect 5580 1818 5598 1836
rect 5580 1836 5598 1854
rect 5580 1854 5598 1872
rect 5580 1872 5598 1890
rect 5580 1890 5598 1908
rect 5580 1908 5598 1926
rect 5580 1926 5598 1944
rect 5580 1944 5598 1962
rect 5580 1962 5598 1980
rect 5580 1980 5598 1998
rect 5580 1998 5598 2016
rect 5580 2016 5598 2034
rect 5580 2034 5598 2052
rect 5580 2052 5598 2070
rect 5580 2070 5598 2088
rect 5580 2088 5598 2106
rect 5580 2106 5598 2124
rect 5580 2124 5598 2142
rect 5580 2142 5598 2160
rect 5580 2160 5598 2178
rect 5580 2178 5598 2196
rect 5580 2196 5598 2214
rect 5580 2214 5598 2232
rect 5580 2232 5598 2250
rect 5580 2250 5598 2268
rect 5580 2268 5598 2286
rect 5580 2286 5598 2304
rect 5580 2304 5598 2322
rect 5580 2322 5598 2340
rect 5580 2340 5598 2358
rect 5580 2358 5598 2376
rect 5580 2376 5598 2394
rect 5580 2394 5598 2412
rect 5580 2412 5598 2430
rect 5580 2430 5598 2448
rect 5580 2448 5598 2466
rect 5580 2466 5598 2484
rect 5580 2484 5598 2502
rect 5580 2502 5598 2520
rect 5580 2520 5598 2538
rect 5580 2538 5598 2556
rect 5580 2772 5598 2790
rect 5580 2790 5598 2808
rect 5580 2808 5598 2826
rect 5580 2826 5598 2844
rect 5580 2844 5598 2862
rect 5580 2862 5598 2880
rect 5580 2880 5598 2898
rect 5580 2898 5598 2916
rect 5580 2916 5598 2934
rect 5580 2934 5598 2952
rect 5580 2952 5598 2970
rect 5580 2970 5598 2988
rect 5580 2988 5598 3006
rect 5580 3006 5598 3024
rect 5580 3024 5598 3042
rect 5580 3042 5598 3060
rect 5580 3060 5598 3078
rect 5580 3078 5598 3096
rect 5580 3096 5598 3114
rect 5580 3114 5598 3132
rect 5580 3132 5598 3150
rect 5580 3150 5598 3168
rect 5580 3168 5598 3186
rect 5580 3186 5598 3204
rect 5580 3204 5598 3222
rect 5580 3222 5598 3240
rect 5580 3240 5598 3258
rect 5580 3258 5598 3276
rect 5580 3276 5598 3294
rect 5580 3294 5598 3312
rect 5580 3312 5598 3330
rect 5580 3330 5598 3348
rect 5580 3348 5598 3366
rect 5580 3366 5598 3384
rect 5580 3384 5598 3402
rect 5580 3402 5598 3420
rect 5580 3420 5598 3438
rect 5580 3438 5598 3456
rect 5580 3456 5598 3474
rect 5580 3474 5598 3492
rect 5580 3492 5598 3510
rect 5580 3510 5598 3528
rect 5580 3528 5598 3546
rect 5580 3546 5598 3564
rect 5580 3564 5598 3582
rect 5580 3582 5598 3600
rect 5580 3600 5598 3618
rect 5580 3618 5598 3636
rect 5580 3636 5598 3654
rect 5580 3654 5598 3672
rect 5580 3672 5598 3690
rect 5580 3690 5598 3708
rect 5580 3708 5598 3726
rect 5580 3726 5598 3744
rect 5580 3744 5598 3762
rect 5580 3762 5598 3780
rect 5580 3780 5598 3798
rect 5580 3798 5598 3816
rect 5580 3816 5598 3834
rect 5580 3834 5598 3852
rect 5580 3852 5598 3870
rect 5580 3870 5598 3888
rect 5580 3888 5598 3906
rect 5580 3906 5598 3924
rect 5580 3924 5598 3942
rect 5580 3942 5598 3960
rect 5580 3960 5598 3978
rect 5580 3978 5598 3996
rect 5580 3996 5598 4014
rect 5580 4014 5598 4032
rect 5580 4032 5598 4050
rect 5580 4050 5598 4068
rect 5580 4068 5598 4086
rect 5580 4086 5598 4104
rect 5580 4104 5598 4122
rect 5580 4122 5598 4140
rect 5580 4140 5598 4158
rect 5580 4158 5598 4176
rect 5580 4176 5598 4194
rect 5580 4194 5598 4212
rect 5580 4212 5598 4230
rect 5580 4230 5598 4248
rect 5580 4248 5598 4266
rect 5580 4266 5598 4284
rect 5580 4284 5598 4302
rect 5580 4302 5598 4320
rect 5580 4320 5598 4338
rect 5580 4338 5598 4356
rect 5580 4356 5598 4374
rect 5580 4374 5598 4392
rect 5580 4392 5598 4410
rect 5580 4410 5598 4428
rect 5580 4428 5598 4446
rect 5580 4446 5598 4464
rect 5580 4464 5598 4482
rect 5580 4482 5598 4500
rect 5580 4500 5598 4518
rect 5580 4518 5598 4536
rect 5580 4536 5598 4554
rect 5580 4554 5598 4572
rect 5580 4572 5598 4590
rect 5580 4590 5598 4608
rect 5580 4608 5598 4626
rect 5580 4626 5598 4644
rect 5580 4644 5598 4662
rect 5580 4662 5598 4680
rect 5580 4680 5598 4698
rect 5580 4698 5598 4716
rect 5580 4716 5598 4734
rect 5580 4734 5598 4752
rect 5580 4752 5598 4770
rect 5580 4770 5598 4788
rect 5580 4788 5598 4806
rect 5580 4806 5598 4824
rect 5580 4824 5598 4842
rect 5580 4842 5598 4860
rect 5580 4860 5598 4878
rect 5580 4878 5598 4896
rect 5580 4896 5598 4914
rect 5580 4914 5598 4932
rect 5580 4932 5598 4950
rect 5580 4950 5598 4968
rect 5580 4968 5598 4986
rect 5580 5202 5598 5220
rect 5580 5220 5598 5238
rect 5580 5238 5598 5256
rect 5580 5256 5598 5274
rect 5580 5274 5598 5292
rect 5580 5292 5598 5310
rect 5580 5310 5598 5328
rect 5580 5328 5598 5346
rect 5580 5346 5598 5364
rect 5580 5364 5598 5382
rect 5580 5382 5598 5400
rect 5580 5400 5598 5418
rect 5580 5418 5598 5436
rect 5580 5436 5598 5454
rect 5580 5454 5598 5472
rect 5580 5472 5598 5490
rect 5580 5490 5598 5508
rect 5580 5508 5598 5526
rect 5580 5526 5598 5544
rect 5580 5544 5598 5562
rect 5580 5562 5598 5580
rect 5580 5580 5598 5598
rect 5580 5598 5598 5616
rect 5580 5616 5598 5634
rect 5580 5634 5598 5652
rect 5580 5652 5598 5670
rect 5580 5670 5598 5688
rect 5580 5688 5598 5706
rect 5580 5706 5598 5724
rect 5580 5724 5598 5742
rect 5580 5742 5598 5760
rect 5580 5760 5598 5778
rect 5580 5778 5598 5796
rect 5580 5796 5598 5814
rect 5580 5814 5598 5832
rect 5580 5832 5598 5850
rect 5580 5850 5598 5868
rect 5580 5868 5598 5886
rect 5580 5886 5598 5904
rect 5580 5904 5598 5922
rect 5580 5922 5598 5940
rect 5580 5940 5598 5958
rect 5580 5958 5598 5976
rect 5580 5976 5598 5994
rect 5580 5994 5598 6012
rect 5580 6012 5598 6030
rect 5580 6030 5598 6048
rect 5580 6048 5598 6066
rect 5580 6066 5598 6084
rect 5580 6084 5598 6102
rect 5580 6102 5598 6120
rect 5580 6120 5598 6138
rect 5580 6138 5598 6156
rect 5580 6156 5598 6174
rect 5580 6174 5598 6192
rect 5580 6192 5598 6210
rect 5580 6210 5598 6228
rect 5580 6228 5598 6246
rect 5580 6246 5598 6264
rect 5580 6264 5598 6282
rect 5580 6282 5598 6300
rect 5580 6300 5598 6318
rect 5580 6318 5598 6336
rect 5580 6336 5598 6354
rect 5580 6354 5598 6372
rect 5580 6372 5598 6390
rect 5580 6390 5598 6408
rect 5580 6408 5598 6426
rect 5580 6426 5598 6444
rect 5580 6444 5598 6462
rect 5580 6462 5598 6480
rect 5580 6480 5598 6498
rect 5580 6498 5598 6516
rect 5580 6516 5598 6534
rect 5580 6534 5598 6552
rect 5580 6552 5598 6570
rect 5580 6570 5598 6588
rect 5580 6588 5598 6606
rect 5580 6606 5598 6624
rect 5580 6624 5598 6642
rect 5580 6642 5598 6660
rect 5580 6660 5598 6678
rect 5580 6678 5598 6696
rect 5580 6696 5598 6714
rect 5580 6714 5598 6732
rect 5580 6732 5598 6750
rect 5580 6750 5598 6768
rect 5580 6768 5598 6786
rect 5580 6786 5598 6804
rect 5580 6804 5598 6822
rect 5580 6822 5598 6840
rect 5580 6840 5598 6858
rect 5580 6858 5598 6876
rect 5580 6876 5598 6894
rect 5580 6894 5598 6912
rect 5580 6912 5598 6930
rect 5580 6930 5598 6948
rect 5580 6948 5598 6966
rect 5580 6966 5598 6984
rect 5580 6984 5598 7002
rect 5580 7002 5598 7020
rect 5580 7020 5598 7038
rect 5580 7038 5598 7056
rect 5580 7056 5598 7074
rect 5580 7074 5598 7092
rect 5580 7092 5598 7110
rect 5580 7110 5598 7128
rect 5580 7128 5598 7146
rect 5580 7146 5598 7164
rect 5580 7164 5598 7182
rect 5580 7182 5598 7200
rect 5580 7200 5598 7218
rect 5580 7218 5598 7236
rect 5580 7236 5598 7254
rect 5580 7254 5598 7272
rect 5580 7272 5598 7290
rect 5580 7290 5598 7308
rect 5580 7308 5598 7326
rect 5580 7326 5598 7344
rect 5580 7344 5598 7362
rect 5580 7362 5598 7380
rect 5580 7380 5598 7398
rect 5580 7398 5598 7416
rect 5580 7416 5598 7434
rect 5580 7434 5598 7452
rect 5580 7452 5598 7470
rect 5580 7470 5598 7488
rect 5580 7488 5598 7506
rect 5580 7506 5598 7524
rect 5580 7524 5598 7542
rect 5580 7542 5598 7560
rect 5580 7560 5598 7578
rect 5580 7578 5598 7596
rect 5580 7596 5598 7614
rect 5580 7614 5598 7632
rect 5580 7632 5598 7650
rect 5580 7650 5598 7668
rect 5580 7668 5598 7686
rect 5580 7686 5598 7704
rect 5580 7704 5598 7722
rect 5580 7722 5598 7740
rect 5580 7740 5598 7758
rect 5580 7758 5598 7776
rect 5580 7776 5598 7794
rect 5580 7794 5598 7812
rect 5580 7812 5598 7830
rect 5580 7830 5598 7848
rect 5580 7848 5598 7866
rect 5580 7866 5598 7884
rect 5580 7884 5598 7902
rect 5580 7902 5598 7920
rect 5580 7920 5598 7938
rect 5580 7938 5598 7956
rect 5580 7956 5598 7974
rect 5580 7974 5598 7992
rect 5580 7992 5598 8010
rect 5580 8010 5598 8028
rect 5580 8028 5598 8046
rect 5580 8046 5598 8064
rect 5580 8064 5598 8082
rect 5580 8082 5598 8100
rect 5580 8100 5598 8118
rect 5580 8118 5598 8136
rect 5580 8136 5598 8154
rect 5580 8154 5598 8172
rect 5580 8172 5598 8190
rect 5580 8190 5598 8208
rect 5580 8208 5598 8226
rect 5580 8226 5598 8244
rect 5580 8244 5598 8262
rect 5580 8262 5598 8280
rect 5580 8280 5598 8298
rect 5580 8298 5598 8316
rect 5580 8316 5598 8334
rect 5580 8334 5598 8352
rect 5580 8352 5598 8370
rect 5580 8370 5598 8388
rect 5580 8388 5598 8406
rect 5580 8406 5598 8424
rect 5580 8424 5598 8442
rect 5580 8442 5598 8460
rect 5580 8460 5598 8478
rect 5580 8478 5598 8496
rect 5580 8496 5598 8514
rect 5580 8514 5598 8532
rect 5580 8532 5598 8550
rect 5580 8550 5598 8568
rect 5580 8568 5598 8586
rect 5580 8586 5598 8604
rect 5580 8604 5598 8622
rect 5580 8622 5598 8640
rect 5580 8640 5598 8658
rect 5580 8658 5598 8676
rect 5598 594 5616 612
rect 5598 612 5616 630
rect 5598 630 5616 648
rect 5598 648 5616 666
rect 5598 666 5616 684
rect 5598 684 5616 702
rect 5598 702 5616 720
rect 5598 720 5616 738
rect 5598 738 5616 756
rect 5598 756 5616 774
rect 5598 774 5616 792
rect 5598 792 5616 810
rect 5598 810 5616 828
rect 5598 828 5616 846
rect 5598 846 5616 864
rect 5598 864 5616 882
rect 5598 882 5616 900
rect 5598 900 5616 918
rect 5598 918 5616 936
rect 5598 936 5616 954
rect 5598 1098 5616 1116
rect 5598 1116 5616 1134
rect 5598 1134 5616 1152
rect 5598 1152 5616 1170
rect 5598 1170 5616 1188
rect 5598 1188 5616 1206
rect 5598 1206 5616 1224
rect 5598 1224 5616 1242
rect 5598 1242 5616 1260
rect 5598 1260 5616 1278
rect 5598 1278 5616 1296
rect 5598 1296 5616 1314
rect 5598 1314 5616 1332
rect 5598 1332 5616 1350
rect 5598 1350 5616 1368
rect 5598 1368 5616 1386
rect 5598 1386 5616 1404
rect 5598 1404 5616 1422
rect 5598 1422 5616 1440
rect 5598 1440 5616 1458
rect 5598 1458 5616 1476
rect 5598 1476 5616 1494
rect 5598 1494 5616 1512
rect 5598 1512 5616 1530
rect 5598 1530 5616 1548
rect 5598 1548 5616 1566
rect 5598 1566 5616 1584
rect 5598 1584 5616 1602
rect 5598 1602 5616 1620
rect 5598 1620 5616 1638
rect 5598 1638 5616 1656
rect 5598 1656 5616 1674
rect 5598 1674 5616 1692
rect 5598 1692 5616 1710
rect 5598 1710 5616 1728
rect 5598 1728 5616 1746
rect 5598 1746 5616 1764
rect 5598 1764 5616 1782
rect 5598 1782 5616 1800
rect 5598 1800 5616 1818
rect 5598 1818 5616 1836
rect 5598 1836 5616 1854
rect 5598 1854 5616 1872
rect 5598 1872 5616 1890
rect 5598 1890 5616 1908
rect 5598 1908 5616 1926
rect 5598 1926 5616 1944
rect 5598 1944 5616 1962
rect 5598 1962 5616 1980
rect 5598 1980 5616 1998
rect 5598 1998 5616 2016
rect 5598 2016 5616 2034
rect 5598 2034 5616 2052
rect 5598 2052 5616 2070
rect 5598 2070 5616 2088
rect 5598 2088 5616 2106
rect 5598 2106 5616 2124
rect 5598 2124 5616 2142
rect 5598 2142 5616 2160
rect 5598 2160 5616 2178
rect 5598 2178 5616 2196
rect 5598 2196 5616 2214
rect 5598 2214 5616 2232
rect 5598 2232 5616 2250
rect 5598 2250 5616 2268
rect 5598 2268 5616 2286
rect 5598 2286 5616 2304
rect 5598 2304 5616 2322
rect 5598 2322 5616 2340
rect 5598 2340 5616 2358
rect 5598 2358 5616 2376
rect 5598 2376 5616 2394
rect 5598 2394 5616 2412
rect 5598 2412 5616 2430
rect 5598 2430 5616 2448
rect 5598 2448 5616 2466
rect 5598 2466 5616 2484
rect 5598 2484 5616 2502
rect 5598 2502 5616 2520
rect 5598 2520 5616 2538
rect 5598 2538 5616 2556
rect 5598 2556 5616 2574
rect 5598 2772 5616 2790
rect 5598 2790 5616 2808
rect 5598 2808 5616 2826
rect 5598 2826 5616 2844
rect 5598 2844 5616 2862
rect 5598 2862 5616 2880
rect 5598 2880 5616 2898
rect 5598 2898 5616 2916
rect 5598 2916 5616 2934
rect 5598 2934 5616 2952
rect 5598 2952 5616 2970
rect 5598 2970 5616 2988
rect 5598 2988 5616 3006
rect 5598 3006 5616 3024
rect 5598 3024 5616 3042
rect 5598 3042 5616 3060
rect 5598 3060 5616 3078
rect 5598 3078 5616 3096
rect 5598 3096 5616 3114
rect 5598 3114 5616 3132
rect 5598 3132 5616 3150
rect 5598 3150 5616 3168
rect 5598 3168 5616 3186
rect 5598 3186 5616 3204
rect 5598 3204 5616 3222
rect 5598 3222 5616 3240
rect 5598 3240 5616 3258
rect 5598 3258 5616 3276
rect 5598 3276 5616 3294
rect 5598 3294 5616 3312
rect 5598 3312 5616 3330
rect 5598 3330 5616 3348
rect 5598 3348 5616 3366
rect 5598 3366 5616 3384
rect 5598 3384 5616 3402
rect 5598 3402 5616 3420
rect 5598 3420 5616 3438
rect 5598 3438 5616 3456
rect 5598 3456 5616 3474
rect 5598 3474 5616 3492
rect 5598 3492 5616 3510
rect 5598 3510 5616 3528
rect 5598 3528 5616 3546
rect 5598 3546 5616 3564
rect 5598 3564 5616 3582
rect 5598 3582 5616 3600
rect 5598 3600 5616 3618
rect 5598 3618 5616 3636
rect 5598 3636 5616 3654
rect 5598 3654 5616 3672
rect 5598 3672 5616 3690
rect 5598 3690 5616 3708
rect 5598 3708 5616 3726
rect 5598 3726 5616 3744
rect 5598 3744 5616 3762
rect 5598 3762 5616 3780
rect 5598 3780 5616 3798
rect 5598 3798 5616 3816
rect 5598 3816 5616 3834
rect 5598 3834 5616 3852
rect 5598 3852 5616 3870
rect 5598 3870 5616 3888
rect 5598 3888 5616 3906
rect 5598 3906 5616 3924
rect 5598 3924 5616 3942
rect 5598 3942 5616 3960
rect 5598 3960 5616 3978
rect 5598 3978 5616 3996
rect 5598 3996 5616 4014
rect 5598 4014 5616 4032
rect 5598 4032 5616 4050
rect 5598 4050 5616 4068
rect 5598 4068 5616 4086
rect 5598 4086 5616 4104
rect 5598 4104 5616 4122
rect 5598 4122 5616 4140
rect 5598 4140 5616 4158
rect 5598 4158 5616 4176
rect 5598 4176 5616 4194
rect 5598 4194 5616 4212
rect 5598 4212 5616 4230
rect 5598 4230 5616 4248
rect 5598 4248 5616 4266
rect 5598 4266 5616 4284
rect 5598 4284 5616 4302
rect 5598 4302 5616 4320
rect 5598 4320 5616 4338
rect 5598 4338 5616 4356
rect 5598 4356 5616 4374
rect 5598 4374 5616 4392
rect 5598 4392 5616 4410
rect 5598 4410 5616 4428
rect 5598 4428 5616 4446
rect 5598 4446 5616 4464
rect 5598 4464 5616 4482
rect 5598 4482 5616 4500
rect 5598 4500 5616 4518
rect 5598 4518 5616 4536
rect 5598 4536 5616 4554
rect 5598 4554 5616 4572
rect 5598 4572 5616 4590
rect 5598 4590 5616 4608
rect 5598 4608 5616 4626
rect 5598 4626 5616 4644
rect 5598 4644 5616 4662
rect 5598 4662 5616 4680
rect 5598 4680 5616 4698
rect 5598 4698 5616 4716
rect 5598 4716 5616 4734
rect 5598 4734 5616 4752
rect 5598 4752 5616 4770
rect 5598 4770 5616 4788
rect 5598 4788 5616 4806
rect 5598 4806 5616 4824
rect 5598 4824 5616 4842
rect 5598 4842 5616 4860
rect 5598 4860 5616 4878
rect 5598 4878 5616 4896
rect 5598 4896 5616 4914
rect 5598 4914 5616 4932
rect 5598 4932 5616 4950
rect 5598 4950 5616 4968
rect 5598 4968 5616 4986
rect 5598 4986 5616 5004
rect 5598 5220 5616 5238
rect 5598 5238 5616 5256
rect 5598 5256 5616 5274
rect 5598 5274 5616 5292
rect 5598 5292 5616 5310
rect 5598 5310 5616 5328
rect 5598 5328 5616 5346
rect 5598 5346 5616 5364
rect 5598 5364 5616 5382
rect 5598 5382 5616 5400
rect 5598 5400 5616 5418
rect 5598 5418 5616 5436
rect 5598 5436 5616 5454
rect 5598 5454 5616 5472
rect 5598 5472 5616 5490
rect 5598 5490 5616 5508
rect 5598 5508 5616 5526
rect 5598 5526 5616 5544
rect 5598 5544 5616 5562
rect 5598 5562 5616 5580
rect 5598 5580 5616 5598
rect 5598 5598 5616 5616
rect 5598 5616 5616 5634
rect 5598 5634 5616 5652
rect 5598 5652 5616 5670
rect 5598 5670 5616 5688
rect 5598 5688 5616 5706
rect 5598 5706 5616 5724
rect 5598 5724 5616 5742
rect 5598 5742 5616 5760
rect 5598 5760 5616 5778
rect 5598 5778 5616 5796
rect 5598 5796 5616 5814
rect 5598 5814 5616 5832
rect 5598 5832 5616 5850
rect 5598 5850 5616 5868
rect 5598 5868 5616 5886
rect 5598 5886 5616 5904
rect 5598 5904 5616 5922
rect 5598 5922 5616 5940
rect 5598 5940 5616 5958
rect 5598 5958 5616 5976
rect 5598 5976 5616 5994
rect 5598 5994 5616 6012
rect 5598 6012 5616 6030
rect 5598 6030 5616 6048
rect 5598 6048 5616 6066
rect 5598 6066 5616 6084
rect 5598 6084 5616 6102
rect 5598 6102 5616 6120
rect 5598 6120 5616 6138
rect 5598 6138 5616 6156
rect 5598 6156 5616 6174
rect 5598 6174 5616 6192
rect 5598 6192 5616 6210
rect 5598 6210 5616 6228
rect 5598 6228 5616 6246
rect 5598 6246 5616 6264
rect 5598 6264 5616 6282
rect 5598 6282 5616 6300
rect 5598 6300 5616 6318
rect 5598 6318 5616 6336
rect 5598 6336 5616 6354
rect 5598 6354 5616 6372
rect 5598 6372 5616 6390
rect 5598 6390 5616 6408
rect 5598 6408 5616 6426
rect 5598 6426 5616 6444
rect 5598 6444 5616 6462
rect 5598 6462 5616 6480
rect 5598 6480 5616 6498
rect 5598 6498 5616 6516
rect 5598 6516 5616 6534
rect 5598 6534 5616 6552
rect 5598 6552 5616 6570
rect 5598 6570 5616 6588
rect 5598 6588 5616 6606
rect 5598 6606 5616 6624
rect 5598 6624 5616 6642
rect 5598 6642 5616 6660
rect 5598 6660 5616 6678
rect 5598 6678 5616 6696
rect 5598 6696 5616 6714
rect 5598 6714 5616 6732
rect 5598 6732 5616 6750
rect 5598 6750 5616 6768
rect 5598 6768 5616 6786
rect 5598 6786 5616 6804
rect 5598 6804 5616 6822
rect 5598 6822 5616 6840
rect 5598 6840 5616 6858
rect 5598 6858 5616 6876
rect 5598 6876 5616 6894
rect 5598 6894 5616 6912
rect 5598 6912 5616 6930
rect 5598 6930 5616 6948
rect 5598 6948 5616 6966
rect 5598 6966 5616 6984
rect 5598 6984 5616 7002
rect 5598 7002 5616 7020
rect 5598 7020 5616 7038
rect 5598 7038 5616 7056
rect 5598 7056 5616 7074
rect 5598 7074 5616 7092
rect 5598 7092 5616 7110
rect 5598 7110 5616 7128
rect 5598 7128 5616 7146
rect 5598 7146 5616 7164
rect 5598 7164 5616 7182
rect 5598 7182 5616 7200
rect 5598 7200 5616 7218
rect 5598 7218 5616 7236
rect 5598 7236 5616 7254
rect 5598 7254 5616 7272
rect 5598 7272 5616 7290
rect 5598 7290 5616 7308
rect 5598 7308 5616 7326
rect 5598 7326 5616 7344
rect 5598 7344 5616 7362
rect 5598 7362 5616 7380
rect 5598 7380 5616 7398
rect 5598 7398 5616 7416
rect 5598 7416 5616 7434
rect 5598 7434 5616 7452
rect 5598 7452 5616 7470
rect 5598 7470 5616 7488
rect 5598 7488 5616 7506
rect 5598 7506 5616 7524
rect 5598 7524 5616 7542
rect 5598 7542 5616 7560
rect 5598 7560 5616 7578
rect 5598 7578 5616 7596
rect 5598 7596 5616 7614
rect 5598 7614 5616 7632
rect 5598 7632 5616 7650
rect 5598 7650 5616 7668
rect 5598 7668 5616 7686
rect 5598 7686 5616 7704
rect 5598 7704 5616 7722
rect 5598 7722 5616 7740
rect 5598 7740 5616 7758
rect 5598 7758 5616 7776
rect 5598 7776 5616 7794
rect 5598 7794 5616 7812
rect 5598 7812 5616 7830
rect 5598 7830 5616 7848
rect 5598 7848 5616 7866
rect 5598 7866 5616 7884
rect 5598 7884 5616 7902
rect 5598 7902 5616 7920
rect 5598 7920 5616 7938
rect 5598 7938 5616 7956
rect 5598 7956 5616 7974
rect 5598 7974 5616 7992
rect 5598 7992 5616 8010
rect 5598 8010 5616 8028
rect 5598 8028 5616 8046
rect 5598 8046 5616 8064
rect 5598 8064 5616 8082
rect 5598 8082 5616 8100
rect 5598 8100 5616 8118
rect 5598 8118 5616 8136
rect 5598 8136 5616 8154
rect 5598 8154 5616 8172
rect 5598 8172 5616 8190
rect 5598 8190 5616 8208
rect 5598 8208 5616 8226
rect 5598 8226 5616 8244
rect 5598 8244 5616 8262
rect 5598 8262 5616 8280
rect 5598 8280 5616 8298
rect 5598 8298 5616 8316
rect 5598 8316 5616 8334
rect 5598 8334 5616 8352
rect 5598 8352 5616 8370
rect 5598 8370 5616 8388
rect 5598 8388 5616 8406
rect 5598 8406 5616 8424
rect 5598 8424 5616 8442
rect 5598 8442 5616 8460
rect 5598 8460 5616 8478
rect 5598 8478 5616 8496
rect 5598 8496 5616 8514
rect 5598 8514 5616 8532
rect 5598 8532 5616 8550
rect 5598 8550 5616 8568
rect 5598 8568 5616 8586
rect 5598 8586 5616 8604
rect 5598 8604 5616 8622
rect 5598 8622 5616 8640
rect 5598 8640 5616 8658
rect 5598 8658 5616 8676
rect 5598 8676 5616 8694
rect 5616 594 5634 612
rect 5616 612 5634 630
rect 5616 630 5634 648
rect 5616 648 5634 666
rect 5616 666 5634 684
rect 5616 684 5634 702
rect 5616 702 5634 720
rect 5616 720 5634 738
rect 5616 738 5634 756
rect 5616 756 5634 774
rect 5616 774 5634 792
rect 5616 792 5634 810
rect 5616 810 5634 828
rect 5616 828 5634 846
rect 5616 846 5634 864
rect 5616 864 5634 882
rect 5616 882 5634 900
rect 5616 900 5634 918
rect 5616 918 5634 936
rect 5616 936 5634 954
rect 5616 954 5634 972
rect 5616 1098 5634 1116
rect 5616 1116 5634 1134
rect 5616 1134 5634 1152
rect 5616 1152 5634 1170
rect 5616 1170 5634 1188
rect 5616 1188 5634 1206
rect 5616 1206 5634 1224
rect 5616 1224 5634 1242
rect 5616 1242 5634 1260
rect 5616 1260 5634 1278
rect 5616 1278 5634 1296
rect 5616 1296 5634 1314
rect 5616 1314 5634 1332
rect 5616 1332 5634 1350
rect 5616 1350 5634 1368
rect 5616 1368 5634 1386
rect 5616 1386 5634 1404
rect 5616 1404 5634 1422
rect 5616 1422 5634 1440
rect 5616 1440 5634 1458
rect 5616 1458 5634 1476
rect 5616 1476 5634 1494
rect 5616 1494 5634 1512
rect 5616 1512 5634 1530
rect 5616 1530 5634 1548
rect 5616 1548 5634 1566
rect 5616 1566 5634 1584
rect 5616 1584 5634 1602
rect 5616 1602 5634 1620
rect 5616 1620 5634 1638
rect 5616 1638 5634 1656
rect 5616 1656 5634 1674
rect 5616 1674 5634 1692
rect 5616 1692 5634 1710
rect 5616 1710 5634 1728
rect 5616 1728 5634 1746
rect 5616 1746 5634 1764
rect 5616 1764 5634 1782
rect 5616 1782 5634 1800
rect 5616 1800 5634 1818
rect 5616 1818 5634 1836
rect 5616 1836 5634 1854
rect 5616 1854 5634 1872
rect 5616 1872 5634 1890
rect 5616 1890 5634 1908
rect 5616 1908 5634 1926
rect 5616 1926 5634 1944
rect 5616 1944 5634 1962
rect 5616 1962 5634 1980
rect 5616 1980 5634 1998
rect 5616 1998 5634 2016
rect 5616 2016 5634 2034
rect 5616 2034 5634 2052
rect 5616 2052 5634 2070
rect 5616 2070 5634 2088
rect 5616 2088 5634 2106
rect 5616 2106 5634 2124
rect 5616 2124 5634 2142
rect 5616 2142 5634 2160
rect 5616 2160 5634 2178
rect 5616 2178 5634 2196
rect 5616 2196 5634 2214
rect 5616 2214 5634 2232
rect 5616 2232 5634 2250
rect 5616 2250 5634 2268
rect 5616 2268 5634 2286
rect 5616 2286 5634 2304
rect 5616 2304 5634 2322
rect 5616 2322 5634 2340
rect 5616 2340 5634 2358
rect 5616 2358 5634 2376
rect 5616 2376 5634 2394
rect 5616 2394 5634 2412
rect 5616 2412 5634 2430
rect 5616 2430 5634 2448
rect 5616 2448 5634 2466
rect 5616 2466 5634 2484
rect 5616 2484 5634 2502
rect 5616 2502 5634 2520
rect 5616 2520 5634 2538
rect 5616 2538 5634 2556
rect 5616 2556 5634 2574
rect 5616 2790 5634 2808
rect 5616 2808 5634 2826
rect 5616 2826 5634 2844
rect 5616 2844 5634 2862
rect 5616 2862 5634 2880
rect 5616 2880 5634 2898
rect 5616 2898 5634 2916
rect 5616 2916 5634 2934
rect 5616 2934 5634 2952
rect 5616 2952 5634 2970
rect 5616 2970 5634 2988
rect 5616 2988 5634 3006
rect 5616 3006 5634 3024
rect 5616 3024 5634 3042
rect 5616 3042 5634 3060
rect 5616 3060 5634 3078
rect 5616 3078 5634 3096
rect 5616 3096 5634 3114
rect 5616 3114 5634 3132
rect 5616 3132 5634 3150
rect 5616 3150 5634 3168
rect 5616 3168 5634 3186
rect 5616 3186 5634 3204
rect 5616 3204 5634 3222
rect 5616 3222 5634 3240
rect 5616 3240 5634 3258
rect 5616 3258 5634 3276
rect 5616 3276 5634 3294
rect 5616 3294 5634 3312
rect 5616 3312 5634 3330
rect 5616 3330 5634 3348
rect 5616 3348 5634 3366
rect 5616 3366 5634 3384
rect 5616 3384 5634 3402
rect 5616 3402 5634 3420
rect 5616 3420 5634 3438
rect 5616 3438 5634 3456
rect 5616 3456 5634 3474
rect 5616 3474 5634 3492
rect 5616 3492 5634 3510
rect 5616 3510 5634 3528
rect 5616 3528 5634 3546
rect 5616 3546 5634 3564
rect 5616 3564 5634 3582
rect 5616 3582 5634 3600
rect 5616 3600 5634 3618
rect 5616 3618 5634 3636
rect 5616 3636 5634 3654
rect 5616 3654 5634 3672
rect 5616 3672 5634 3690
rect 5616 3690 5634 3708
rect 5616 3708 5634 3726
rect 5616 3726 5634 3744
rect 5616 3744 5634 3762
rect 5616 3762 5634 3780
rect 5616 3780 5634 3798
rect 5616 3798 5634 3816
rect 5616 3816 5634 3834
rect 5616 3834 5634 3852
rect 5616 3852 5634 3870
rect 5616 3870 5634 3888
rect 5616 3888 5634 3906
rect 5616 3906 5634 3924
rect 5616 3924 5634 3942
rect 5616 3942 5634 3960
rect 5616 3960 5634 3978
rect 5616 3978 5634 3996
rect 5616 3996 5634 4014
rect 5616 4014 5634 4032
rect 5616 4032 5634 4050
rect 5616 4050 5634 4068
rect 5616 4068 5634 4086
rect 5616 4086 5634 4104
rect 5616 4104 5634 4122
rect 5616 4122 5634 4140
rect 5616 4140 5634 4158
rect 5616 4158 5634 4176
rect 5616 4176 5634 4194
rect 5616 4194 5634 4212
rect 5616 4212 5634 4230
rect 5616 4230 5634 4248
rect 5616 4248 5634 4266
rect 5616 4266 5634 4284
rect 5616 4284 5634 4302
rect 5616 4302 5634 4320
rect 5616 4320 5634 4338
rect 5616 4338 5634 4356
rect 5616 4356 5634 4374
rect 5616 4374 5634 4392
rect 5616 4392 5634 4410
rect 5616 4410 5634 4428
rect 5616 4428 5634 4446
rect 5616 4446 5634 4464
rect 5616 4464 5634 4482
rect 5616 4482 5634 4500
rect 5616 4500 5634 4518
rect 5616 4518 5634 4536
rect 5616 4536 5634 4554
rect 5616 4554 5634 4572
rect 5616 4572 5634 4590
rect 5616 4590 5634 4608
rect 5616 4608 5634 4626
rect 5616 4626 5634 4644
rect 5616 4644 5634 4662
rect 5616 4662 5634 4680
rect 5616 4680 5634 4698
rect 5616 4698 5634 4716
rect 5616 4716 5634 4734
rect 5616 4734 5634 4752
rect 5616 4752 5634 4770
rect 5616 4770 5634 4788
rect 5616 4788 5634 4806
rect 5616 4806 5634 4824
rect 5616 4824 5634 4842
rect 5616 4842 5634 4860
rect 5616 4860 5634 4878
rect 5616 4878 5634 4896
rect 5616 4896 5634 4914
rect 5616 4914 5634 4932
rect 5616 4932 5634 4950
rect 5616 4950 5634 4968
rect 5616 4968 5634 4986
rect 5616 4986 5634 5004
rect 5616 5004 5634 5022
rect 5616 5238 5634 5256
rect 5616 5256 5634 5274
rect 5616 5274 5634 5292
rect 5616 5292 5634 5310
rect 5616 5310 5634 5328
rect 5616 5328 5634 5346
rect 5616 5346 5634 5364
rect 5616 5364 5634 5382
rect 5616 5382 5634 5400
rect 5616 5400 5634 5418
rect 5616 5418 5634 5436
rect 5616 5436 5634 5454
rect 5616 5454 5634 5472
rect 5616 5472 5634 5490
rect 5616 5490 5634 5508
rect 5616 5508 5634 5526
rect 5616 5526 5634 5544
rect 5616 5544 5634 5562
rect 5616 5562 5634 5580
rect 5616 5580 5634 5598
rect 5616 5598 5634 5616
rect 5616 5616 5634 5634
rect 5616 5634 5634 5652
rect 5616 5652 5634 5670
rect 5616 5670 5634 5688
rect 5616 5688 5634 5706
rect 5616 5706 5634 5724
rect 5616 5724 5634 5742
rect 5616 5742 5634 5760
rect 5616 5760 5634 5778
rect 5616 5778 5634 5796
rect 5616 5796 5634 5814
rect 5616 5814 5634 5832
rect 5616 5832 5634 5850
rect 5616 5850 5634 5868
rect 5616 5868 5634 5886
rect 5616 5886 5634 5904
rect 5616 5904 5634 5922
rect 5616 5922 5634 5940
rect 5616 5940 5634 5958
rect 5616 5958 5634 5976
rect 5616 5976 5634 5994
rect 5616 5994 5634 6012
rect 5616 6012 5634 6030
rect 5616 6030 5634 6048
rect 5616 6048 5634 6066
rect 5616 6066 5634 6084
rect 5616 6084 5634 6102
rect 5616 6102 5634 6120
rect 5616 6120 5634 6138
rect 5616 6138 5634 6156
rect 5616 6156 5634 6174
rect 5616 6174 5634 6192
rect 5616 6192 5634 6210
rect 5616 6210 5634 6228
rect 5616 6228 5634 6246
rect 5616 6246 5634 6264
rect 5616 6264 5634 6282
rect 5616 6282 5634 6300
rect 5616 6300 5634 6318
rect 5616 6318 5634 6336
rect 5616 6336 5634 6354
rect 5616 6354 5634 6372
rect 5616 6372 5634 6390
rect 5616 6390 5634 6408
rect 5616 6408 5634 6426
rect 5616 6426 5634 6444
rect 5616 6444 5634 6462
rect 5616 6462 5634 6480
rect 5616 6480 5634 6498
rect 5616 6498 5634 6516
rect 5616 6516 5634 6534
rect 5616 6534 5634 6552
rect 5616 6552 5634 6570
rect 5616 6570 5634 6588
rect 5616 6588 5634 6606
rect 5616 6606 5634 6624
rect 5616 6624 5634 6642
rect 5616 6642 5634 6660
rect 5616 6660 5634 6678
rect 5616 6678 5634 6696
rect 5616 6696 5634 6714
rect 5616 6714 5634 6732
rect 5616 6732 5634 6750
rect 5616 6750 5634 6768
rect 5616 6768 5634 6786
rect 5616 6786 5634 6804
rect 5616 6804 5634 6822
rect 5616 6822 5634 6840
rect 5616 6840 5634 6858
rect 5616 6858 5634 6876
rect 5616 6876 5634 6894
rect 5616 6894 5634 6912
rect 5616 6912 5634 6930
rect 5616 6930 5634 6948
rect 5616 6948 5634 6966
rect 5616 6966 5634 6984
rect 5616 6984 5634 7002
rect 5616 7002 5634 7020
rect 5616 7020 5634 7038
rect 5616 7038 5634 7056
rect 5616 7056 5634 7074
rect 5616 7074 5634 7092
rect 5616 7092 5634 7110
rect 5616 7110 5634 7128
rect 5616 7128 5634 7146
rect 5616 7146 5634 7164
rect 5616 7164 5634 7182
rect 5616 7182 5634 7200
rect 5616 7200 5634 7218
rect 5616 7218 5634 7236
rect 5616 7236 5634 7254
rect 5616 7254 5634 7272
rect 5616 7272 5634 7290
rect 5616 7290 5634 7308
rect 5616 7308 5634 7326
rect 5616 7326 5634 7344
rect 5616 7344 5634 7362
rect 5616 7362 5634 7380
rect 5616 7380 5634 7398
rect 5616 7398 5634 7416
rect 5616 7416 5634 7434
rect 5616 7434 5634 7452
rect 5616 7452 5634 7470
rect 5616 7470 5634 7488
rect 5616 7488 5634 7506
rect 5616 7506 5634 7524
rect 5616 7524 5634 7542
rect 5616 7542 5634 7560
rect 5616 7560 5634 7578
rect 5616 7578 5634 7596
rect 5616 7596 5634 7614
rect 5616 7614 5634 7632
rect 5616 7632 5634 7650
rect 5616 7650 5634 7668
rect 5616 7668 5634 7686
rect 5616 7686 5634 7704
rect 5616 7704 5634 7722
rect 5616 7722 5634 7740
rect 5616 7740 5634 7758
rect 5616 7758 5634 7776
rect 5616 7776 5634 7794
rect 5616 7794 5634 7812
rect 5616 7812 5634 7830
rect 5616 7830 5634 7848
rect 5616 7848 5634 7866
rect 5616 7866 5634 7884
rect 5616 7884 5634 7902
rect 5616 7902 5634 7920
rect 5616 7920 5634 7938
rect 5616 7938 5634 7956
rect 5616 7956 5634 7974
rect 5616 7974 5634 7992
rect 5616 7992 5634 8010
rect 5616 8010 5634 8028
rect 5616 8028 5634 8046
rect 5616 8046 5634 8064
rect 5616 8064 5634 8082
rect 5616 8082 5634 8100
rect 5616 8100 5634 8118
rect 5616 8118 5634 8136
rect 5616 8136 5634 8154
rect 5616 8154 5634 8172
rect 5616 8172 5634 8190
rect 5616 8190 5634 8208
rect 5616 8208 5634 8226
rect 5616 8226 5634 8244
rect 5616 8244 5634 8262
rect 5616 8262 5634 8280
rect 5616 8280 5634 8298
rect 5616 8298 5634 8316
rect 5616 8316 5634 8334
rect 5616 8334 5634 8352
rect 5616 8352 5634 8370
rect 5616 8370 5634 8388
rect 5616 8388 5634 8406
rect 5616 8406 5634 8424
rect 5616 8424 5634 8442
rect 5616 8442 5634 8460
rect 5616 8460 5634 8478
rect 5616 8478 5634 8496
rect 5616 8496 5634 8514
rect 5616 8514 5634 8532
rect 5616 8532 5634 8550
rect 5616 8550 5634 8568
rect 5616 8568 5634 8586
rect 5616 8586 5634 8604
rect 5616 8604 5634 8622
rect 5616 8622 5634 8640
rect 5616 8640 5634 8658
rect 5616 8658 5634 8676
rect 5616 8676 5634 8694
rect 5616 8694 5634 8712
rect 5616 8712 5634 8730
rect 5634 612 5652 630
rect 5634 630 5652 648
rect 5634 648 5652 666
rect 5634 666 5652 684
rect 5634 684 5652 702
rect 5634 702 5652 720
rect 5634 720 5652 738
rect 5634 738 5652 756
rect 5634 756 5652 774
rect 5634 774 5652 792
rect 5634 792 5652 810
rect 5634 810 5652 828
rect 5634 828 5652 846
rect 5634 846 5652 864
rect 5634 864 5652 882
rect 5634 882 5652 900
rect 5634 900 5652 918
rect 5634 918 5652 936
rect 5634 936 5652 954
rect 5634 954 5652 972
rect 5634 1116 5652 1134
rect 5634 1134 5652 1152
rect 5634 1152 5652 1170
rect 5634 1170 5652 1188
rect 5634 1188 5652 1206
rect 5634 1206 5652 1224
rect 5634 1224 5652 1242
rect 5634 1242 5652 1260
rect 5634 1260 5652 1278
rect 5634 1278 5652 1296
rect 5634 1296 5652 1314
rect 5634 1314 5652 1332
rect 5634 1332 5652 1350
rect 5634 1350 5652 1368
rect 5634 1368 5652 1386
rect 5634 1386 5652 1404
rect 5634 1404 5652 1422
rect 5634 1422 5652 1440
rect 5634 1440 5652 1458
rect 5634 1458 5652 1476
rect 5634 1476 5652 1494
rect 5634 1494 5652 1512
rect 5634 1512 5652 1530
rect 5634 1530 5652 1548
rect 5634 1548 5652 1566
rect 5634 1566 5652 1584
rect 5634 1584 5652 1602
rect 5634 1602 5652 1620
rect 5634 1620 5652 1638
rect 5634 1638 5652 1656
rect 5634 1656 5652 1674
rect 5634 1674 5652 1692
rect 5634 1692 5652 1710
rect 5634 1710 5652 1728
rect 5634 1728 5652 1746
rect 5634 1746 5652 1764
rect 5634 1764 5652 1782
rect 5634 1782 5652 1800
rect 5634 1800 5652 1818
rect 5634 1818 5652 1836
rect 5634 1836 5652 1854
rect 5634 1854 5652 1872
rect 5634 1872 5652 1890
rect 5634 1890 5652 1908
rect 5634 1908 5652 1926
rect 5634 1926 5652 1944
rect 5634 1944 5652 1962
rect 5634 1962 5652 1980
rect 5634 1980 5652 1998
rect 5634 1998 5652 2016
rect 5634 2016 5652 2034
rect 5634 2034 5652 2052
rect 5634 2052 5652 2070
rect 5634 2070 5652 2088
rect 5634 2088 5652 2106
rect 5634 2106 5652 2124
rect 5634 2124 5652 2142
rect 5634 2142 5652 2160
rect 5634 2160 5652 2178
rect 5634 2178 5652 2196
rect 5634 2196 5652 2214
rect 5634 2214 5652 2232
rect 5634 2232 5652 2250
rect 5634 2250 5652 2268
rect 5634 2268 5652 2286
rect 5634 2286 5652 2304
rect 5634 2304 5652 2322
rect 5634 2322 5652 2340
rect 5634 2340 5652 2358
rect 5634 2358 5652 2376
rect 5634 2376 5652 2394
rect 5634 2394 5652 2412
rect 5634 2412 5652 2430
rect 5634 2430 5652 2448
rect 5634 2448 5652 2466
rect 5634 2466 5652 2484
rect 5634 2484 5652 2502
rect 5634 2502 5652 2520
rect 5634 2520 5652 2538
rect 5634 2538 5652 2556
rect 5634 2556 5652 2574
rect 5634 2574 5652 2592
rect 5634 2790 5652 2808
rect 5634 2808 5652 2826
rect 5634 2826 5652 2844
rect 5634 2844 5652 2862
rect 5634 2862 5652 2880
rect 5634 2880 5652 2898
rect 5634 2898 5652 2916
rect 5634 2916 5652 2934
rect 5634 2934 5652 2952
rect 5634 2952 5652 2970
rect 5634 2970 5652 2988
rect 5634 2988 5652 3006
rect 5634 3006 5652 3024
rect 5634 3024 5652 3042
rect 5634 3042 5652 3060
rect 5634 3060 5652 3078
rect 5634 3078 5652 3096
rect 5634 3096 5652 3114
rect 5634 3114 5652 3132
rect 5634 3132 5652 3150
rect 5634 3150 5652 3168
rect 5634 3168 5652 3186
rect 5634 3186 5652 3204
rect 5634 3204 5652 3222
rect 5634 3222 5652 3240
rect 5634 3240 5652 3258
rect 5634 3258 5652 3276
rect 5634 3276 5652 3294
rect 5634 3294 5652 3312
rect 5634 3312 5652 3330
rect 5634 3330 5652 3348
rect 5634 3348 5652 3366
rect 5634 3366 5652 3384
rect 5634 3384 5652 3402
rect 5634 3402 5652 3420
rect 5634 3420 5652 3438
rect 5634 3438 5652 3456
rect 5634 3456 5652 3474
rect 5634 3474 5652 3492
rect 5634 3492 5652 3510
rect 5634 3510 5652 3528
rect 5634 3528 5652 3546
rect 5634 3546 5652 3564
rect 5634 3564 5652 3582
rect 5634 3582 5652 3600
rect 5634 3600 5652 3618
rect 5634 3618 5652 3636
rect 5634 3636 5652 3654
rect 5634 3654 5652 3672
rect 5634 3672 5652 3690
rect 5634 3690 5652 3708
rect 5634 3708 5652 3726
rect 5634 3726 5652 3744
rect 5634 3744 5652 3762
rect 5634 3762 5652 3780
rect 5634 3780 5652 3798
rect 5634 3798 5652 3816
rect 5634 3816 5652 3834
rect 5634 3834 5652 3852
rect 5634 3852 5652 3870
rect 5634 3870 5652 3888
rect 5634 3888 5652 3906
rect 5634 3906 5652 3924
rect 5634 3924 5652 3942
rect 5634 3942 5652 3960
rect 5634 3960 5652 3978
rect 5634 3978 5652 3996
rect 5634 3996 5652 4014
rect 5634 4014 5652 4032
rect 5634 4032 5652 4050
rect 5634 4050 5652 4068
rect 5634 4068 5652 4086
rect 5634 4086 5652 4104
rect 5634 4104 5652 4122
rect 5634 4122 5652 4140
rect 5634 4140 5652 4158
rect 5634 4158 5652 4176
rect 5634 4176 5652 4194
rect 5634 4194 5652 4212
rect 5634 4212 5652 4230
rect 5634 4230 5652 4248
rect 5634 4248 5652 4266
rect 5634 4266 5652 4284
rect 5634 4284 5652 4302
rect 5634 4302 5652 4320
rect 5634 4320 5652 4338
rect 5634 4338 5652 4356
rect 5634 4356 5652 4374
rect 5634 4374 5652 4392
rect 5634 4392 5652 4410
rect 5634 4410 5652 4428
rect 5634 4428 5652 4446
rect 5634 4446 5652 4464
rect 5634 4464 5652 4482
rect 5634 4482 5652 4500
rect 5634 4500 5652 4518
rect 5634 4518 5652 4536
rect 5634 4536 5652 4554
rect 5634 4554 5652 4572
rect 5634 4572 5652 4590
rect 5634 4590 5652 4608
rect 5634 4608 5652 4626
rect 5634 4626 5652 4644
rect 5634 4644 5652 4662
rect 5634 4662 5652 4680
rect 5634 4680 5652 4698
rect 5634 4698 5652 4716
rect 5634 4716 5652 4734
rect 5634 4734 5652 4752
rect 5634 4752 5652 4770
rect 5634 4770 5652 4788
rect 5634 4788 5652 4806
rect 5634 4806 5652 4824
rect 5634 4824 5652 4842
rect 5634 4842 5652 4860
rect 5634 4860 5652 4878
rect 5634 4878 5652 4896
rect 5634 4896 5652 4914
rect 5634 4914 5652 4932
rect 5634 4932 5652 4950
rect 5634 4950 5652 4968
rect 5634 4968 5652 4986
rect 5634 4986 5652 5004
rect 5634 5004 5652 5022
rect 5634 5022 5652 5040
rect 5634 5256 5652 5274
rect 5634 5274 5652 5292
rect 5634 5292 5652 5310
rect 5634 5310 5652 5328
rect 5634 5328 5652 5346
rect 5634 5346 5652 5364
rect 5634 5364 5652 5382
rect 5634 5382 5652 5400
rect 5634 5400 5652 5418
rect 5634 5418 5652 5436
rect 5634 5436 5652 5454
rect 5634 5454 5652 5472
rect 5634 5472 5652 5490
rect 5634 5490 5652 5508
rect 5634 5508 5652 5526
rect 5634 5526 5652 5544
rect 5634 5544 5652 5562
rect 5634 5562 5652 5580
rect 5634 5580 5652 5598
rect 5634 5598 5652 5616
rect 5634 5616 5652 5634
rect 5634 5634 5652 5652
rect 5634 5652 5652 5670
rect 5634 5670 5652 5688
rect 5634 5688 5652 5706
rect 5634 5706 5652 5724
rect 5634 5724 5652 5742
rect 5634 5742 5652 5760
rect 5634 5760 5652 5778
rect 5634 5778 5652 5796
rect 5634 5796 5652 5814
rect 5634 5814 5652 5832
rect 5634 5832 5652 5850
rect 5634 5850 5652 5868
rect 5634 5868 5652 5886
rect 5634 5886 5652 5904
rect 5634 5904 5652 5922
rect 5634 5922 5652 5940
rect 5634 5940 5652 5958
rect 5634 5958 5652 5976
rect 5634 5976 5652 5994
rect 5634 5994 5652 6012
rect 5634 6012 5652 6030
rect 5634 6030 5652 6048
rect 5634 6048 5652 6066
rect 5634 6066 5652 6084
rect 5634 6084 5652 6102
rect 5634 6102 5652 6120
rect 5634 6120 5652 6138
rect 5634 6138 5652 6156
rect 5634 6156 5652 6174
rect 5634 6174 5652 6192
rect 5634 6192 5652 6210
rect 5634 6210 5652 6228
rect 5634 6228 5652 6246
rect 5634 6246 5652 6264
rect 5634 6264 5652 6282
rect 5634 6282 5652 6300
rect 5634 6300 5652 6318
rect 5634 6318 5652 6336
rect 5634 6336 5652 6354
rect 5634 6354 5652 6372
rect 5634 6372 5652 6390
rect 5634 6390 5652 6408
rect 5634 6408 5652 6426
rect 5634 6426 5652 6444
rect 5634 6444 5652 6462
rect 5634 6462 5652 6480
rect 5634 6480 5652 6498
rect 5634 6498 5652 6516
rect 5634 6516 5652 6534
rect 5634 6534 5652 6552
rect 5634 6552 5652 6570
rect 5634 6570 5652 6588
rect 5634 6588 5652 6606
rect 5634 6606 5652 6624
rect 5634 6624 5652 6642
rect 5634 6642 5652 6660
rect 5634 6660 5652 6678
rect 5634 6678 5652 6696
rect 5634 6696 5652 6714
rect 5634 6714 5652 6732
rect 5634 6732 5652 6750
rect 5634 6750 5652 6768
rect 5634 6768 5652 6786
rect 5634 6786 5652 6804
rect 5634 6804 5652 6822
rect 5634 6822 5652 6840
rect 5634 6840 5652 6858
rect 5634 6858 5652 6876
rect 5634 6876 5652 6894
rect 5634 6894 5652 6912
rect 5634 6912 5652 6930
rect 5634 6930 5652 6948
rect 5634 6948 5652 6966
rect 5634 6966 5652 6984
rect 5634 6984 5652 7002
rect 5634 7002 5652 7020
rect 5634 7020 5652 7038
rect 5634 7038 5652 7056
rect 5634 7056 5652 7074
rect 5634 7074 5652 7092
rect 5634 7092 5652 7110
rect 5634 7110 5652 7128
rect 5634 7128 5652 7146
rect 5634 7146 5652 7164
rect 5634 7164 5652 7182
rect 5634 7182 5652 7200
rect 5634 7200 5652 7218
rect 5634 7218 5652 7236
rect 5634 7236 5652 7254
rect 5634 7254 5652 7272
rect 5634 7272 5652 7290
rect 5634 7290 5652 7308
rect 5634 7308 5652 7326
rect 5634 7326 5652 7344
rect 5634 7344 5652 7362
rect 5634 7362 5652 7380
rect 5634 7380 5652 7398
rect 5634 7398 5652 7416
rect 5634 7416 5652 7434
rect 5634 7434 5652 7452
rect 5634 7452 5652 7470
rect 5634 7470 5652 7488
rect 5634 7488 5652 7506
rect 5634 7506 5652 7524
rect 5634 7524 5652 7542
rect 5634 7542 5652 7560
rect 5634 7560 5652 7578
rect 5634 7578 5652 7596
rect 5634 7596 5652 7614
rect 5634 7614 5652 7632
rect 5634 7632 5652 7650
rect 5634 7650 5652 7668
rect 5634 7668 5652 7686
rect 5634 7686 5652 7704
rect 5634 7704 5652 7722
rect 5634 7722 5652 7740
rect 5634 7740 5652 7758
rect 5634 7758 5652 7776
rect 5634 7776 5652 7794
rect 5634 7794 5652 7812
rect 5634 7812 5652 7830
rect 5634 7830 5652 7848
rect 5634 7848 5652 7866
rect 5634 7866 5652 7884
rect 5634 7884 5652 7902
rect 5634 7902 5652 7920
rect 5634 7920 5652 7938
rect 5634 7938 5652 7956
rect 5634 7956 5652 7974
rect 5634 7974 5652 7992
rect 5634 7992 5652 8010
rect 5634 8010 5652 8028
rect 5634 8028 5652 8046
rect 5634 8046 5652 8064
rect 5634 8064 5652 8082
rect 5634 8082 5652 8100
rect 5634 8100 5652 8118
rect 5634 8118 5652 8136
rect 5634 8136 5652 8154
rect 5634 8154 5652 8172
rect 5634 8172 5652 8190
rect 5634 8190 5652 8208
rect 5634 8208 5652 8226
rect 5634 8226 5652 8244
rect 5634 8244 5652 8262
rect 5634 8262 5652 8280
rect 5634 8280 5652 8298
rect 5634 8298 5652 8316
rect 5634 8316 5652 8334
rect 5634 8334 5652 8352
rect 5634 8352 5652 8370
rect 5634 8370 5652 8388
rect 5634 8388 5652 8406
rect 5634 8406 5652 8424
rect 5634 8424 5652 8442
rect 5634 8442 5652 8460
rect 5634 8460 5652 8478
rect 5634 8478 5652 8496
rect 5634 8496 5652 8514
rect 5634 8514 5652 8532
rect 5634 8532 5652 8550
rect 5634 8550 5652 8568
rect 5634 8568 5652 8586
rect 5634 8586 5652 8604
rect 5634 8604 5652 8622
rect 5634 8622 5652 8640
rect 5634 8640 5652 8658
rect 5634 8658 5652 8676
rect 5634 8676 5652 8694
rect 5634 8694 5652 8712
rect 5634 8712 5652 8730
rect 5634 8730 5652 8748
rect 5652 630 5670 648
rect 5652 648 5670 666
rect 5652 666 5670 684
rect 5652 684 5670 702
rect 5652 702 5670 720
rect 5652 720 5670 738
rect 5652 738 5670 756
rect 5652 756 5670 774
rect 5652 774 5670 792
rect 5652 792 5670 810
rect 5652 810 5670 828
rect 5652 828 5670 846
rect 5652 846 5670 864
rect 5652 864 5670 882
rect 5652 882 5670 900
rect 5652 900 5670 918
rect 5652 918 5670 936
rect 5652 936 5670 954
rect 5652 954 5670 972
rect 5652 1116 5670 1134
rect 5652 1134 5670 1152
rect 5652 1152 5670 1170
rect 5652 1170 5670 1188
rect 5652 1188 5670 1206
rect 5652 1206 5670 1224
rect 5652 1224 5670 1242
rect 5652 1242 5670 1260
rect 5652 1260 5670 1278
rect 5652 1278 5670 1296
rect 5652 1296 5670 1314
rect 5652 1314 5670 1332
rect 5652 1332 5670 1350
rect 5652 1350 5670 1368
rect 5652 1368 5670 1386
rect 5652 1386 5670 1404
rect 5652 1404 5670 1422
rect 5652 1422 5670 1440
rect 5652 1440 5670 1458
rect 5652 1458 5670 1476
rect 5652 1476 5670 1494
rect 5652 1494 5670 1512
rect 5652 1512 5670 1530
rect 5652 1530 5670 1548
rect 5652 1548 5670 1566
rect 5652 1566 5670 1584
rect 5652 1584 5670 1602
rect 5652 1602 5670 1620
rect 5652 1620 5670 1638
rect 5652 1638 5670 1656
rect 5652 1656 5670 1674
rect 5652 1674 5670 1692
rect 5652 1692 5670 1710
rect 5652 1710 5670 1728
rect 5652 1728 5670 1746
rect 5652 1746 5670 1764
rect 5652 1764 5670 1782
rect 5652 1782 5670 1800
rect 5652 1800 5670 1818
rect 5652 1818 5670 1836
rect 5652 1836 5670 1854
rect 5652 1854 5670 1872
rect 5652 1872 5670 1890
rect 5652 1890 5670 1908
rect 5652 1908 5670 1926
rect 5652 1926 5670 1944
rect 5652 1944 5670 1962
rect 5652 1962 5670 1980
rect 5652 1980 5670 1998
rect 5652 1998 5670 2016
rect 5652 2016 5670 2034
rect 5652 2034 5670 2052
rect 5652 2052 5670 2070
rect 5652 2070 5670 2088
rect 5652 2088 5670 2106
rect 5652 2106 5670 2124
rect 5652 2124 5670 2142
rect 5652 2142 5670 2160
rect 5652 2160 5670 2178
rect 5652 2178 5670 2196
rect 5652 2196 5670 2214
rect 5652 2214 5670 2232
rect 5652 2232 5670 2250
rect 5652 2250 5670 2268
rect 5652 2268 5670 2286
rect 5652 2286 5670 2304
rect 5652 2304 5670 2322
rect 5652 2322 5670 2340
rect 5652 2340 5670 2358
rect 5652 2358 5670 2376
rect 5652 2376 5670 2394
rect 5652 2394 5670 2412
rect 5652 2412 5670 2430
rect 5652 2430 5670 2448
rect 5652 2448 5670 2466
rect 5652 2466 5670 2484
rect 5652 2484 5670 2502
rect 5652 2502 5670 2520
rect 5652 2520 5670 2538
rect 5652 2538 5670 2556
rect 5652 2556 5670 2574
rect 5652 2574 5670 2592
rect 5652 2808 5670 2826
rect 5652 2826 5670 2844
rect 5652 2844 5670 2862
rect 5652 2862 5670 2880
rect 5652 2880 5670 2898
rect 5652 2898 5670 2916
rect 5652 2916 5670 2934
rect 5652 2934 5670 2952
rect 5652 2952 5670 2970
rect 5652 2970 5670 2988
rect 5652 2988 5670 3006
rect 5652 3006 5670 3024
rect 5652 3024 5670 3042
rect 5652 3042 5670 3060
rect 5652 3060 5670 3078
rect 5652 3078 5670 3096
rect 5652 3096 5670 3114
rect 5652 3114 5670 3132
rect 5652 3132 5670 3150
rect 5652 3150 5670 3168
rect 5652 3168 5670 3186
rect 5652 3186 5670 3204
rect 5652 3204 5670 3222
rect 5652 3222 5670 3240
rect 5652 3240 5670 3258
rect 5652 3258 5670 3276
rect 5652 3276 5670 3294
rect 5652 3294 5670 3312
rect 5652 3312 5670 3330
rect 5652 3330 5670 3348
rect 5652 3348 5670 3366
rect 5652 3366 5670 3384
rect 5652 3384 5670 3402
rect 5652 3402 5670 3420
rect 5652 3420 5670 3438
rect 5652 3438 5670 3456
rect 5652 3456 5670 3474
rect 5652 3474 5670 3492
rect 5652 3492 5670 3510
rect 5652 3510 5670 3528
rect 5652 3528 5670 3546
rect 5652 3546 5670 3564
rect 5652 3564 5670 3582
rect 5652 3582 5670 3600
rect 5652 3600 5670 3618
rect 5652 3618 5670 3636
rect 5652 3636 5670 3654
rect 5652 3654 5670 3672
rect 5652 3672 5670 3690
rect 5652 3690 5670 3708
rect 5652 3708 5670 3726
rect 5652 3726 5670 3744
rect 5652 3744 5670 3762
rect 5652 3762 5670 3780
rect 5652 3780 5670 3798
rect 5652 3798 5670 3816
rect 5652 3816 5670 3834
rect 5652 3834 5670 3852
rect 5652 3852 5670 3870
rect 5652 3870 5670 3888
rect 5652 3888 5670 3906
rect 5652 3906 5670 3924
rect 5652 3924 5670 3942
rect 5652 3942 5670 3960
rect 5652 3960 5670 3978
rect 5652 3978 5670 3996
rect 5652 3996 5670 4014
rect 5652 4014 5670 4032
rect 5652 4032 5670 4050
rect 5652 4050 5670 4068
rect 5652 4068 5670 4086
rect 5652 4086 5670 4104
rect 5652 4104 5670 4122
rect 5652 4122 5670 4140
rect 5652 4140 5670 4158
rect 5652 4158 5670 4176
rect 5652 4176 5670 4194
rect 5652 4194 5670 4212
rect 5652 4212 5670 4230
rect 5652 4230 5670 4248
rect 5652 4248 5670 4266
rect 5652 4266 5670 4284
rect 5652 4284 5670 4302
rect 5652 4302 5670 4320
rect 5652 4320 5670 4338
rect 5652 4338 5670 4356
rect 5652 4356 5670 4374
rect 5652 4374 5670 4392
rect 5652 4392 5670 4410
rect 5652 4410 5670 4428
rect 5652 4428 5670 4446
rect 5652 4446 5670 4464
rect 5652 4464 5670 4482
rect 5652 4482 5670 4500
rect 5652 4500 5670 4518
rect 5652 4518 5670 4536
rect 5652 4536 5670 4554
rect 5652 4554 5670 4572
rect 5652 4572 5670 4590
rect 5652 4590 5670 4608
rect 5652 4608 5670 4626
rect 5652 4626 5670 4644
rect 5652 4644 5670 4662
rect 5652 4662 5670 4680
rect 5652 4680 5670 4698
rect 5652 4698 5670 4716
rect 5652 4716 5670 4734
rect 5652 4734 5670 4752
rect 5652 4752 5670 4770
rect 5652 4770 5670 4788
rect 5652 4788 5670 4806
rect 5652 4806 5670 4824
rect 5652 4824 5670 4842
rect 5652 4842 5670 4860
rect 5652 4860 5670 4878
rect 5652 4878 5670 4896
rect 5652 4896 5670 4914
rect 5652 4914 5670 4932
rect 5652 4932 5670 4950
rect 5652 4950 5670 4968
rect 5652 4968 5670 4986
rect 5652 4986 5670 5004
rect 5652 5004 5670 5022
rect 5652 5022 5670 5040
rect 5652 5040 5670 5058
rect 5652 5274 5670 5292
rect 5652 5292 5670 5310
rect 5652 5310 5670 5328
rect 5652 5328 5670 5346
rect 5652 5346 5670 5364
rect 5652 5364 5670 5382
rect 5652 5382 5670 5400
rect 5652 5400 5670 5418
rect 5652 5418 5670 5436
rect 5652 5436 5670 5454
rect 5652 5454 5670 5472
rect 5652 5472 5670 5490
rect 5652 5490 5670 5508
rect 5652 5508 5670 5526
rect 5652 5526 5670 5544
rect 5652 5544 5670 5562
rect 5652 5562 5670 5580
rect 5652 5580 5670 5598
rect 5652 5598 5670 5616
rect 5652 5616 5670 5634
rect 5652 5634 5670 5652
rect 5652 5652 5670 5670
rect 5652 5670 5670 5688
rect 5652 5688 5670 5706
rect 5652 5706 5670 5724
rect 5652 5724 5670 5742
rect 5652 5742 5670 5760
rect 5652 5760 5670 5778
rect 5652 5778 5670 5796
rect 5652 5796 5670 5814
rect 5652 5814 5670 5832
rect 5652 5832 5670 5850
rect 5652 5850 5670 5868
rect 5652 5868 5670 5886
rect 5652 5886 5670 5904
rect 5652 5904 5670 5922
rect 5652 5922 5670 5940
rect 5652 5940 5670 5958
rect 5652 5958 5670 5976
rect 5652 5976 5670 5994
rect 5652 5994 5670 6012
rect 5652 6012 5670 6030
rect 5652 6030 5670 6048
rect 5652 6048 5670 6066
rect 5652 6066 5670 6084
rect 5652 6084 5670 6102
rect 5652 6102 5670 6120
rect 5652 6120 5670 6138
rect 5652 6138 5670 6156
rect 5652 6156 5670 6174
rect 5652 6174 5670 6192
rect 5652 6192 5670 6210
rect 5652 6210 5670 6228
rect 5652 6228 5670 6246
rect 5652 6246 5670 6264
rect 5652 6264 5670 6282
rect 5652 6282 5670 6300
rect 5652 6300 5670 6318
rect 5652 6318 5670 6336
rect 5652 6336 5670 6354
rect 5652 6354 5670 6372
rect 5652 6372 5670 6390
rect 5652 6390 5670 6408
rect 5652 6408 5670 6426
rect 5652 6426 5670 6444
rect 5652 6444 5670 6462
rect 5652 6462 5670 6480
rect 5652 6480 5670 6498
rect 5652 6498 5670 6516
rect 5652 6516 5670 6534
rect 5652 6534 5670 6552
rect 5652 6552 5670 6570
rect 5652 6570 5670 6588
rect 5652 6588 5670 6606
rect 5652 6606 5670 6624
rect 5652 6624 5670 6642
rect 5652 6642 5670 6660
rect 5652 6660 5670 6678
rect 5652 6678 5670 6696
rect 5652 6696 5670 6714
rect 5652 6714 5670 6732
rect 5652 6732 5670 6750
rect 5652 6750 5670 6768
rect 5652 6768 5670 6786
rect 5652 6786 5670 6804
rect 5652 6804 5670 6822
rect 5652 6822 5670 6840
rect 5652 6840 5670 6858
rect 5652 6858 5670 6876
rect 5652 6876 5670 6894
rect 5652 6894 5670 6912
rect 5652 6912 5670 6930
rect 5652 6930 5670 6948
rect 5652 6948 5670 6966
rect 5652 6966 5670 6984
rect 5652 6984 5670 7002
rect 5652 7002 5670 7020
rect 5652 7020 5670 7038
rect 5652 7038 5670 7056
rect 5652 7056 5670 7074
rect 5652 7074 5670 7092
rect 5652 7092 5670 7110
rect 5652 7110 5670 7128
rect 5652 7128 5670 7146
rect 5652 7146 5670 7164
rect 5652 7164 5670 7182
rect 5652 7182 5670 7200
rect 5652 7200 5670 7218
rect 5652 7218 5670 7236
rect 5652 7236 5670 7254
rect 5652 7254 5670 7272
rect 5652 7272 5670 7290
rect 5652 7290 5670 7308
rect 5652 7308 5670 7326
rect 5652 7326 5670 7344
rect 5652 7344 5670 7362
rect 5652 7362 5670 7380
rect 5652 7380 5670 7398
rect 5652 7398 5670 7416
rect 5652 7416 5670 7434
rect 5652 7434 5670 7452
rect 5652 7452 5670 7470
rect 5652 7470 5670 7488
rect 5652 7488 5670 7506
rect 5652 7506 5670 7524
rect 5652 7524 5670 7542
rect 5652 7542 5670 7560
rect 5652 7560 5670 7578
rect 5652 7578 5670 7596
rect 5652 7596 5670 7614
rect 5652 7614 5670 7632
rect 5652 7632 5670 7650
rect 5652 7650 5670 7668
rect 5652 7668 5670 7686
rect 5652 7686 5670 7704
rect 5652 7704 5670 7722
rect 5652 7722 5670 7740
rect 5652 7740 5670 7758
rect 5652 7758 5670 7776
rect 5652 7776 5670 7794
rect 5652 7794 5670 7812
rect 5652 7812 5670 7830
rect 5652 7830 5670 7848
rect 5652 7848 5670 7866
rect 5652 7866 5670 7884
rect 5652 7884 5670 7902
rect 5652 7902 5670 7920
rect 5652 7920 5670 7938
rect 5652 7938 5670 7956
rect 5652 7956 5670 7974
rect 5652 7974 5670 7992
rect 5652 7992 5670 8010
rect 5652 8010 5670 8028
rect 5652 8028 5670 8046
rect 5652 8046 5670 8064
rect 5652 8064 5670 8082
rect 5652 8082 5670 8100
rect 5652 8100 5670 8118
rect 5652 8118 5670 8136
rect 5652 8136 5670 8154
rect 5652 8154 5670 8172
rect 5652 8172 5670 8190
rect 5652 8190 5670 8208
rect 5652 8208 5670 8226
rect 5652 8226 5670 8244
rect 5652 8244 5670 8262
rect 5652 8262 5670 8280
rect 5652 8280 5670 8298
rect 5652 8298 5670 8316
rect 5652 8316 5670 8334
rect 5652 8334 5670 8352
rect 5652 8352 5670 8370
rect 5652 8370 5670 8388
rect 5652 8388 5670 8406
rect 5652 8406 5670 8424
rect 5652 8424 5670 8442
rect 5652 8442 5670 8460
rect 5652 8460 5670 8478
rect 5652 8478 5670 8496
rect 5652 8496 5670 8514
rect 5652 8514 5670 8532
rect 5652 8532 5670 8550
rect 5652 8550 5670 8568
rect 5652 8568 5670 8586
rect 5652 8586 5670 8604
rect 5652 8604 5670 8622
rect 5652 8622 5670 8640
rect 5652 8640 5670 8658
rect 5652 8658 5670 8676
rect 5652 8676 5670 8694
rect 5652 8694 5670 8712
rect 5652 8712 5670 8730
rect 5652 8730 5670 8748
rect 5652 8748 5670 8766
rect 5670 630 5688 648
rect 5670 648 5688 666
rect 5670 666 5688 684
rect 5670 684 5688 702
rect 5670 702 5688 720
rect 5670 720 5688 738
rect 5670 738 5688 756
rect 5670 756 5688 774
rect 5670 774 5688 792
rect 5670 792 5688 810
rect 5670 810 5688 828
rect 5670 828 5688 846
rect 5670 846 5688 864
rect 5670 864 5688 882
rect 5670 882 5688 900
rect 5670 900 5688 918
rect 5670 918 5688 936
rect 5670 936 5688 954
rect 5670 954 5688 972
rect 5670 972 5688 990
rect 5670 1116 5688 1134
rect 5670 1134 5688 1152
rect 5670 1152 5688 1170
rect 5670 1170 5688 1188
rect 5670 1188 5688 1206
rect 5670 1206 5688 1224
rect 5670 1224 5688 1242
rect 5670 1242 5688 1260
rect 5670 1260 5688 1278
rect 5670 1278 5688 1296
rect 5670 1296 5688 1314
rect 5670 1314 5688 1332
rect 5670 1332 5688 1350
rect 5670 1350 5688 1368
rect 5670 1368 5688 1386
rect 5670 1386 5688 1404
rect 5670 1404 5688 1422
rect 5670 1422 5688 1440
rect 5670 1440 5688 1458
rect 5670 1458 5688 1476
rect 5670 1476 5688 1494
rect 5670 1494 5688 1512
rect 5670 1512 5688 1530
rect 5670 1530 5688 1548
rect 5670 1548 5688 1566
rect 5670 1566 5688 1584
rect 5670 1584 5688 1602
rect 5670 1602 5688 1620
rect 5670 1620 5688 1638
rect 5670 1638 5688 1656
rect 5670 1656 5688 1674
rect 5670 1674 5688 1692
rect 5670 1692 5688 1710
rect 5670 1710 5688 1728
rect 5670 1728 5688 1746
rect 5670 1746 5688 1764
rect 5670 1764 5688 1782
rect 5670 1782 5688 1800
rect 5670 1800 5688 1818
rect 5670 1818 5688 1836
rect 5670 1836 5688 1854
rect 5670 1854 5688 1872
rect 5670 1872 5688 1890
rect 5670 1890 5688 1908
rect 5670 1908 5688 1926
rect 5670 1926 5688 1944
rect 5670 1944 5688 1962
rect 5670 1962 5688 1980
rect 5670 1980 5688 1998
rect 5670 1998 5688 2016
rect 5670 2016 5688 2034
rect 5670 2034 5688 2052
rect 5670 2052 5688 2070
rect 5670 2070 5688 2088
rect 5670 2088 5688 2106
rect 5670 2106 5688 2124
rect 5670 2124 5688 2142
rect 5670 2142 5688 2160
rect 5670 2160 5688 2178
rect 5670 2178 5688 2196
rect 5670 2196 5688 2214
rect 5670 2214 5688 2232
rect 5670 2232 5688 2250
rect 5670 2250 5688 2268
rect 5670 2268 5688 2286
rect 5670 2286 5688 2304
rect 5670 2304 5688 2322
rect 5670 2322 5688 2340
rect 5670 2340 5688 2358
rect 5670 2358 5688 2376
rect 5670 2376 5688 2394
rect 5670 2394 5688 2412
rect 5670 2412 5688 2430
rect 5670 2430 5688 2448
rect 5670 2448 5688 2466
rect 5670 2466 5688 2484
rect 5670 2484 5688 2502
rect 5670 2502 5688 2520
rect 5670 2520 5688 2538
rect 5670 2538 5688 2556
rect 5670 2556 5688 2574
rect 5670 2574 5688 2592
rect 5670 2592 5688 2610
rect 5670 2808 5688 2826
rect 5670 2826 5688 2844
rect 5670 2844 5688 2862
rect 5670 2862 5688 2880
rect 5670 2880 5688 2898
rect 5670 2898 5688 2916
rect 5670 2916 5688 2934
rect 5670 2934 5688 2952
rect 5670 2952 5688 2970
rect 5670 2970 5688 2988
rect 5670 2988 5688 3006
rect 5670 3006 5688 3024
rect 5670 3024 5688 3042
rect 5670 3042 5688 3060
rect 5670 3060 5688 3078
rect 5670 3078 5688 3096
rect 5670 3096 5688 3114
rect 5670 3114 5688 3132
rect 5670 3132 5688 3150
rect 5670 3150 5688 3168
rect 5670 3168 5688 3186
rect 5670 3186 5688 3204
rect 5670 3204 5688 3222
rect 5670 3222 5688 3240
rect 5670 3240 5688 3258
rect 5670 3258 5688 3276
rect 5670 3276 5688 3294
rect 5670 3294 5688 3312
rect 5670 3312 5688 3330
rect 5670 3330 5688 3348
rect 5670 3348 5688 3366
rect 5670 3366 5688 3384
rect 5670 3384 5688 3402
rect 5670 3402 5688 3420
rect 5670 3420 5688 3438
rect 5670 3438 5688 3456
rect 5670 3456 5688 3474
rect 5670 3474 5688 3492
rect 5670 3492 5688 3510
rect 5670 3510 5688 3528
rect 5670 3528 5688 3546
rect 5670 3546 5688 3564
rect 5670 3564 5688 3582
rect 5670 3582 5688 3600
rect 5670 3600 5688 3618
rect 5670 3618 5688 3636
rect 5670 3636 5688 3654
rect 5670 3654 5688 3672
rect 5670 3672 5688 3690
rect 5670 3690 5688 3708
rect 5670 3708 5688 3726
rect 5670 3726 5688 3744
rect 5670 3744 5688 3762
rect 5670 3762 5688 3780
rect 5670 3780 5688 3798
rect 5670 3798 5688 3816
rect 5670 3816 5688 3834
rect 5670 3834 5688 3852
rect 5670 3852 5688 3870
rect 5670 3870 5688 3888
rect 5670 3888 5688 3906
rect 5670 3906 5688 3924
rect 5670 3924 5688 3942
rect 5670 3942 5688 3960
rect 5670 3960 5688 3978
rect 5670 3978 5688 3996
rect 5670 3996 5688 4014
rect 5670 4014 5688 4032
rect 5670 4032 5688 4050
rect 5670 4050 5688 4068
rect 5670 4068 5688 4086
rect 5670 4086 5688 4104
rect 5670 4104 5688 4122
rect 5670 4122 5688 4140
rect 5670 4140 5688 4158
rect 5670 4158 5688 4176
rect 5670 4176 5688 4194
rect 5670 4194 5688 4212
rect 5670 4212 5688 4230
rect 5670 4230 5688 4248
rect 5670 4248 5688 4266
rect 5670 4266 5688 4284
rect 5670 4284 5688 4302
rect 5670 4302 5688 4320
rect 5670 4320 5688 4338
rect 5670 4338 5688 4356
rect 5670 4356 5688 4374
rect 5670 4374 5688 4392
rect 5670 4392 5688 4410
rect 5670 4410 5688 4428
rect 5670 4428 5688 4446
rect 5670 4446 5688 4464
rect 5670 4464 5688 4482
rect 5670 4482 5688 4500
rect 5670 4500 5688 4518
rect 5670 4518 5688 4536
rect 5670 4536 5688 4554
rect 5670 4554 5688 4572
rect 5670 4572 5688 4590
rect 5670 4590 5688 4608
rect 5670 4608 5688 4626
rect 5670 4626 5688 4644
rect 5670 4644 5688 4662
rect 5670 4662 5688 4680
rect 5670 4680 5688 4698
rect 5670 4698 5688 4716
rect 5670 4716 5688 4734
rect 5670 4734 5688 4752
rect 5670 4752 5688 4770
rect 5670 4770 5688 4788
rect 5670 4788 5688 4806
rect 5670 4806 5688 4824
rect 5670 4824 5688 4842
rect 5670 4842 5688 4860
rect 5670 4860 5688 4878
rect 5670 4878 5688 4896
rect 5670 4896 5688 4914
rect 5670 4914 5688 4932
rect 5670 4932 5688 4950
rect 5670 4950 5688 4968
rect 5670 4968 5688 4986
rect 5670 4986 5688 5004
rect 5670 5004 5688 5022
rect 5670 5022 5688 5040
rect 5670 5040 5688 5058
rect 5670 5058 5688 5076
rect 5670 5292 5688 5310
rect 5670 5310 5688 5328
rect 5670 5328 5688 5346
rect 5670 5346 5688 5364
rect 5670 5364 5688 5382
rect 5670 5382 5688 5400
rect 5670 5400 5688 5418
rect 5670 5418 5688 5436
rect 5670 5436 5688 5454
rect 5670 5454 5688 5472
rect 5670 5472 5688 5490
rect 5670 5490 5688 5508
rect 5670 5508 5688 5526
rect 5670 5526 5688 5544
rect 5670 5544 5688 5562
rect 5670 5562 5688 5580
rect 5670 5580 5688 5598
rect 5670 5598 5688 5616
rect 5670 5616 5688 5634
rect 5670 5634 5688 5652
rect 5670 5652 5688 5670
rect 5670 5670 5688 5688
rect 5670 5688 5688 5706
rect 5670 5706 5688 5724
rect 5670 5724 5688 5742
rect 5670 5742 5688 5760
rect 5670 5760 5688 5778
rect 5670 5778 5688 5796
rect 5670 5796 5688 5814
rect 5670 5814 5688 5832
rect 5670 5832 5688 5850
rect 5670 5850 5688 5868
rect 5670 5868 5688 5886
rect 5670 5886 5688 5904
rect 5670 5904 5688 5922
rect 5670 5922 5688 5940
rect 5670 5940 5688 5958
rect 5670 5958 5688 5976
rect 5670 5976 5688 5994
rect 5670 5994 5688 6012
rect 5670 6012 5688 6030
rect 5670 6030 5688 6048
rect 5670 6048 5688 6066
rect 5670 6066 5688 6084
rect 5670 6084 5688 6102
rect 5670 6102 5688 6120
rect 5670 6120 5688 6138
rect 5670 6138 5688 6156
rect 5670 6156 5688 6174
rect 5670 6174 5688 6192
rect 5670 6192 5688 6210
rect 5670 6210 5688 6228
rect 5670 6228 5688 6246
rect 5670 6246 5688 6264
rect 5670 6264 5688 6282
rect 5670 6282 5688 6300
rect 5670 6300 5688 6318
rect 5670 6318 5688 6336
rect 5670 6336 5688 6354
rect 5670 6354 5688 6372
rect 5670 6372 5688 6390
rect 5670 6390 5688 6408
rect 5670 6408 5688 6426
rect 5670 6426 5688 6444
rect 5670 6444 5688 6462
rect 5670 6462 5688 6480
rect 5670 6480 5688 6498
rect 5670 6498 5688 6516
rect 5670 6516 5688 6534
rect 5670 6534 5688 6552
rect 5670 6552 5688 6570
rect 5670 6570 5688 6588
rect 5670 6588 5688 6606
rect 5670 6606 5688 6624
rect 5670 6624 5688 6642
rect 5670 6642 5688 6660
rect 5670 6660 5688 6678
rect 5670 6678 5688 6696
rect 5670 6696 5688 6714
rect 5670 6714 5688 6732
rect 5670 6732 5688 6750
rect 5670 6750 5688 6768
rect 5670 6768 5688 6786
rect 5670 6786 5688 6804
rect 5670 6804 5688 6822
rect 5670 6822 5688 6840
rect 5670 6840 5688 6858
rect 5670 6858 5688 6876
rect 5670 6876 5688 6894
rect 5670 6894 5688 6912
rect 5670 6912 5688 6930
rect 5670 6930 5688 6948
rect 5670 6948 5688 6966
rect 5670 6966 5688 6984
rect 5670 6984 5688 7002
rect 5670 7002 5688 7020
rect 5670 7020 5688 7038
rect 5670 7038 5688 7056
rect 5670 7056 5688 7074
rect 5670 7074 5688 7092
rect 5670 7092 5688 7110
rect 5670 7110 5688 7128
rect 5670 7128 5688 7146
rect 5670 7146 5688 7164
rect 5670 7164 5688 7182
rect 5670 7182 5688 7200
rect 5670 7200 5688 7218
rect 5670 7218 5688 7236
rect 5670 7236 5688 7254
rect 5670 7254 5688 7272
rect 5670 7272 5688 7290
rect 5670 7290 5688 7308
rect 5670 7308 5688 7326
rect 5670 7326 5688 7344
rect 5670 7344 5688 7362
rect 5670 7362 5688 7380
rect 5670 7380 5688 7398
rect 5670 7398 5688 7416
rect 5670 7416 5688 7434
rect 5670 7434 5688 7452
rect 5670 7452 5688 7470
rect 5670 7470 5688 7488
rect 5670 7488 5688 7506
rect 5670 7506 5688 7524
rect 5670 7524 5688 7542
rect 5670 7542 5688 7560
rect 5670 7560 5688 7578
rect 5670 7578 5688 7596
rect 5670 7596 5688 7614
rect 5670 7614 5688 7632
rect 5670 7632 5688 7650
rect 5670 7650 5688 7668
rect 5670 7668 5688 7686
rect 5670 7686 5688 7704
rect 5670 7704 5688 7722
rect 5670 7722 5688 7740
rect 5670 7740 5688 7758
rect 5670 7758 5688 7776
rect 5670 7776 5688 7794
rect 5670 7794 5688 7812
rect 5670 7812 5688 7830
rect 5670 7830 5688 7848
rect 5670 7848 5688 7866
rect 5670 7866 5688 7884
rect 5670 7884 5688 7902
rect 5670 7902 5688 7920
rect 5670 7920 5688 7938
rect 5670 7938 5688 7956
rect 5670 7956 5688 7974
rect 5670 7974 5688 7992
rect 5670 7992 5688 8010
rect 5670 8010 5688 8028
rect 5670 8028 5688 8046
rect 5670 8046 5688 8064
rect 5670 8064 5688 8082
rect 5670 8082 5688 8100
rect 5670 8100 5688 8118
rect 5670 8118 5688 8136
rect 5670 8136 5688 8154
rect 5670 8154 5688 8172
rect 5670 8172 5688 8190
rect 5670 8190 5688 8208
rect 5670 8208 5688 8226
rect 5670 8226 5688 8244
rect 5670 8244 5688 8262
rect 5670 8262 5688 8280
rect 5670 8280 5688 8298
rect 5670 8298 5688 8316
rect 5670 8316 5688 8334
rect 5670 8334 5688 8352
rect 5670 8352 5688 8370
rect 5670 8370 5688 8388
rect 5670 8388 5688 8406
rect 5670 8406 5688 8424
rect 5670 8424 5688 8442
rect 5670 8442 5688 8460
rect 5670 8460 5688 8478
rect 5670 8478 5688 8496
rect 5670 8496 5688 8514
rect 5670 8514 5688 8532
rect 5670 8532 5688 8550
rect 5670 8550 5688 8568
rect 5670 8568 5688 8586
rect 5670 8586 5688 8604
rect 5670 8604 5688 8622
rect 5670 8622 5688 8640
rect 5670 8640 5688 8658
rect 5670 8658 5688 8676
rect 5670 8676 5688 8694
rect 5670 8694 5688 8712
rect 5670 8712 5688 8730
rect 5670 8730 5688 8748
rect 5670 8748 5688 8766
rect 5670 8766 5688 8784
rect 5670 8784 5688 8802
rect 5688 648 5706 666
rect 5688 666 5706 684
rect 5688 684 5706 702
rect 5688 702 5706 720
rect 5688 720 5706 738
rect 5688 738 5706 756
rect 5688 756 5706 774
rect 5688 774 5706 792
rect 5688 792 5706 810
rect 5688 810 5706 828
rect 5688 828 5706 846
rect 5688 846 5706 864
rect 5688 864 5706 882
rect 5688 882 5706 900
rect 5688 900 5706 918
rect 5688 918 5706 936
rect 5688 936 5706 954
rect 5688 954 5706 972
rect 5688 972 5706 990
rect 5688 1134 5706 1152
rect 5688 1152 5706 1170
rect 5688 1170 5706 1188
rect 5688 1188 5706 1206
rect 5688 1206 5706 1224
rect 5688 1224 5706 1242
rect 5688 1242 5706 1260
rect 5688 1260 5706 1278
rect 5688 1278 5706 1296
rect 5688 1296 5706 1314
rect 5688 1314 5706 1332
rect 5688 1332 5706 1350
rect 5688 1350 5706 1368
rect 5688 1368 5706 1386
rect 5688 1386 5706 1404
rect 5688 1404 5706 1422
rect 5688 1422 5706 1440
rect 5688 1440 5706 1458
rect 5688 1458 5706 1476
rect 5688 1476 5706 1494
rect 5688 1494 5706 1512
rect 5688 1512 5706 1530
rect 5688 1530 5706 1548
rect 5688 1548 5706 1566
rect 5688 1566 5706 1584
rect 5688 1584 5706 1602
rect 5688 1602 5706 1620
rect 5688 1620 5706 1638
rect 5688 1638 5706 1656
rect 5688 1656 5706 1674
rect 5688 1674 5706 1692
rect 5688 1692 5706 1710
rect 5688 1710 5706 1728
rect 5688 1728 5706 1746
rect 5688 1746 5706 1764
rect 5688 1764 5706 1782
rect 5688 1782 5706 1800
rect 5688 1800 5706 1818
rect 5688 1818 5706 1836
rect 5688 1836 5706 1854
rect 5688 1854 5706 1872
rect 5688 1872 5706 1890
rect 5688 1890 5706 1908
rect 5688 1908 5706 1926
rect 5688 1926 5706 1944
rect 5688 1944 5706 1962
rect 5688 1962 5706 1980
rect 5688 1980 5706 1998
rect 5688 1998 5706 2016
rect 5688 2016 5706 2034
rect 5688 2034 5706 2052
rect 5688 2052 5706 2070
rect 5688 2070 5706 2088
rect 5688 2088 5706 2106
rect 5688 2106 5706 2124
rect 5688 2124 5706 2142
rect 5688 2142 5706 2160
rect 5688 2160 5706 2178
rect 5688 2178 5706 2196
rect 5688 2196 5706 2214
rect 5688 2214 5706 2232
rect 5688 2232 5706 2250
rect 5688 2250 5706 2268
rect 5688 2268 5706 2286
rect 5688 2286 5706 2304
rect 5688 2304 5706 2322
rect 5688 2322 5706 2340
rect 5688 2340 5706 2358
rect 5688 2358 5706 2376
rect 5688 2376 5706 2394
rect 5688 2394 5706 2412
rect 5688 2412 5706 2430
rect 5688 2430 5706 2448
rect 5688 2448 5706 2466
rect 5688 2466 5706 2484
rect 5688 2484 5706 2502
rect 5688 2502 5706 2520
rect 5688 2520 5706 2538
rect 5688 2538 5706 2556
rect 5688 2556 5706 2574
rect 5688 2574 5706 2592
rect 5688 2592 5706 2610
rect 5688 2826 5706 2844
rect 5688 2844 5706 2862
rect 5688 2862 5706 2880
rect 5688 2880 5706 2898
rect 5688 2898 5706 2916
rect 5688 2916 5706 2934
rect 5688 2934 5706 2952
rect 5688 2952 5706 2970
rect 5688 2970 5706 2988
rect 5688 2988 5706 3006
rect 5688 3006 5706 3024
rect 5688 3024 5706 3042
rect 5688 3042 5706 3060
rect 5688 3060 5706 3078
rect 5688 3078 5706 3096
rect 5688 3096 5706 3114
rect 5688 3114 5706 3132
rect 5688 3132 5706 3150
rect 5688 3150 5706 3168
rect 5688 3168 5706 3186
rect 5688 3186 5706 3204
rect 5688 3204 5706 3222
rect 5688 3222 5706 3240
rect 5688 3240 5706 3258
rect 5688 3258 5706 3276
rect 5688 3276 5706 3294
rect 5688 3294 5706 3312
rect 5688 3312 5706 3330
rect 5688 3330 5706 3348
rect 5688 3348 5706 3366
rect 5688 3366 5706 3384
rect 5688 3384 5706 3402
rect 5688 3402 5706 3420
rect 5688 3420 5706 3438
rect 5688 3438 5706 3456
rect 5688 3456 5706 3474
rect 5688 3474 5706 3492
rect 5688 3492 5706 3510
rect 5688 3510 5706 3528
rect 5688 3528 5706 3546
rect 5688 3546 5706 3564
rect 5688 3564 5706 3582
rect 5688 3582 5706 3600
rect 5688 3600 5706 3618
rect 5688 3618 5706 3636
rect 5688 3636 5706 3654
rect 5688 3654 5706 3672
rect 5688 3672 5706 3690
rect 5688 3690 5706 3708
rect 5688 3708 5706 3726
rect 5688 3726 5706 3744
rect 5688 3744 5706 3762
rect 5688 3762 5706 3780
rect 5688 3780 5706 3798
rect 5688 3798 5706 3816
rect 5688 3816 5706 3834
rect 5688 3834 5706 3852
rect 5688 3852 5706 3870
rect 5688 3870 5706 3888
rect 5688 3888 5706 3906
rect 5688 3906 5706 3924
rect 5688 3924 5706 3942
rect 5688 3942 5706 3960
rect 5688 3960 5706 3978
rect 5688 3978 5706 3996
rect 5688 3996 5706 4014
rect 5688 4014 5706 4032
rect 5688 4032 5706 4050
rect 5688 4050 5706 4068
rect 5688 4068 5706 4086
rect 5688 4086 5706 4104
rect 5688 4104 5706 4122
rect 5688 4122 5706 4140
rect 5688 4140 5706 4158
rect 5688 4158 5706 4176
rect 5688 4176 5706 4194
rect 5688 4194 5706 4212
rect 5688 4212 5706 4230
rect 5688 4230 5706 4248
rect 5688 4248 5706 4266
rect 5688 4266 5706 4284
rect 5688 4284 5706 4302
rect 5688 4302 5706 4320
rect 5688 4320 5706 4338
rect 5688 4338 5706 4356
rect 5688 4356 5706 4374
rect 5688 4374 5706 4392
rect 5688 4392 5706 4410
rect 5688 4410 5706 4428
rect 5688 4428 5706 4446
rect 5688 4446 5706 4464
rect 5688 4464 5706 4482
rect 5688 4482 5706 4500
rect 5688 4500 5706 4518
rect 5688 4518 5706 4536
rect 5688 4536 5706 4554
rect 5688 4554 5706 4572
rect 5688 4572 5706 4590
rect 5688 4590 5706 4608
rect 5688 4608 5706 4626
rect 5688 4626 5706 4644
rect 5688 4644 5706 4662
rect 5688 4662 5706 4680
rect 5688 4680 5706 4698
rect 5688 4698 5706 4716
rect 5688 4716 5706 4734
rect 5688 4734 5706 4752
rect 5688 4752 5706 4770
rect 5688 4770 5706 4788
rect 5688 4788 5706 4806
rect 5688 4806 5706 4824
rect 5688 4824 5706 4842
rect 5688 4842 5706 4860
rect 5688 4860 5706 4878
rect 5688 4878 5706 4896
rect 5688 4896 5706 4914
rect 5688 4914 5706 4932
rect 5688 4932 5706 4950
rect 5688 4950 5706 4968
rect 5688 4968 5706 4986
rect 5688 4986 5706 5004
rect 5688 5004 5706 5022
rect 5688 5022 5706 5040
rect 5688 5040 5706 5058
rect 5688 5058 5706 5076
rect 5688 5076 5706 5094
rect 5688 5310 5706 5328
rect 5688 5328 5706 5346
rect 5688 5346 5706 5364
rect 5688 5364 5706 5382
rect 5688 5382 5706 5400
rect 5688 5400 5706 5418
rect 5688 5418 5706 5436
rect 5688 5436 5706 5454
rect 5688 5454 5706 5472
rect 5688 5472 5706 5490
rect 5688 5490 5706 5508
rect 5688 5508 5706 5526
rect 5688 5526 5706 5544
rect 5688 5544 5706 5562
rect 5688 5562 5706 5580
rect 5688 5580 5706 5598
rect 5688 5598 5706 5616
rect 5688 5616 5706 5634
rect 5688 5634 5706 5652
rect 5688 5652 5706 5670
rect 5688 5670 5706 5688
rect 5688 5688 5706 5706
rect 5688 5706 5706 5724
rect 5688 5724 5706 5742
rect 5688 5742 5706 5760
rect 5688 5760 5706 5778
rect 5688 5778 5706 5796
rect 5688 5796 5706 5814
rect 5688 5814 5706 5832
rect 5688 5832 5706 5850
rect 5688 5850 5706 5868
rect 5688 5868 5706 5886
rect 5688 5886 5706 5904
rect 5688 5904 5706 5922
rect 5688 5922 5706 5940
rect 5688 5940 5706 5958
rect 5688 5958 5706 5976
rect 5688 5976 5706 5994
rect 5688 5994 5706 6012
rect 5688 6012 5706 6030
rect 5688 6030 5706 6048
rect 5688 6048 5706 6066
rect 5688 6066 5706 6084
rect 5688 6084 5706 6102
rect 5688 6102 5706 6120
rect 5688 6120 5706 6138
rect 5688 6138 5706 6156
rect 5688 6156 5706 6174
rect 5688 6174 5706 6192
rect 5688 6192 5706 6210
rect 5688 6210 5706 6228
rect 5688 6228 5706 6246
rect 5688 6246 5706 6264
rect 5688 6264 5706 6282
rect 5688 6282 5706 6300
rect 5688 6300 5706 6318
rect 5688 6318 5706 6336
rect 5688 6336 5706 6354
rect 5688 6354 5706 6372
rect 5688 6372 5706 6390
rect 5688 6390 5706 6408
rect 5688 6408 5706 6426
rect 5688 6426 5706 6444
rect 5688 6444 5706 6462
rect 5688 6462 5706 6480
rect 5688 6480 5706 6498
rect 5688 6498 5706 6516
rect 5688 6516 5706 6534
rect 5688 6534 5706 6552
rect 5688 6552 5706 6570
rect 5688 6570 5706 6588
rect 5688 6588 5706 6606
rect 5688 6606 5706 6624
rect 5688 6624 5706 6642
rect 5688 6642 5706 6660
rect 5688 6660 5706 6678
rect 5688 6678 5706 6696
rect 5688 6696 5706 6714
rect 5688 6714 5706 6732
rect 5688 6732 5706 6750
rect 5688 6750 5706 6768
rect 5688 6768 5706 6786
rect 5688 6786 5706 6804
rect 5688 6804 5706 6822
rect 5688 6822 5706 6840
rect 5688 6840 5706 6858
rect 5688 6858 5706 6876
rect 5688 6876 5706 6894
rect 5688 6894 5706 6912
rect 5688 6912 5706 6930
rect 5688 6930 5706 6948
rect 5688 6948 5706 6966
rect 5688 6966 5706 6984
rect 5688 6984 5706 7002
rect 5688 7002 5706 7020
rect 5688 7020 5706 7038
rect 5688 7038 5706 7056
rect 5688 7056 5706 7074
rect 5688 7074 5706 7092
rect 5688 7092 5706 7110
rect 5688 7110 5706 7128
rect 5688 7128 5706 7146
rect 5688 7146 5706 7164
rect 5688 7164 5706 7182
rect 5688 7182 5706 7200
rect 5688 7200 5706 7218
rect 5688 7218 5706 7236
rect 5688 7236 5706 7254
rect 5688 7254 5706 7272
rect 5688 7272 5706 7290
rect 5688 7290 5706 7308
rect 5688 7308 5706 7326
rect 5688 7326 5706 7344
rect 5688 7344 5706 7362
rect 5688 7362 5706 7380
rect 5688 7380 5706 7398
rect 5688 7398 5706 7416
rect 5688 7416 5706 7434
rect 5688 7434 5706 7452
rect 5688 7452 5706 7470
rect 5688 7470 5706 7488
rect 5688 7488 5706 7506
rect 5688 7506 5706 7524
rect 5688 7524 5706 7542
rect 5688 7542 5706 7560
rect 5688 7560 5706 7578
rect 5688 7578 5706 7596
rect 5688 7596 5706 7614
rect 5688 7614 5706 7632
rect 5688 7632 5706 7650
rect 5688 7650 5706 7668
rect 5688 7668 5706 7686
rect 5688 7686 5706 7704
rect 5688 7704 5706 7722
rect 5688 7722 5706 7740
rect 5688 7740 5706 7758
rect 5688 7758 5706 7776
rect 5688 7776 5706 7794
rect 5688 7794 5706 7812
rect 5688 7812 5706 7830
rect 5688 7830 5706 7848
rect 5688 7848 5706 7866
rect 5688 7866 5706 7884
rect 5688 7884 5706 7902
rect 5688 7902 5706 7920
rect 5688 7920 5706 7938
rect 5688 7938 5706 7956
rect 5688 7956 5706 7974
rect 5688 7974 5706 7992
rect 5688 7992 5706 8010
rect 5688 8010 5706 8028
rect 5688 8028 5706 8046
rect 5688 8046 5706 8064
rect 5688 8064 5706 8082
rect 5688 8082 5706 8100
rect 5688 8100 5706 8118
rect 5688 8118 5706 8136
rect 5688 8136 5706 8154
rect 5688 8154 5706 8172
rect 5688 8172 5706 8190
rect 5688 8190 5706 8208
rect 5688 8208 5706 8226
rect 5688 8226 5706 8244
rect 5688 8244 5706 8262
rect 5688 8262 5706 8280
rect 5688 8280 5706 8298
rect 5688 8298 5706 8316
rect 5688 8316 5706 8334
rect 5688 8334 5706 8352
rect 5688 8352 5706 8370
rect 5688 8370 5706 8388
rect 5688 8388 5706 8406
rect 5688 8406 5706 8424
rect 5688 8424 5706 8442
rect 5688 8442 5706 8460
rect 5688 8460 5706 8478
rect 5688 8478 5706 8496
rect 5688 8496 5706 8514
rect 5688 8514 5706 8532
rect 5688 8532 5706 8550
rect 5688 8550 5706 8568
rect 5688 8568 5706 8586
rect 5688 8586 5706 8604
rect 5688 8604 5706 8622
rect 5688 8622 5706 8640
rect 5688 8640 5706 8658
rect 5688 8658 5706 8676
rect 5688 8676 5706 8694
rect 5688 8694 5706 8712
rect 5688 8712 5706 8730
rect 5688 8730 5706 8748
rect 5688 8748 5706 8766
rect 5688 8766 5706 8784
rect 5688 8784 5706 8802
rect 5688 8802 5706 8820
rect 5706 666 5724 684
rect 5706 684 5724 702
rect 5706 702 5724 720
rect 5706 720 5724 738
rect 5706 738 5724 756
rect 5706 756 5724 774
rect 5706 774 5724 792
rect 5706 792 5724 810
rect 5706 810 5724 828
rect 5706 828 5724 846
rect 5706 846 5724 864
rect 5706 864 5724 882
rect 5706 882 5724 900
rect 5706 900 5724 918
rect 5706 918 5724 936
rect 5706 936 5724 954
rect 5706 954 5724 972
rect 5706 972 5724 990
rect 5706 1134 5724 1152
rect 5706 1152 5724 1170
rect 5706 1170 5724 1188
rect 5706 1188 5724 1206
rect 5706 1206 5724 1224
rect 5706 1224 5724 1242
rect 5706 1242 5724 1260
rect 5706 1260 5724 1278
rect 5706 1278 5724 1296
rect 5706 1296 5724 1314
rect 5706 1314 5724 1332
rect 5706 1332 5724 1350
rect 5706 1350 5724 1368
rect 5706 1368 5724 1386
rect 5706 1386 5724 1404
rect 5706 1404 5724 1422
rect 5706 1422 5724 1440
rect 5706 1440 5724 1458
rect 5706 1458 5724 1476
rect 5706 1476 5724 1494
rect 5706 1494 5724 1512
rect 5706 1512 5724 1530
rect 5706 1530 5724 1548
rect 5706 1548 5724 1566
rect 5706 1566 5724 1584
rect 5706 1584 5724 1602
rect 5706 1602 5724 1620
rect 5706 1620 5724 1638
rect 5706 1638 5724 1656
rect 5706 1656 5724 1674
rect 5706 1674 5724 1692
rect 5706 1692 5724 1710
rect 5706 1710 5724 1728
rect 5706 1728 5724 1746
rect 5706 1746 5724 1764
rect 5706 1764 5724 1782
rect 5706 1782 5724 1800
rect 5706 1800 5724 1818
rect 5706 1818 5724 1836
rect 5706 1836 5724 1854
rect 5706 1854 5724 1872
rect 5706 1872 5724 1890
rect 5706 1890 5724 1908
rect 5706 1908 5724 1926
rect 5706 1926 5724 1944
rect 5706 1944 5724 1962
rect 5706 1962 5724 1980
rect 5706 1980 5724 1998
rect 5706 1998 5724 2016
rect 5706 2016 5724 2034
rect 5706 2034 5724 2052
rect 5706 2052 5724 2070
rect 5706 2070 5724 2088
rect 5706 2088 5724 2106
rect 5706 2106 5724 2124
rect 5706 2124 5724 2142
rect 5706 2142 5724 2160
rect 5706 2160 5724 2178
rect 5706 2178 5724 2196
rect 5706 2196 5724 2214
rect 5706 2214 5724 2232
rect 5706 2232 5724 2250
rect 5706 2250 5724 2268
rect 5706 2268 5724 2286
rect 5706 2286 5724 2304
rect 5706 2304 5724 2322
rect 5706 2322 5724 2340
rect 5706 2340 5724 2358
rect 5706 2358 5724 2376
rect 5706 2376 5724 2394
rect 5706 2394 5724 2412
rect 5706 2412 5724 2430
rect 5706 2430 5724 2448
rect 5706 2448 5724 2466
rect 5706 2466 5724 2484
rect 5706 2484 5724 2502
rect 5706 2502 5724 2520
rect 5706 2520 5724 2538
rect 5706 2538 5724 2556
rect 5706 2556 5724 2574
rect 5706 2574 5724 2592
rect 5706 2592 5724 2610
rect 5706 2610 5724 2628
rect 5706 2826 5724 2844
rect 5706 2844 5724 2862
rect 5706 2862 5724 2880
rect 5706 2880 5724 2898
rect 5706 2898 5724 2916
rect 5706 2916 5724 2934
rect 5706 2934 5724 2952
rect 5706 2952 5724 2970
rect 5706 2970 5724 2988
rect 5706 2988 5724 3006
rect 5706 3006 5724 3024
rect 5706 3024 5724 3042
rect 5706 3042 5724 3060
rect 5706 3060 5724 3078
rect 5706 3078 5724 3096
rect 5706 3096 5724 3114
rect 5706 3114 5724 3132
rect 5706 3132 5724 3150
rect 5706 3150 5724 3168
rect 5706 3168 5724 3186
rect 5706 3186 5724 3204
rect 5706 3204 5724 3222
rect 5706 3222 5724 3240
rect 5706 3240 5724 3258
rect 5706 3258 5724 3276
rect 5706 3276 5724 3294
rect 5706 3294 5724 3312
rect 5706 3312 5724 3330
rect 5706 3330 5724 3348
rect 5706 3348 5724 3366
rect 5706 3366 5724 3384
rect 5706 3384 5724 3402
rect 5706 3402 5724 3420
rect 5706 3420 5724 3438
rect 5706 3438 5724 3456
rect 5706 3456 5724 3474
rect 5706 3474 5724 3492
rect 5706 3492 5724 3510
rect 5706 3510 5724 3528
rect 5706 3528 5724 3546
rect 5706 3546 5724 3564
rect 5706 3564 5724 3582
rect 5706 3582 5724 3600
rect 5706 3600 5724 3618
rect 5706 3618 5724 3636
rect 5706 3636 5724 3654
rect 5706 3654 5724 3672
rect 5706 3672 5724 3690
rect 5706 3690 5724 3708
rect 5706 3708 5724 3726
rect 5706 3726 5724 3744
rect 5706 3744 5724 3762
rect 5706 3762 5724 3780
rect 5706 3780 5724 3798
rect 5706 3798 5724 3816
rect 5706 3816 5724 3834
rect 5706 3834 5724 3852
rect 5706 3852 5724 3870
rect 5706 3870 5724 3888
rect 5706 3888 5724 3906
rect 5706 3906 5724 3924
rect 5706 3924 5724 3942
rect 5706 3942 5724 3960
rect 5706 3960 5724 3978
rect 5706 3978 5724 3996
rect 5706 3996 5724 4014
rect 5706 4014 5724 4032
rect 5706 4032 5724 4050
rect 5706 4050 5724 4068
rect 5706 4068 5724 4086
rect 5706 4086 5724 4104
rect 5706 4104 5724 4122
rect 5706 4122 5724 4140
rect 5706 4140 5724 4158
rect 5706 4158 5724 4176
rect 5706 4176 5724 4194
rect 5706 4194 5724 4212
rect 5706 4212 5724 4230
rect 5706 4230 5724 4248
rect 5706 4248 5724 4266
rect 5706 4266 5724 4284
rect 5706 4284 5724 4302
rect 5706 4302 5724 4320
rect 5706 4320 5724 4338
rect 5706 4338 5724 4356
rect 5706 4356 5724 4374
rect 5706 4374 5724 4392
rect 5706 4392 5724 4410
rect 5706 4410 5724 4428
rect 5706 4428 5724 4446
rect 5706 4446 5724 4464
rect 5706 4464 5724 4482
rect 5706 4482 5724 4500
rect 5706 4500 5724 4518
rect 5706 4518 5724 4536
rect 5706 4536 5724 4554
rect 5706 4554 5724 4572
rect 5706 4572 5724 4590
rect 5706 4590 5724 4608
rect 5706 4608 5724 4626
rect 5706 4626 5724 4644
rect 5706 4644 5724 4662
rect 5706 4662 5724 4680
rect 5706 4680 5724 4698
rect 5706 4698 5724 4716
rect 5706 4716 5724 4734
rect 5706 4734 5724 4752
rect 5706 4752 5724 4770
rect 5706 4770 5724 4788
rect 5706 4788 5724 4806
rect 5706 4806 5724 4824
rect 5706 4824 5724 4842
rect 5706 4842 5724 4860
rect 5706 4860 5724 4878
rect 5706 4878 5724 4896
rect 5706 4896 5724 4914
rect 5706 4914 5724 4932
rect 5706 4932 5724 4950
rect 5706 4950 5724 4968
rect 5706 4968 5724 4986
rect 5706 4986 5724 5004
rect 5706 5004 5724 5022
rect 5706 5022 5724 5040
rect 5706 5040 5724 5058
rect 5706 5058 5724 5076
rect 5706 5076 5724 5094
rect 5706 5094 5724 5112
rect 5706 5328 5724 5346
rect 5706 5346 5724 5364
rect 5706 5364 5724 5382
rect 5706 5382 5724 5400
rect 5706 5400 5724 5418
rect 5706 5418 5724 5436
rect 5706 5436 5724 5454
rect 5706 5454 5724 5472
rect 5706 5472 5724 5490
rect 5706 5490 5724 5508
rect 5706 5508 5724 5526
rect 5706 5526 5724 5544
rect 5706 5544 5724 5562
rect 5706 5562 5724 5580
rect 5706 5580 5724 5598
rect 5706 5598 5724 5616
rect 5706 5616 5724 5634
rect 5706 5634 5724 5652
rect 5706 5652 5724 5670
rect 5706 5670 5724 5688
rect 5706 5688 5724 5706
rect 5706 5706 5724 5724
rect 5706 5724 5724 5742
rect 5706 5742 5724 5760
rect 5706 5760 5724 5778
rect 5706 5778 5724 5796
rect 5706 5796 5724 5814
rect 5706 5814 5724 5832
rect 5706 5832 5724 5850
rect 5706 5850 5724 5868
rect 5706 5868 5724 5886
rect 5706 5886 5724 5904
rect 5706 5904 5724 5922
rect 5706 5922 5724 5940
rect 5706 5940 5724 5958
rect 5706 5958 5724 5976
rect 5706 5976 5724 5994
rect 5706 5994 5724 6012
rect 5706 6012 5724 6030
rect 5706 6030 5724 6048
rect 5706 6048 5724 6066
rect 5706 6066 5724 6084
rect 5706 6084 5724 6102
rect 5706 6102 5724 6120
rect 5706 6120 5724 6138
rect 5706 6138 5724 6156
rect 5706 6156 5724 6174
rect 5706 6174 5724 6192
rect 5706 6192 5724 6210
rect 5706 6210 5724 6228
rect 5706 6228 5724 6246
rect 5706 6246 5724 6264
rect 5706 6264 5724 6282
rect 5706 6282 5724 6300
rect 5706 6300 5724 6318
rect 5706 6318 5724 6336
rect 5706 6336 5724 6354
rect 5706 6354 5724 6372
rect 5706 6372 5724 6390
rect 5706 6390 5724 6408
rect 5706 6408 5724 6426
rect 5706 6426 5724 6444
rect 5706 6444 5724 6462
rect 5706 6462 5724 6480
rect 5706 6480 5724 6498
rect 5706 6498 5724 6516
rect 5706 6516 5724 6534
rect 5706 6534 5724 6552
rect 5706 6552 5724 6570
rect 5706 6570 5724 6588
rect 5706 6588 5724 6606
rect 5706 6606 5724 6624
rect 5706 6624 5724 6642
rect 5706 6642 5724 6660
rect 5706 6660 5724 6678
rect 5706 6678 5724 6696
rect 5706 6696 5724 6714
rect 5706 6714 5724 6732
rect 5706 6732 5724 6750
rect 5706 6750 5724 6768
rect 5706 6768 5724 6786
rect 5706 6786 5724 6804
rect 5706 6804 5724 6822
rect 5706 6822 5724 6840
rect 5706 6840 5724 6858
rect 5706 6858 5724 6876
rect 5706 6876 5724 6894
rect 5706 6894 5724 6912
rect 5706 6912 5724 6930
rect 5706 6930 5724 6948
rect 5706 6948 5724 6966
rect 5706 6966 5724 6984
rect 5706 6984 5724 7002
rect 5706 7002 5724 7020
rect 5706 7020 5724 7038
rect 5706 7038 5724 7056
rect 5706 7056 5724 7074
rect 5706 7074 5724 7092
rect 5706 7092 5724 7110
rect 5706 7110 5724 7128
rect 5706 7128 5724 7146
rect 5706 7146 5724 7164
rect 5706 7164 5724 7182
rect 5706 7182 5724 7200
rect 5706 7200 5724 7218
rect 5706 7218 5724 7236
rect 5706 7236 5724 7254
rect 5706 7254 5724 7272
rect 5706 7272 5724 7290
rect 5706 7290 5724 7308
rect 5706 7308 5724 7326
rect 5706 7326 5724 7344
rect 5706 7344 5724 7362
rect 5706 7362 5724 7380
rect 5706 7380 5724 7398
rect 5706 7398 5724 7416
rect 5706 7416 5724 7434
rect 5706 7434 5724 7452
rect 5706 7452 5724 7470
rect 5706 7470 5724 7488
rect 5706 7488 5724 7506
rect 5706 7506 5724 7524
rect 5706 7524 5724 7542
rect 5706 7542 5724 7560
rect 5706 7560 5724 7578
rect 5706 7578 5724 7596
rect 5706 7596 5724 7614
rect 5706 7614 5724 7632
rect 5706 7632 5724 7650
rect 5706 7650 5724 7668
rect 5706 7668 5724 7686
rect 5706 7686 5724 7704
rect 5706 7704 5724 7722
rect 5706 7722 5724 7740
rect 5706 7740 5724 7758
rect 5706 7758 5724 7776
rect 5706 7776 5724 7794
rect 5706 7794 5724 7812
rect 5706 7812 5724 7830
rect 5706 7830 5724 7848
rect 5706 7848 5724 7866
rect 5706 7866 5724 7884
rect 5706 7884 5724 7902
rect 5706 7902 5724 7920
rect 5706 7920 5724 7938
rect 5706 7938 5724 7956
rect 5706 7956 5724 7974
rect 5706 7974 5724 7992
rect 5706 7992 5724 8010
rect 5706 8010 5724 8028
rect 5706 8028 5724 8046
rect 5706 8046 5724 8064
rect 5706 8064 5724 8082
rect 5706 8082 5724 8100
rect 5706 8100 5724 8118
rect 5706 8118 5724 8136
rect 5706 8136 5724 8154
rect 5706 8154 5724 8172
rect 5706 8172 5724 8190
rect 5706 8190 5724 8208
rect 5706 8208 5724 8226
rect 5706 8226 5724 8244
rect 5706 8244 5724 8262
rect 5706 8262 5724 8280
rect 5706 8280 5724 8298
rect 5706 8298 5724 8316
rect 5706 8316 5724 8334
rect 5706 8334 5724 8352
rect 5706 8352 5724 8370
rect 5706 8370 5724 8388
rect 5706 8388 5724 8406
rect 5706 8406 5724 8424
rect 5706 8424 5724 8442
rect 5706 8442 5724 8460
rect 5706 8460 5724 8478
rect 5706 8478 5724 8496
rect 5706 8496 5724 8514
rect 5706 8514 5724 8532
rect 5706 8532 5724 8550
rect 5706 8550 5724 8568
rect 5706 8568 5724 8586
rect 5706 8586 5724 8604
rect 5706 8604 5724 8622
rect 5706 8622 5724 8640
rect 5706 8640 5724 8658
rect 5706 8658 5724 8676
rect 5706 8676 5724 8694
rect 5706 8694 5724 8712
rect 5706 8712 5724 8730
rect 5706 8730 5724 8748
rect 5706 8748 5724 8766
rect 5706 8766 5724 8784
rect 5706 8784 5724 8802
rect 5706 8802 5724 8820
rect 5706 8820 5724 8838
rect 5724 684 5742 702
rect 5724 702 5742 720
rect 5724 720 5742 738
rect 5724 738 5742 756
rect 5724 756 5742 774
rect 5724 774 5742 792
rect 5724 792 5742 810
rect 5724 810 5742 828
rect 5724 828 5742 846
rect 5724 846 5742 864
rect 5724 864 5742 882
rect 5724 882 5742 900
rect 5724 900 5742 918
rect 5724 918 5742 936
rect 5724 936 5742 954
rect 5724 954 5742 972
rect 5724 972 5742 990
rect 5724 990 5742 1008
rect 5724 1152 5742 1170
rect 5724 1170 5742 1188
rect 5724 1188 5742 1206
rect 5724 1206 5742 1224
rect 5724 1224 5742 1242
rect 5724 1242 5742 1260
rect 5724 1260 5742 1278
rect 5724 1278 5742 1296
rect 5724 1296 5742 1314
rect 5724 1314 5742 1332
rect 5724 1332 5742 1350
rect 5724 1350 5742 1368
rect 5724 1368 5742 1386
rect 5724 1386 5742 1404
rect 5724 1404 5742 1422
rect 5724 1422 5742 1440
rect 5724 1440 5742 1458
rect 5724 1458 5742 1476
rect 5724 1476 5742 1494
rect 5724 1494 5742 1512
rect 5724 1512 5742 1530
rect 5724 1530 5742 1548
rect 5724 1548 5742 1566
rect 5724 1566 5742 1584
rect 5724 1584 5742 1602
rect 5724 1602 5742 1620
rect 5724 1620 5742 1638
rect 5724 1638 5742 1656
rect 5724 1656 5742 1674
rect 5724 1674 5742 1692
rect 5724 1692 5742 1710
rect 5724 1710 5742 1728
rect 5724 1728 5742 1746
rect 5724 1746 5742 1764
rect 5724 1764 5742 1782
rect 5724 1782 5742 1800
rect 5724 1800 5742 1818
rect 5724 1818 5742 1836
rect 5724 1836 5742 1854
rect 5724 1854 5742 1872
rect 5724 1872 5742 1890
rect 5724 1890 5742 1908
rect 5724 1908 5742 1926
rect 5724 1926 5742 1944
rect 5724 1944 5742 1962
rect 5724 1962 5742 1980
rect 5724 1980 5742 1998
rect 5724 1998 5742 2016
rect 5724 2016 5742 2034
rect 5724 2034 5742 2052
rect 5724 2052 5742 2070
rect 5724 2070 5742 2088
rect 5724 2088 5742 2106
rect 5724 2106 5742 2124
rect 5724 2124 5742 2142
rect 5724 2142 5742 2160
rect 5724 2160 5742 2178
rect 5724 2178 5742 2196
rect 5724 2196 5742 2214
rect 5724 2214 5742 2232
rect 5724 2232 5742 2250
rect 5724 2250 5742 2268
rect 5724 2268 5742 2286
rect 5724 2286 5742 2304
rect 5724 2304 5742 2322
rect 5724 2322 5742 2340
rect 5724 2340 5742 2358
rect 5724 2358 5742 2376
rect 5724 2376 5742 2394
rect 5724 2394 5742 2412
rect 5724 2412 5742 2430
rect 5724 2430 5742 2448
rect 5724 2448 5742 2466
rect 5724 2466 5742 2484
rect 5724 2484 5742 2502
rect 5724 2502 5742 2520
rect 5724 2520 5742 2538
rect 5724 2538 5742 2556
rect 5724 2556 5742 2574
rect 5724 2574 5742 2592
rect 5724 2592 5742 2610
rect 5724 2610 5742 2628
rect 5724 2844 5742 2862
rect 5724 2862 5742 2880
rect 5724 2880 5742 2898
rect 5724 2898 5742 2916
rect 5724 2916 5742 2934
rect 5724 2934 5742 2952
rect 5724 2952 5742 2970
rect 5724 2970 5742 2988
rect 5724 2988 5742 3006
rect 5724 3006 5742 3024
rect 5724 3024 5742 3042
rect 5724 3042 5742 3060
rect 5724 3060 5742 3078
rect 5724 3078 5742 3096
rect 5724 3096 5742 3114
rect 5724 3114 5742 3132
rect 5724 3132 5742 3150
rect 5724 3150 5742 3168
rect 5724 3168 5742 3186
rect 5724 3186 5742 3204
rect 5724 3204 5742 3222
rect 5724 3222 5742 3240
rect 5724 3240 5742 3258
rect 5724 3258 5742 3276
rect 5724 3276 5742 3294
rect 5724 3294 5742 3312
rect 5724 3312 5742 3330
rect 5724 3330 5742 3348
rect 5724 3348 5742 3366
rect 5724 3366 5742 3384
rect 5724 3384 5742 3402
rect 5724 3402 5742 3420
rect 5724 3420 5742 3438
rect 5724 3438 5742 3456
rect 5724 3456 5742 3474
rect 5724 3474 5742 3492
rect 5724 3492 5742 3510
rect 5724 3510 5742 3528
rect 5724 3528 5742 3546
rect 5724 3546 5742 3564
rect 5724 3564 5742 3582
rect 5724 3582 5742 3600
rect 5724 3600 5742 3618
rect 5724 3618 5742 3636
rect 5724 3636 5742 3654
rect 5724 3654 5742 3672
rect 5724 3672 5742 3690
rect 5724 3690 5742 3708
rect 5724 3708 5742 3726
rect 5724 3726 5742 3744
rect 5724 3744 5742 3762
rect 5724 3762 5742 3780
rect 5724 3780 5742 3798
rect 5724 3798 5742 3816
rect 5724 3816 5742 3834
rect 5724 3834 5742 3852
rect 5724 3852 5742 3870
rect 5724 3870 5742 3888
rect 5724 3888 5742 3906
rect 5724 3906 5742 3924
rect 5724 3924 5742 3942
rect 5724 3942 5742 3960
rect 5724 3960 5742 3978
rect 5724 3978 5742 3996
rect 5724 3996 5742 4014
rect 5724 4014 5742 4032
rect 5724 4032 5742 4050
rect 5724 4050 5742 4068
rect 5724 4068 5742 4086
rect 5724 4086 5742 4104
rect 5724 4104 5742 4122
rect 5724 4122 5742 4140
rect 5724 4140 5742 4158
rect 5724 4158 5742 4176
rect 5724 4176 5742 4194
rect 5724 4194 5742 4212
rect 5724 4212 5742 4230
rect 5724 4230 5742 4248
rect 5724 4248 5742 4266
rect 5724 4266 5742 4284
rect 5724 4284 5742 4302
rect 5724 4302 5742 4320
rect 5724 4320 5742 4338
rect 5724 4338 5742 4356
rect 5724 4356 5742 4374
rect 5724 4374 5742 4392
rect 5724 4392 5742 4410
rect 5724 4410 5742 4428
rect 5724 4428 5742 4446
rect 5724 4446 5742 4464
rect 5724 4464 5742 4482
rect 5724 4482 5742 4500
rect 5724 4500 5742 4518
rect 5724 4518 5742 4536
rect 5724 4536 5742 4554
rect 5724 4554 5742 4572
rect 5724 4572 5742 4590
rect 5724 4590 5742 4608
rect 5724 4608 5742 4626
rect 5724 4626 5742 4644
rect 5724 4644 5742 4662
rect 5724 4662 5742 4680
rect 5724 4680 5742 4698
rect 5724 4698 5742 4716
rect 5724 4716 5742 4734
rect 5724 4734 5742 4752
rect 5724 4752 5742 4770
rect 5724 4770 5742 4788
rect 5724 4788 5742 4806
rect 5724 4806 5742 4824
rect 5724 4824 5742 4842
rect 5724 4842 5742 4860
rect 5724 4860 5742 4878
rect 5724 4878 5742 4896
rect 5724 4896 5742 4914
rect 5724 4914 5742 4932
rect 5724 4932 5742 4950
rect 5724 4950 5742 4968
rect 5724 4968 5742 4986
rect 5724 4986 5742 5004
rect 5724 5004 5742 5022
rect 5724 5022 5742 5040
rect 5724 5040 5742 5058
rect 5724 5058 5742 5076
rect 5724 5076 5742 5094
rect 5724 5094 5742 5112
rect 5724 5112 5742 5130
rect 5724 5346 5742 5364
rect 5724 5364 5742 5382
rect 5724 5382 5742 5400
rect 5724 5400 5742 5418
rect 5724 5418 5742 5436
rect 5724 5436 5742 5454
rect 5724 5454 5742 5472
rect 5724 5472 5742 5490
rect 5724 5490 5742 5508
rect 5724 5508 5742 5526
rect 5724 5526 5742 5544
rect 5724 5544 5742 5562
rect 5724 5562 5742 5580
rect 5724 5580 5742 5598
rect 5724 5598 5742 5616
rect 5724 5616 5742 5634
rect 5724 5634 5742 5652
rect 5724 5652 5742 5670
rect 5724 5670 5742 5688
rect 5724 5688 5742 5706
rect 5724 5706 5742 5724
rect 5724 5724 5742 5742
rect 5724 5742 5742 5760
rect 5724 5760 5742 5778
rect 5724 5778 5742 5796
rect 5724 5796 5742 5814
rect 5724 5814 5742 5832
rect 5724 5832 5742 5850
rect 5724 5850 5742 5868
rect 5724 5868 5742 5886
rect 5724 5886 5742 5904
rect 5724 5904 5742 5922
rect 5724 5922 5742 5940
rect 5724 5940 5742 5958
rect 5724 5958 5742 5976
rect 5724 5976 5742 5994
rect 5724 5994 5742 6012
rect 5724 6012 5742 6030
rect 5724 6030 5742 6048
rect 5724 6048 5742 6066
rect 5724 6066 5742 6084
rect 5724 6084 5742 6102
rect 5724 6102 5742 6120
rect 5724 6120 5742 6138
rect 5724 6138 5742 6156
rect 5724 6156 5742 6174
rect 5724 6174 5742 6192
rect 5724 6192 5742 6210
rect 5724 6210 5742 6228
rect 5724 6228 5742 6246
rect 5724 6246 5742 6264
rect 5724 6264 5742 6282
rect 5724 6282 5742 6300
rect 5724 6300 5742 6318
rect 5724 6318 5742 6336
rect 5724 6336 5742 6354
rect 5724 6354 5742 6372
rect 5724 6372 5742 6390
rect 5724 6390 5742 6408
rect 5724 6408 5742 6426
rect 5724 6426 5742 6444
rect 5724 6444 5742 6462
rect 5724 6462 5742 6480
rect 5724 6480 5742 6498
rect 5724 6498 5742 6516
rect 5724 6516 5742 6534
rect 5724 6534 5742 6552
rect 5724 6552 5742 6570
rect 5724 6570 5742 6588
rect 5724 6588 5742 6606
rect 5724 6606 5742 6624
rect 5724 6624 5742 6642
rect 5724 6642 5742 6660
rect 5724 6660 5742 6678
rect 5724 6678 5742 6696
rect 5724 6696 5742 6714
rect 5724 6714 5742 6732
rect 5724 6732 5742 6750
rect 5724 6750 5742 6768
rect 5724 6768 5742 6786
rect 5724 6786 5742 6804
rect 5724 6804 5742 6822
rect 5724 6822 5742 6840
rect 5724 6840 5742 6858
rect 5724 6858 5742 6876
rect 5724 6876 5742 6894
rect 5724 6894 5742 6912
rect 5724 6912 5742 6930
rect 5724 6930 5742 6948
rect 5724 6948 5742 6966
rect 5724 6966 5742 6984
rect 5724 6984 5742 7002
rect 5724 7002 5742 7020
rect 5724 7020 5742 7038
rect 5724 7038 5742 7056
rect 5724 7056 5742 7074
rect 5724 7074 5742 7092
rect 5724 7092 5742 7110
rect 5724 7110 5742 7128
rect 5724 7128 5742 7146
rect 5724 7146 5742 7164
rect 5724 7164 5742 7182
rect 5724 7182 5742 7200
rect 5724 7200 5742 7218
rect 5724 7218 5742 7236
rect 5724 7236 5742 7254
rect 5724 7254 5742 7272
rect 5724 7272 5742 7290
rect 5724 7290 5742 7308
rect 5724 7308 5742 7326
rect 5724 7326 5742 7344
rect 5724 7344 5742 7362
rect 5724 7362 5742 7380
rect 5724 7380 5742 7398
rect 5724 7398 5742 7416
rect 5724 7416 5742 7434
rect 5724 7434 5742 7452
rect 5724 7452 5742 7470
rect 5724 7470 5742 7488
rect 5724 7488 5742 7506
rect 5724 7506 5742 7524
rect 5724 7524 5742 7542
rect 5724 7542 5742 7560
rect 5724 7560 5742 7578
rect 5724 7578 5742 7596
rect 5724 7596 5742 7614
rect 5724 7614 5742 7632
rect 5724 7632 5742 7650
rect 5724 7650 5742 7668
rect 5724 7668 5742 7686
rect 5724 7686 5742 7704
rect 5724 7704 5742 7722
rect 5724 7722 5742 7740
rect 5724 7740 5742 7758
rect 5724 7758 5742 7776
rect 5724 7776 5742 7794
rect 5724 7794 5742 7812
rect 5724 7812 5742 7830
rect 5724 7830 5742 7848
rect 5724 7848 5742 7866
rect 5724 7866 5742 7884
rect 5724 7884 5742 7902
rect 5724 7902 5742 7920
rect 5724 7920 5742 7938
rect 5724 7938 5742 7956
rect 5724 7956 5742 7974
rect 5724 7974 5742 7992
rect 5724 7992 5742 8010
rect 5724 8010 5742 8028
rect 5724 8028 5742 8046
rect 5724 8046 5742 8064
rect 5724 8064 5742 8082
rect 5724 8082 5742 8100
rect 5724 8100 5742 8118
rect 5724 8118 5742 8136
rect 5724 8136 5742 8154
rect 5724 8154 5742 8172
rect 5724 8172 5742 8190
rect 5724 8190 5742 8208
rect 5724 8208 5742 8226
rect 5724 8226 5742 8244
rect 5724 8244 5742 8262
rect 5724 8262 5742 8280
rect 5724 8280 5742 8298
rect 5724 8298 5742 8316
rect 5724 8316 5742 8334
rect 5724 8334 5742 8352
rect 5724 8352 5742 8370
rect 5724 8370 5742 8388
rect 5724 8388 5742 8406
rect 5724 8406 5742 8424
rect 5724 8424 5742 8442
rect 5724 8442 5742 8460
rect 5724 8460 5742 8478
rect 5724 8478 5742 8496
rect 5724 8496 5742 8514
rect 5724 8514 5742 8532
rect 5724 8532 5742 8550
rect 5724 8550 5742 8568
rect 5724 8568 5742 8586
rect 5724 8586 5742 8604
rect 5724 8604 5742 8622
rect 5724 8622 5742 8640
rect 5724 8640 5742 8658
rect 5724 8658 5742 8676
rect 5724 8676 5742 8694
rect 5724 8694 5742 8712
rect 5724 8712 5742 8730
rect 5724 8730 5742 8748
rect 5724 8748 5742 8766
rect 5724 8766 5742 8784
rect 5724 8784 5742 8802
rect 5724 8802 5742 8820
rect 5724 8820 5742 8838
rect 5724 8838 5742 8856
rect 5724 8856 5742 8874
rect 5742 702 5760 720
rect 5742 720 5760 738
rect 5742 738 5760 756
rect 5742 756 5760 774
rect 5742 774 5760 792
rect 5742 792 5760 810
rect 5742 810 5760 828
rect 5742 828 5760 846
rect 5742 846 5760 864
rect 5742 864 5760 882
rect 5742 882 5760 900
rect 5742 900 5760 918
rect 5742 918 5760 936
rect 5742 936 5760 954
rect 5742 954 5760 972
rect 5742 972 5760 990
rect 5742 990 5760 1008
rect 5742 1152 5760 1170
rect 5742 1170 5760 1188
rect 5742 1188 5760 1206
rect 5742 1206 5760 1224
rect 5742 1224 5760 1242
rect 5742 1242 5760 1260
rect 5742 1260 5760 1278
rect 5742 1278 5760 1296
rect 5742 1296 5760 1314
rect 5742 1314 5760 1332
rect 5742 1332 5760 1350
rect 5742 1350 5760 1368
rect 5742 1368 5760 1386
rect 5742 1386 5760 1404
rect 5742 1404 5760 1422
rect 5742 1422 5760 1440
rect 5742 1440 5760 1458
rect 5742 1458 5760 1476
rect 5742 1476 5760 1494
rect 5742 1494 5760 1512
rect 5742 1512 5760 1530
rect 5742 1530 5760 1548
rect 5742 1548 5760 1566
rect 5742 1566 5760 1584
rect 5742 1584 5760 1602
rect 5742 1602 5760 1620
rect 5742 1620 5760 1638
rect 5742 1638 5760 1656
rect 5742 1656 5760 1674
rect 5742 1674 5760 1692
rect 5742 1692 5760 1710
rect 5742 1710 5760 1728
rect 5742 1728 5760 1746
rect 5742 1746 5760 1764
rect 5742 1764 5760 1782
rect 5742 1782 5760 1800
rect 5742 1800 5760 1818
rect 5742 1818 5760 1836
rect 5742 1836 5760 1854
rect 5742 1854 5760 1872
rect 5742 1872 5760 1890
rect 5742 1890 5760 1908
rect 5742 1908 5760 1926
rect 5742 1926 5760 1944
rect 5742 1944 5760 1962
rect 5742 1962 5760 1980
rect 5742 1980 5760 1998
rect 5742 1998 5760 2016
rect 5742 2016 5760 2034
rect 5742 2034 5760 2052
rect 5742 2052 5760 2070
rect 5742 2070 5760 2088
rect 5742 2088 5760 2106
rect 5742 2106 5760 2124
rect 5742 2124 5760 2142
rect 5742 2142 5760 2160
rect 5742 2160 5760 2178
rect 5742 2178 5760 2196
rect 5742 2196 5760 2214
rect 5742 2214 5760 2232
rect 5742 2232 5760 2250
rect 5742 2250 5760 2268
rect 5742 2268 5760 2286
rect 5742 2286 5760 2304
rect 5742 2304 5760 2322
rect 5742 2322 5760 2340
rect 5742 2340 5760 2358
rect 5742 2358 5760 2376
rect 5742 2376 5760 2394
rect 5742 2394 5760 2412
rect 5742 2412 5760 2430
rect 5742 2430 5760 2448
rect 5742 2448 5760 2466
rect 5742 2466 5760 2484
rect 5742 2484 5760 2502
rect 5742 2502 5760 2520
rect 5742 2520 5760 2538
rect 5742 2538 5760 2556
rect 5742 2556 5760 2574
rect 5742 2574 5760 2592
rect 5742 2592 5760 2610
rect 5742 2610 5760 2628
rect 5742 2844 5760 2862
rect 5742 2862 5760 2880
rect 5742 2880 5760 2898
rect 5742 2898 5760 2916
rect 5742 2916 5760 2934
rect 5742 2934 5760 2952
rect 5742 2952 5760 2970
rect 5742 2970 5760 2988
rect 5742 2988 5760 3006
rect 5742 3006 5760 3024
rect 5742 3024 5760 3042
rect 5742 3042 5760 3060
rect 5742 3060 5760 3078
rect 5742 3078 5760 3096
rect 5742 3096 5760 3114
rect 5742 3114 5760 3132
rect 5742 3132 5760 3150
rect 5742 3150 5760 3168
rect 5742 3168 5760 3186
rect 5742 3186 5760 3204
rect 5742 3204 5760 3222
rect 5742 3222 5760 3240
rect 5742 3240 5760 3258
rect 5742 3258 5760 3276
rect 5742 3276 5760 3294
rect 5742 3294 5760 3312
rect 5742 3312 5760 3330
rect 5742 3330 5760 3348
rect 5742 3348 5760 3366
rect 5742 3366 5760 3384
rect 5742 3384 5760 3402
rect 5742 3402 5760 3420
rect 5742 3420 5760 3438
rect 5742 3438 5760 3456
rect 5742 3456 5760 3474
rect 5742 3474 5760 3492
rect 5742 3492 5760 3510
rect 5742 3510 5760 3528
rect 5742 3528 5760 3546
rect 5742 3546 5760 3564
rect 5742 3564 5760 3582
rect 5742 3582 5760 3600
rect 5742 3600 5760 3618
rect 5742 3618 5760 3636
rect 5742 3636 5760 3654
rect 5742 3654 5760 3672
rect 5742 3672 5760 3690
rect 5742 3690 5760 3708
rect 5742 3708 5760 3726
rect 5742 3726 5760 3744
rect 5742 3744 5760 3762
rect 5742 3762 5760 3780
rect 5742 3780 5760 3798
rect 5742 3798 5760 3816
rect 5742 3816 5760 3834
rect 5742 3834 5760 3852
rect 5742 3852 5760 3870
rect 5742 3870 5760 3888
rect 5742 3888 5760 3906
rect 5742 3906 5760 3924
rect 5742 3924 5760 3942
rect 5742 3942 5760 3960
rect 5742 3960 5760 3978
rect 5742 3978 5760 3996
rect 5742 3996 5760 4014
rect 5742 4014 5760 4032
rect 5742 4032 5760 4050
rect 5742 4050 5760 4068
rect 5742 4068 5760 4086
rect 5742 4086 5760 4104
rect 5742 4104 5760 4122
rect 5742 4122 5760 4140
rect 5742 4140 5760 4158
rect 5742 4158 5760 4176
rect 5742 4176 5760 4194
rect 5742 4194 5760 4212
rect 5742 4212 5760 4230
rect 5742 4230 5760 4248
rect 5742 4248 5760 4266
rect 5742 4266 5760 4284
rect 5742 4284 5760 4302
rect 5742 4302 5760 4320
rect 5742 4320 5760 4338
rect 5742 4338 5760 4356
rect 5742 4356 5760 4374
rect 5742 4374 5760 4392
rect 5742 4392 5760 4410
rect 5742 4410 5760 4428
rect 5742 4428 5760 4446
rect 5742 4446 5760 4464
rect 5742 4464 5760 4482
rect 5742 4482 5760 4500
rect 5742 4500 5760 4518
rect 5742 4518 5760 4536
rect 5742 4536 5760 4554
rect 5742 4554 5760 4572
rect 5742 4572 5760 4590
rect 5742 4590 5760 4608
rect 5742 4608 5760 4626
rect 5742 4626 5760 4644
rect 5742 4644 5760 4662
rect 5742 4662 5760 4680
rect 5742 4680 5760 4698
rect 5742 4698 5760 4716
rect 5742 4716 5760 4734
rect 5742 4734 5760 4752
rect 5742 4752 5760 4770
rect 5742 4770 5760 4788
rect 5742 4788 5760 4806
rect 5742 4806 5760 4824
rect 5742 4824 5760 4842
rect 5742 4842 5760 4860
rect 5742 4860 5760 4878
rect 5742 4878 5760 4896
rect 5742 4896 5760 4914
rect 5742 4914 5760 4932
rect 5742 4932 5760 4950
rect 5742 4950 5760 4968
rect 5742 4968 5760 4986
rect 5742 4986 5760 5004
rect 5742 5004 5760 5022
rect 5742 5022 5760 5040
rect 5742 5040 5760 5058
rect 5742 5058 5760 5076
rect 5742 5076 5760 5094
rect 5742 5094 5760 5112
rect 5742 5112 5760 5130
rect 5742 5364 5760 5382
rect 5742 5382 5760 5400
rect 5742 5400 5760 5418
rect 5742 5418 5760 5436
rect 5742 5436 5760 5454
rect 5742 5454 5760 5472
rect 5742 5472 5760 5490
rect 5742 5490 5760 5508
rect 5742 5508 5760 5526
rect 5742 5526 5760 5544
rect 5742 5544 5760 5562
rect 5742 5562 5760 5580
rect 5742 5580 5760 5598
rect 5742 5598 5760 5616
rect 5742 5616 5760 5634
rect 5742 5634 5760 5652
rect 5742 5652 5760 5670
rect 5742 5670 5760 5688
rect 5742 5688 5760 5706
rect 5742 5706 5760 5724
rect 5742 5724 5760 5742
rect 5742 5742 5760 5760
rect 5742 5760 5760 5778
rect 5742 5778 5760 5796
rect 5742 5796 5760 5814
rect 5742 5814 5760 5832
rect 5742 5832 5760 5850
rect 5742 5850 5760 5868
rect 5742 5868 5760 5886
rect 5742 5886 5760 5904
rect 5742 5904 5760 5922
rect 5742 5922 5760 5940
rect 5742 5940 5760 5958
rect 5742 5958 5760 5976
rect 5742 5976 5760 5994
rect 5742 5994 5760 6012
rect 5742 6012 5760 6030
rect 5742 6030 5760 6048
rect 5742 6048 5760 6066
rect 5742 6066 5760 6084
rect 5742 6084 5760 6102
rect 5742 6102 5760 6120
rect 5742 6120 5760 6138
rect 5742 6138 5760 6156
rect 5742 6156 5760 6174
rect 5742 6174 5760 6192
rect 5742 6192 5760 6210
rect 5742 6210 5760 6228
rect 5742 6228 5760 6246
rect 5742 6246 5760 6264
rect 5742 6264 5760 6282
rect 5742 6282 5760 6300
rect 5742 6300 5760 6318
rect 5742 6318 5760 6336
rect 5742 6336 5760 6354
rect 5742 6354 5760 6372
rect 5742 6372 5760 6390
rect 5742 6390 5760 6408
rect 5742 6408 5760 6426
rect 5742 6426 5760 6444
rect 5742 6444 5760 6462
rect 5742 6462 5760 6480
rect 5742 6480 5760 6498
rect 5742 6498 5760 6516
rect 5742 6516 5760 6534
rect 5742 6534 5760 6552
rect 5742 6552 5760 6570
rect 5742 6570 5760 6588
rect 5742 6588 5760 6606
rect 5742 6606 5760 6624
rect 5742 6624 5760 6642
rect 5742 6642 5760 6660
rect 5742 6660 5760 6678
rect 5742 6678 5760 6696
rect 5742 6696 5760 6714
rect 5742 6714 5760 6732
rect 5742 6732 5760 6750
rect 5742 6750 5760 6768
rect 5742 6768 5760 6786
rect 5742 6786 5760 6804
rect 5742 6804 5760 6822
rect 5742 6822 5760 6840
rect 5742 6840 5760 6858
rect 5742 6858 5760 6876
rect 5742 6876 5760 6894
rect 5742 6894 5760 6912
rect 5742 6912 5760 6930
rect 5742 6930 5760 6948
rect 5742 6948 5760 6966
rect 5742 6966 5760 6984
rect 5742 6984 5760 7002
rect 5742 7002 5760 7020
rect 5742 7020 5760 7038
rect 5742 7038 5760 7056
rect 5742 7056 5760 7074
rect 5742 7074 5760 7092
rect 5742 7092 5760 7110
rect 5742 7110 5760 7128
rect 5742 7128 5760 7146
rect 5742 7146 5760 7164
rect 5742 7164 5760 7182
rect 5742 7182 5760 7200
rect 5742 7200 5760 7218
rect 5742 7218 5760 7236
rect 5742 7236 5760 7254
rect 5742 7254 5760 7272
rect 5742 7272 5760 7290
rect 5742 7290 5760 7308
rect 5742 7308 5760 7326
rect 5742 7326 5760 7344
rect 5742 7344 5760 7362
rect 5742 7362 5760 7380
rect 5742 7380 5760 7398
rect 5742 7398 5760 7416
rect 5742 7416 5760 7434
rect 5742 7434 5760 7452
rect 5742 7452 5760 7470
rect 5742 7470 5760 7488
rect 5742 7488 5760 7506
rect 5742 7506 5760 7524
rect 5742 7524 5760 7542
rect 5742 7542 5760 7560
rect 5742 7560 5760 7578
rect 5742 7578 5760 7596
rect 5742 7596 5760 7614
rect 5742 7614 5760 7632
rect 5742 7632 5760 7650
rect 5742 7650 5760 7668
rect 5742 7668 5760 7686
rect 5742 7686 5760 7704
rect 5742 7704 5760 7722
rect 5742 7722 5760 7740
rect 5742 7740 5760 7758
rect 5742 7758 5760 7776
rect 5742 7776 5760 7794
rect 5742 7794 5760 7812
rect 5742 7812 5760 7830
rect 5742 7830 5760 7848
rect 5742 7848 5760 7866
rect 5742 7866 5760 7884
rect 5742 7884 5760 7902
rect 5742 7902 5760 7920
rect 5742 7920 5760 7938
rect 5742 7938 5760 7956
rect 5742 7956 5760 7974
rect 5742 7974 5760 7992
rect 5742 7992 5760 8010
rect 5742 8010 5760 8028
rect 5742 8028 5760 8046
rect 5742 8046 5760 8064
rect 5742 8064 5760 8082
rect 5742 8082 5760 8100
rect 5742 8100 5760 8118
rect 5742 8118 5760 8136
rect 5742 8136 5760 8154
rect 5742 8154 5760 8172
rect 5742 8172 5760 8190
rect 5742 8190 5760 8208
rect 5742 8208 5760 8226
rect 5742 8226 5760 8244
rect 5742 8244 5760 8262
rect 5742 8262 5760 8280
rect 5742 8280 5760 8298
rect 5742 8298 5760 8316
rect 5742 8316 5760 8334
rect 5742 8334 5760 8352
rect 5742 8352 5760 8370
rect 5742 8370 5760 8388
rect 5742 8388 5760 8406
rect 5742 8406 5760 8424
rect 5742 8424 5760 8442
rect 5742 8442 5760 8460
rect 5742 8460 5760 8478
rect 5742 8478 5760 8496
rect 5742 8496 5760 8514
rect 5742 8514 5760 8532
rect 5742 8532 5760 8550
rect 5742 8550 5760 8568
rect 5742 8568 5760 8586
rect 5742 8586 5760 8604
rect 5742 8604 5760 8622
rect 5742 8622 5760 8640
rect 5742 8640 5760 8658
rect 5742 8658 5760 8676
rect 5742 8676 5760 8694
rect 5742 8694 5760 8712
rect 5742 8712 5760 8730
rect 5742 8730 5760 8748
rect 5742 8748 5760 8766
rect 5742 8766 5760 8784
rect 5742 8784 5760 8802
rect 5742 8802 5760 8820
rect 5742 8820 5760 8838
rect 5742 8838 5760 8856
rect 5742 8856 5760 8874
rect 5742 8874 5760 8892
rect 5760 702 5778 720
rect 5760 720 5778 738
rect 5760 738 5778 756
rect 5760 756 5778 774
rect 5760 774 5778 792
rect 5760 792 5778 810
rect 5760 810 5778 828
rect 5760 828 5778 846
rect 5760 846 5778 864
rect 5760 864 5778 882
rect 5760 882 5778 900
rect 5760 900 5778 918
rect 5760 918 5778 936
rect 5760 936 5778 954
rect 5760 954 5778 972
rect 5760 972 5778 990
rect 5760 990 5778 1008
rect 5760 1008 5778 1026
rect 5760 1152 5778 1170
rect 5760 1170 5778 1188
rect 5760 1188 5778 1206
rect 5760 1206 5778 1224
rect 5760 1224 5778 1242
rect 5760 1242 5778 1260
rect 5760 1260 5778 1278
rect 5760 1278 5778 1296
rect 5760 1296 5778 1314
rect 5760 1314 5778 1332
rect 5760 1332 5778 1350
rect 5760 1350 5778 1368
rect 5760 1368 5778 1386
rect 5760 1386 5778 1404
rect 5760 1404 5778 1422
rect 5760 1422 5778 1440
rect 5760 1440 5778 1458
rect 5760 1458 5778 1476
rect 5760 1476 5778 1494
rect 5760 1494 5778 1512
rect 5760 1512 5778 1530
rect 5760 1530 5778 1548
rect 5760 1548 5778 1566
rect 5760 1566 5778 1584
rect 5760 1584 5778 1602
rect 5760 1602 5778 1620
rect 5760 1620 5778 1638
rect 5760 1638 5778 1656
rect 5760 1656 5778 1674
rect 5760 1674 5778 1692
rect 5760 1692 5778 1710
rect 5760 1710 5778 1728
rect 5760 1728 5778 1746
rect 5760 1746 5778 1764
rect 5760 1764 5778 1782
rect 5760 1782 5778 1800
rect 5760 1800 5778 1818
rect 5760 1818 5778 1836
rect 5760 1836 5778 1854
rect 5760 1854 5778 1872
rect 5760 1872 5778 1890
rect 5760 1890 5778 1908
rect 5760 1908 5778 1926
rect 5760 1926 5778 1944
rect 5760 1944 5778 1962
rect 5760 1962 5778 1980
rect 5760 1980 5778 1998
rect 5760 1998 5778 2016
rect 5760 2016 5778 2034
rect 5760 2034 5778 2052
rect 5760 2052 5778 2070
rect 5760 2070 5778 2088
rect 5760 2088 5778 2106
rect 5760 2106 5778 2124
rect 5760 2124 5778 2142
rect 5760 2142 5778 2160
rect 5760 2160 5778 2178
rect 5760 2178 5778 2196
rect 5760 2196 5778 2214
rect 5760 2214 5778 2232
rect 5760 2232 5778 2250
rect 5760 2250 5778 2268
rect 5760 2268 5778 2286
rect 5760 2286 5778 2304
rect 5760 2304 5778 2322
rect 5760 2322 5778 2340
rect 5760 2340 5778 2358
rect 5760 2358 5778 2376
rect 5760 2376 5778 2394
rect 5760 2394 5778 2412
rect 5760 2412 5778 2430
rect 5760 2430 5778 2448
rect 5760 2448 5778 2466
rect 5760 2466 5778 2484
rect 5760 2484 5778 2502
rect 5760 2502 5778 2520
rect 5760 2520 5778 2538
rect 5760 2538 5778 2556
rect 5760 2556 5778 2574
rect 5760 2574 5778 2592
rect 5760 2592 5778 2610
rect 5760 2610 5778 2628
rect 5760 2628 5778 2646
rect 5760 2862 5778 2880
rect 5760 2880 5778 2898
rect 5760 2898 5778 2916
rect 5760 2916 5778 2934
rect 5760 2934 5778 2952
rect 5760 2952 5778 2970
rect 5760 2970 5778 2988
rect 5760 2988 5778 3006
rect 5760 3006 5778 3024
rect 5760 3024 5778 3042
rect 5760 3042 5778 3060
rect 5760 3060 5778 3078
rect 5760 3078 5778 3096
rect 5760 3096 5778 3114
rect 5760 3114 5778 3132
rect 5760 3132 5778 3150
rect 5760 3150 5778 3168
rect 5760 3168 5778 3186
rect 5760 3186 5778 3204
rect 5760 3204 5778 3222
rect 5760 3222 5778 3240
rect 5760 3240 5778 3258
rect 5760 3258 5778 3276
rect 5760 3276 5778 3294
rect 5760 3294 5778 3312
rect 5760 3312 5778 3330
rect 5760 3330 5778 3348
rect 5760 3348 5778 3366
rect 5760 3366 5778 3384
rect 5760 3384 5778 3402
rect 5760 3402 5778 3420
rect 5760 3420 5778 3438
rect 5760 3438 5778 3456
rect 5760 3456 5778 3474
rect 5760 3474 5778 3492
rect 5760 3492 5778 3510
rect 5760 3510 5778 3528
rect 5760 3528 5778 3546
rect 5760 3546 5778 3564
rect 5760 3564 5778 3582
rect 5760 3582 5778 3600
rect 5760 3600 5778 3618
rect 5760 3618 5778 3636
rect 5760 3636 5778 3654
rect 5760 3654 5778 3672
rect 5760 3672 5778 3690
rect 5760 3690 5778 3708
rect 5760 3708 5778 3726
rect 5760 3726 5778 3744
rect 5760 3744 5778 3762
rect 5760 3762 5778 3780
rect 5760 3780 5778 3798
rect 5760 3798 5778 3816
rect 5760 3816 5778 3834
rect 5760 3834 5778 3852
rect 5760 3852 5778 3870
rect 5760 3870 5778 3888
rect 5760 3888 5778 3906
rect 5760 3906 5778 3924
rect 5760 3924 5778 3942
rect 5760 3942 5778 3960
rect 5760 3960 5778 3978
rect 5760 3978 5778 3996
rect 5760 3996 5778 4014
rect 5760 4014 5778 4032
rect 5760 4032 5778 4050
rect 5760 4050 5778 4068
rect 5760 4068 5778 4086
rect 5760 4086 5778 4104
rect 5760 4104 5778 4122
rect 5760 4122 5778 4140
rect 5760 4140 5778 4158
rect 5760 4158 5778 4176
rect 5760 4176 5778 4194
rect 5760 4194 5778 4212
rect 5760 4212 5778 4230
rect 5760 4230 5778 4248
rect 5760 4248 5778 4266
rect 5760 4266 5778 4284
rect 5760 4284 5778 4302
rect 5760 4302 5778 4320
rect 5760 4320 5778 4338
rect 5760 4338 5778 4356
rect 5760 4356 5778 4374
rect 5760 4374 5778 4392
rect 5760 4392 5778 4410
rect 5760 4410 5778 4428
rect 5760 4428 5778 4446
rect 5760 4446 5778 4464
rect 5760 4464 5778 4482
rect 5760 4482 5778 4500
rect 5760 4500 5778 4518
rect 5760 4518 5778 4536
rect 5760 4536 5778 4554
rect 5760 4554 5778 4572
rect 5760 4572 5778 4590
rect 5760 4590 5778 4608
rect 5760 4608 5778 4626
rect 5760 4626 5778 4644
rect 5760 4644 5778 4662
rect 5760 4662 5778 4680
rect 5760 4680 5778 4698
rect 5760 4698 5778 4716
rect 5760 4716 5778 4734
rect 5760 4734 5778 4752
rect 5760 4752 5778 4770
rect 5760 4770 5778 4788
rect 5760 4788 5778 4806
rect 5760 4806 5778 4824
rect 5760 4824 5778 4842
rect 5760 4842 5778 4860
rect 5760 4860 5778 4878
rect 5760 4878 5778 4896
rect 5760 4896 5778 4914
rect 5760 4914 5778 4932
rect 5760 4932 5778 4950
rect 5760 4950 5778 4968
rect 5760 4968 5778 4986
rect 5760 4986 5778 5004
rect 5760 5004 5778 5022
rect 5760 5022 5778 5040
rect 5760 5040 5778 5058
rect 5760 5058 5778 5076
rect 5760 5076 5778 5094
rect 5760 5094 5778 5112
rect 5760 5112 5778 5130
rect 5760 5130 5778 5148
rect 5760 5382 5778 5400
rect 5760 5400 5778 5418
rect 5760 5418 5778 5436
rect 5760 5436 5778 5454
rect 5760 5454 5778 5472
rect 5760 5472 5778 5490
rect 5760 5490 5778 5508
rect 5760 5508 5778 5526
rect 5760 5526 5778 5544
rect 5760 5544 5778 5562
rect 5760 5562 5778 5580
rect 5760 5580 5778 5598
rect 5760 5598 5778 5616
rect 5760 5616 5778 5634
rect 5760 5634 5778 5652
rect 5760 5652 5778 5670
rect 5760 5670 5778 5688
rect 5760 5688 5778 5706
rect 5760 5706 5778 5724
rect 5760 5724 5778 5742
rect 5760 5742 5778 5760
rect 5760 5760 5778 5778
rect 5760 5778 5778 5796
rect 5760 5796 5778 5814
rect 5760 5814 5778 5832
rect 5760 5832 5778 5850
rect 5760 5850 5778 5868
rect 5760 5868 5778 5886
rect 5760 5886 5778 5904
rect 5760 5904 5778 5922
rect 5760 5922 5778 5940
rect 5760 5940 5778 5958
rect 5760 5958 5778 5976
rect 5760 5976 5778 5994
rect 5760 5994 5778 6012
rect 5760 6012 5778 6030
rect 5760 6030 5778 6048
rect 5760 6048 5778 6066
rect 5760 6066 5778 6084
rect 5760 6084 5778 6102
rect 5760 6102 5778 6120
rect 5760 6120 5778 6138
rect 5760 6138 5778 6156
rect 5760 6156 5778 6174
rect 5760 6174 5778 6192
rect 5760 6192 5778 6210
rect 5760 6210 5778 6228
rect 5760 6228 5778 6246
rect 5760 6246 5778 6264
rect 5760 6264 5778 6282
rect 5760 6282 5778 6300
rect 5760 6300 5778 6318
rect 5760 6318 5778 6336
rect 5760 6336 5778 6354
rect 5760 6354 5778 6372
rect 5760 6372 5778 6390
rect 5760 6390 5778 6408
rect 5760 6408 5778 6426
rect 5760 6426 5778 6444
rect 5760 6444 5778 6462
rect 5760 6462 5778 6480
rect 5760 6480 5778 6498
rect 5760 6498 5778 6516
rect 5760 6516 5778 6534
rect 5760 6534 5778 6552
rect 5760 6552 5778 6570
rect 5760 6570 5778 6588
rect 5760 6588 5778 6606
rect 5760 6606 5778 6624
rect 5760 6624 5778 6642
rect 5760 6642 5778 6660
rect 5760 6660 5778 6678
rect 5760 6678 5778 6696
rect 5760 6696 5778 6714
rect 5760 6714 5778 6732
rect 5760 6732 5778 6750
rect 5760 6750 5778 6768
rect 5760 6768 5778 6786
rect 5760 6786 5778 6804
rect 5760 6804 5778 6822
rect 5760 6822 5778 6840
rect 5760 6840 5778 6858
rect 5760 6858 5778 6876
rect 5760 6876 5778 6894
rect 5760 6894 5778 6912
rect 5760 6912 5778 6930
rect 5760 6930 5778 6948
rect 5760 6948 5778 6966
rect 5760 6966 5778 6984
rect 5760 6984 5778 7002
rect 5760 7002 5778 7020
rect 5760 7020 5778 7038
rect 5760 7038 5778 7056
rect 5760 7056 5778 7074
rect 5760 7074 5778 7092
rect 5760 7092 5778 7110
rect 5760 7110 5778 7128
rect 5760 7128 5778 7146
rect 5760 7146 5778 7164
rect 5760 7164 5778 7182
rect 5760 7182 5778 7200
rect 5760 7200 5778 7218
rect 5760 7218 5778 7236
rect 5760 7236 5778 7254
rect 5760 7254 5778 7272
rect 5760 7272 5778 7290
rect 5760 7290 5778 7308
rect 5760 7308 5778 7326
rect 5760 7326 5778 7344
rect 5760 7344 5778 7362
rect 5760 7362 5778 7380
rect 5760 7380 5778 7398
rect 5760 7398 5778 7416
rect 5760 7416 5778 7434
rect 5760 7434 5778 7452
rect 5760 7452 5778 7470
rect 5760 7470 5778 7488
rect 5760 7488 5778 7506
rect 5760 7506 5778 7524
rect 5760 7524 5778 7542
rect 5760 7542 5778 7560
rect 5760 7560 5778 7578
rect 5760 7578 5778 7596
rect 5760 7596 5778 7614
rect 5760 7614 5778 7632
rect 5760 7632 5778 7650
rect 5760 7650 5778 7668
rect 5760 7668 5778 7686
rect 5760 7686 5778 7704
rect 5760 7704 5778 7722
rect 5760 7722 5778 7740
rect 5760 7740 5778 7758
rect 5760 7758 5778 7776
rect 5760 7776 5778 7794
rect 5760 7794 5778 7812
rect 5760 7812 5778 7830
rect 5760 7830 5778 7848
rect 5760 7848 5778 7866
rect 5760 7866 5778 7884
rect 5760 7884 5778 7902
rect 5760 7902 5778 7920
rect 5760 7920 5778 7938
rect 5760 7938 5778 7956
rect 5760 7956 5778 7974
rect 5760 7974 5778 7992
rect 5760 7992 5778 8010
rect 5760 8010 5778 8028
rect 5760 8028 5778 8046
rect 5760 8046 5778 8064
rect 5760 8064 5778 8082
rect 5760 8082 5778 8100
rect 5760 8100 5778 8118
rect 5760 8118 5778 8136
rect 5760 8136 5778 8154
rect 5760 8154 5778 8172
rect 5760 8172 5778 8190
rect 5760 8190 5778 8208
rect 5760 8208 5778 8226
rect 5760 8226 5778 8244
rect 5760 8244 5778 8262
rect 5760 8262 5778 8280
rect 5760 8280 5778 8298
rect 5760 8298 5778 8316
rect 5760 8316 5778 8334
rect 5760 8334 5778 8352
rect 5760 8352 5778 8370
rect 5760 8370 5778 8388
rect 5760 8388 5778 8406
rect 5760 8406 5778 8424
rect 5760 8424 5778 8442
rect 5760 8442 5778 8460
rect 5760 8460 5778 8478
rect 5760 8478 5778 8496
rect 5760 8496 5778 8514
rect 5760 8514 5778 8532
rect 5760 8532 5778 8550
rect 5760 8550 5778 8568
rect 5760 8568 5778 8586
rect 5760 8586 5778 8604
rect 5760 8604 5778 8622
rect 5760 8622 5778 8640
rect 5760 8640 5778 8658
rect 5760 8658 5778 8676
rect 5760 8676 5778 8694
rect 5760 8694 5778 8712
rect 5760 8712 5778 8730
rect 5760 8730 5778 8748
rect 5760 8748 5778 8766
rect 5760 8766 5778 8784
rect 5760 8784 5778 8802
rect 5760 8802 5778 8820
rect 5760 8820 5778 8838
rect 5760 8838 5778 8856
rect 5760 8856 5778 8874
rect 5760 8874 5778 8892
rect 5760 8892 5778 8910
rect 5778 720 5796 738
rect 5778 738 5796 756
rect 5778 756 5796 774
rect 5778 774 5796 792
rect 5778 792 5796 810
rect 5778 810 5796 828
rect 5778 828 5796 846
rect 5778 846 5796 864
rect 5778 864 5796 882
rect 5778 882 5796 900
rect 5778 900 5796 918
rect 5778 918 5796 936
rect 5778 936 5796 954
rect 5778 954 5796 972
rect 5778 972 5796 990
rect 5778 990 5796 1008
rect 5778 1008 5796 1026
rect 5778 1170 5796 1188
rect 5778 1188 5796 1206
rect 5778 1206 5796 1224
rect 5778 1224 5796 1242
rect 5778 1242 5796 1260
rect 5778 1260 5796 1278
rect 5778 1278 5796 1296
rect 5778 1296 5796 1314
rect 5778 1314 5796 1332
rect 5778 1332 5796 1350
rect 5778 1350 5796 1368
rect 5778 1368 5796 1386
rect 5778 1386 5796 1404
rect 5778 1404 5796 1422
rect 5778 1422 5796 1440
rect 5778 1440 5796 1458
rect 5778 1458 5796 1476
rect 5778 1476 5796 1494
rect 5778 1494 5796 1512
rect 5778 1512 5796 1530
rect 5778 1530 5796 1548
rect 5778 1548 5796 1566
rect 5778 1566 5796 1584
rect 5778 1584 5796 1602
rect 5778 1602 5796 1620
rect 5778 1620 5796 1638
rect 5778 1638 5796 1656
rect 5778 1656 5796 1674
rect 5778 1674 5796 1692
rect 5778 1692 5796 1710
rect 5778 1710 5796 1728
rect 5778 1728 5796 1746
rect 5778 1746 5796 1764
rect 5778 1764 5796 1782
rect 5778 1782 5796 1800
rect 5778 1800 5796 1818
rect 5778 1818 5796 1836
rect 5778 1836 5796 1854
rect 5778 1854 5796 1872
rect 5778 1872 5796 1890
rect 5778 1890 5796 1908
rect 5778 1908 5796 1926
rect 5778 1926 5796 1944
rect 5778 1944 5796 1962
rect 5778 1962 5796 1980
rect 5778 1980 5796 1998
rect 5778 1998 5796 2016
rect 5778 2016 5796 2034
rect 5778 2034 5796 2052
rect 5778 2052 5796 2070
rect 5778 2070 5796 2088
rect 5778 2088 5796 2106
rect 5778 2106 5796 2124
rect 5778 2124 5796 2142
rect 5778 2142 5796 2160
rect 5778 2160 5796 2178
rect 5778 2178 5796 2196
rect 5778 2196 5796 2214
rect 5778 2214 5796 2232
rect 5778 2232 5796 2250
rect 5778 2250 5796 2268
rect 5778 2268 5796 2286
rect 5778 2286 5796 2304
rect 5778 2304 5796 2322
rect 5778 2322 5796 2340
rect 5778 2340 5796 2358
rect 5778 2358 5796 2376
rect 5778 2376 5796 2394
rect 5778 2394 5796 2412
rect 5778 2412 5796 2430
rect 5778 2430 5796 2448
rect 5778 2448 5796 2466
rect 5778 2466 5796 2484
rect 5778 2484 5796 2502
rect 5778 2502 5796 2520
rect 5778 2520 5796 2538
rect 5778 2538 5796 2556
rect 5778 2556 5796 2574
rect 5778 2574 5796 2592
rect 5778 2592 5796 2610
rect 5778 2610 5796 2628
rect 5778 2628 5796 2646
rect 5778 2880 5796 2898
rect 5778 2898 5796 2916
rect 5778 2916 5796 2934
rect 5778 2934 5796 2952
rect 5778 2952 5796 2970
rect 5778 2970 5796 2988
rect 5778 2988 5796 3006
rect 5778 3006 5796 3024
rect 5778 3024 5796 3042
rect 5778 3042 5796 3060
rect 5778 3060 5796 3078
rect 5778 3078 5796 3096
rect 5778 3096 5796 3114
rect 5778 3114 5796 3132
rect 5778 3132 5796 3150
rect 5778 3150 5796 3168
rect 5778 3168 5796 3186
rect 5778 3186 5796 3204
rect 5778 3204 5796 3222
rect 5778 3222 5796 3240
rect 5778 3240 5796 3258
rect 5778 3258 5796 3276
rect 5778 3276 5796 3294
rect 5778 3294 5796 3312
rect 5778 3312 5796 3330
rect 5778 3330 5796 3348
rect 5778 3348 5796 3366
rect 5778 3366 5796 3384
rect 5778 3384 5796 3402
rect 5778 3402 5796 3420
rect 5778 3420 5796 3438
rect 5778 3438 5796 3456
rect 5778 3456 5796 3474
rect 5778 3474 5796 3492
rect 5778 3492 5796 3510
rect 5778 3510 5796 3528
rect 5778 3528 5796 3546
rect 5778 3546 5796 3564
rect 5778 3564 5796 3582
rect 5778 3582 5796 3600
rect 5778 3600 5796 3618
rect 5778 3618 5796 3636
rect 5778 3636 5796 3654
rect 5778 3654 5796 3672
rect 5778 3672 5796 3690
rect 5778 3690 5796 3708
rect 5778 3708 5796 3726
rect 5778 3726 5796 3744
rect 5778 3744 5796 3762
rect 5778 3762 5796 3780
rect 5778 3780 5796 3798
rect 5778 3798 5796 3816
rect 5778 3816 5796 3834
rect 5778 3834 5796 3852
rect 5778 3852 5796 3870
rect 5778 3870 5796 3888
rect 5778 3888 5796 3906
rect 5778 3906 5796 3924
rect 5778 3924 5796 3942
rect 5778 3942 5796 3960
rect 5778 3960 5796 3978
rect 5778 3978 5796 3996
rect 5778 3996 5796 4014
rect 5778 4014 5796 4032
rect 5778 4032 5796 4050
rect 5778 4050 5796 4068
rect 5778 4068 5796 4086
rect 5778 4086 5796 4104
rect 5778 4104 5796 4122
rect 5778 4122 5796 4140
rect 5778 4140 5796 4158
rect 5778 4158 5796 4176
rect 5778 4176 5796 4194
rect 5778 4194 5796 4212
rect 5778 4212 5796 4230
rect 5778 4230 5796 4248
rect 5778 4248 5796 4266
rect 5778 4266 5796 4284
rect 5778 4284 5796 4302
rect 5778 4302 5796 4320
rect 5778 4320 5796 4338
rect 5778 4338 5796 4356
rect 5778 4356 5796 4374
rect 5778 4374 5796 4392
rect 5778 4392 5796 4410
rect 5778 4410 5796 4428
rect 5778 4428 5796 4446
rect 5778 4446 5796 4464
rect 5778 4464 5796 4482
rect 5778 4482 5796 4500
rect 5778 4500 5796 4518
rect 5778 4518 5796 4536
rect 5778 4536 5796 4554
rect 5778 4554 5796 4572
rect 5778 4572 5796 4590
rect 5778 4590 5796 4608
rect 5778 4608 5796 4626
rect 5778 4626 5796 4644
rect 5778 4644 5796 4662
rect 5778 4662 5796 4680
rect 5778 4680 5796 4698
rect 5778 4698 5796 4716
rect 5778 4716 5796 4734
rect 5778 4734 5796 4752
rect 5778 4752 5796 4770
rect 5778 4770 5796 4788
rect 5778 4788 5796 4806
rect 5778 4806 5796 4824
rect 5778 4824 5796 4842
rect 5778 4842 5796 4860
rect 5778 4860 5796 4878
rect 5778 4878 5796 4896
rect 5778 4896 5796 4914
rect 5778 4914 5796 4932
rect 5778 4932 5796 4950
rect 5778 4950 5796 4968
rect 5778 4968 5796 4986
rect 5778 4986 5796 5004
rect 5778 5004 5796 5022
rect 5778 5022 5796 5040
rect 5778 5040 5796 5058
rect 5778 5058 5796 5076
rect 5778 5076 5796 5094
rect 5778 5094 5796 5112
rect 5778 5112 5796 5130
rect 5778 5130 5796 5148
rect 5778 5148 5796 5166
rect 5778 5418 5796 5436
rect 5778 5436 5796 5454
rect 5778 5454 5796 5472
rect 5778 5472 5796 5490
rect 5778 5490 5796 5508
rect 5778 5508 5796 5526
rect 5778 5526 5796 5544
rect 5778 5544 5796 5562
rect 5778 5562 5796 5580
rect 5778 5580 5796 5598
rect 5778 5598 5796 5616
rect 5778 5616 5796 5634
rect 5778 5634 5796 5652
rect 5778 5652 5796 5670
rect 5778 5670 5796 5688
rect 5778 5688 5796 5706
rect 5778 5706 5796 5724
rect 5778 5724 5796 5742
rect 5778 5742 5796 5760
rect 5778 5760 5796 5778
rect 5778 5778 5796 5796
rect 5778 5796 5796 5814
rect 5778 5814 5796 5832
rect 5778 5832 5796 5850
rect 5778 5850 5796 5868
rect 5778 5868 5796 5886
rect 5778 5886 5796 5904
rect 5778 5904 5796 5922
rect 5778 5922 5796 5940
rect 5778 5940 5796 5958
rect 5778 5958 5796 5976
rect 5778 5976 5796 5994
rect 5778 5994 5796 6012
rect 5778 6012 5796 6030
rect 5778 6030 5796 6048
rect 5778 6048 5796 6066
rect 5778 6066 5796 6084
rect 5778 6084 5796 6102
rect 5778 6102 5796 6120
rect 5778 6120 5796 6138
rect 5778 6138 5796 6156
rect 5778 6156 5796 6174
rect 5778 6174 5796 6192
rect 5778 6192 5796 6210
rect 5778 6210 5796 6228
rect 5778 6228 5796 6246
rect 5778 6246 5796 6264
rect 5778 6264 5796 6282
rect 5778 6282 5796 6300
rect 5778 6300 5796 6318
rect 5778 6318 5796 6336
rect 5778 6336 5796 6354
rect 5778 6354 5796 6372
rect 5778 6372 5796 6390
rect 5778 6390 5796 6408
rect 5778 6408 5796 6426
rect 5778 6426 5796 6444
rect 5778 6444 5796 6462
rect 5778 6462 5796 6480
rect 5778 6480 5796 6498
rect 5778 6498 5796 6516
rect 5778 6516 5796 6534
rect 5778 6534 5796 6552
rect 5778 6552 5796 6570
rect 5778 6570 5796 6588
rect 5778 6588 5796 6606
rect 5778 6606 5796 6624
rect 5778 6624 5796 6642
rect 5778 6642 5796 6660
rect 5778 6660 5796 6678
rect 5778 6678 5796 6696
rect 5778 6696 5796 6714
rect 5778 6714 5796 6732
rect 5778 6732 5796 6750
rect 5778 6750 5796 6768
rect 5778 6768 5796 6786
rect 5778 6786 5796 6804
rect 5778 6804 5796 6822
rect 5778 6822 5796 6840
rect 5778 6840 5796 6858
rect 5778 6858 5796 6876
rect 5778 6876 5796 6894
rect 5778 6894 5796 6912
rect 5778 6912 5796 6930
rect 5778 6930 5796 6948
rect 5778 6948 5796 6966
rect 5778 6966 5796 6984
rect 5778 6984 5796 7002
rect 5778 7002 5796 7020
rect 5778 7020 5796 7038
rect 5778 7038 5796 7056
rect 5778 7056 5796 7074
rect 5778 7074 5796 7092
rect 5778 7092 5796 7110
rect 5778 7110 5796 7128
rect 5778 7128 5796 7146
rect 5778 7146 5796 7164
rect 5778 7164 5796 7182
rect 5778 7182 5796 7200
rect 5778 7200 5796 7218
rect 5778 7218 5796 7236
rect 5778 7236 5796 7254
rect 5778 7254 5796 7272
rect 5778 7272 5796 7290
rect 5778 7290 5796 7308
rect 5778 7308 5796 7326
rect 5778 7326 5796 7344
rect 5778 7344 5796 7362
rect 5778 7362 5796 7380
rect 5778 7380 5796 7398
rect 5778 7398 5796 7416
rect 5778 7416 5796 7434
rect 5778 7434 5796 7452
rect 5778 7452 5796 7470
rect 5778 7470 5796 7488
rect 5778 7488 5796 7506
rect 5778 7506 5796 7524
rect 5778 7524 5796 7542
rect 5778 7542 5796 7560
rect 5778 7560 5796 7578
rect 5778 7578 5796 7596
rect 5778 7596 5796 7614
rect 5778 7614 5796 7632
rect 5778 7632 5796 7650
rect 5778 7650 5796 7668
rect 5778 7668 5796 7686
rect 5778 7686 5796 7704
rect 5778 7704 5796 7722
rect 5778 7722 5796 7740
rect 5778 7740 5796 7758
rect 5778 7758 5796 7776
rect 5778 7776 5796 7794
rect 5778 7794 5796 7812
rect 5778 7812 5796 7830
rect 5778 7830 5796 7848
rect 5778 7848 5796 7866
rect 5778 7866 5796 7884
rect 5778 7884 5796 7902
rect 5778 7902 5796 7920
rect 5778 7920 5796 7938
rect 5778 7938 5796 7956
rect 5778 7956 5796 7974
rect 5778 7974 5796 7992
rect 5778 7992 5796 8010
rect 5778 8010 5796 8028
rect 5778 8028 5796 8046
rect 5778 8046 5796 8064
rect 5778 8064 5796 8082
rect 5778 8082 5796 8100
rect 5778 8100 5796 8118
rect 5778 8118 5796 8136
rect 5778 8136 5796 8154
rect 5778 8154 5796 8172
rect 5778 8172 5796 8190
rect 5778 8190 5796 8208
rect 5778 8208 5796 8226
rect 5778 8226 5796 8244
rect 5778 8244 5796 8262
rect 5778 8262 5796 8280
rect 5778 8280 5796 8298
rect 5778 8298 5796 8316
rect 5778 8316 5796 8334
rect 5778 8334 5796 8352
rect 5778 8352 5796 8370
rect 5778 8370 5796 8388
rect 5778 8388 5796 8406
rect 5778 8406 5796 8424
rect 5778 8424 5796 8442
rect 5778 8442 5796 8460
rect 5778 8460 5796 8478
rect 5778 8478 5796 8496
rect 5778 8496 5796 8514
rect 5778 8514 5796 8532
rect 5778 8532 5796 8550
rect 5778 8550 5796 8568
rect 5778 8568 5796 8586
rect 5778 8586 5796 8604
rect 5778 8604 5796 8622
rect 5778 8622 5796 8640
rect 5778 8640 5796 8658
rect 5778 8658 5796 8676
rect 5778 8676 5796 8694
rect 5778 8694 5796 8712
rect 5778 8712 5796 8730
rect 5778 8730 5796 8748
rect 5778 8748 5796 8766
rect 5778 8766 5796 8784
rect 5778 8784 5796 8802
rect 5778 8802 5796 8820
rect 5778 8820 5796 8838
rect 5778 8838 5796 8856
rect 5778 8856 5796 8874
rect 5778 8874 5796 8892
rect 5778 8892 5796 8910
rect 5778 8910 5796 8928
rect 5778 8928 5796 8946
rect 5796 738 5814 756
rect 5796 756 5814 774
rect 5796 774 5814 792
rect 5796 792 5814 810
rect 5796 810 5814 828
rect 5796 828 5814 846
rect 5796 846 5814 864
rect 5796 864 5814 882
rect 5796 882 5814 900
rect 5796 900 5814 918
rect 5796 918 5814 936
rect 5796 936 5814 954
rect 5796 954 5814 972
rect 5796 972 5814 990
rect 5796 990 5814 1008
rect 5796 1008 5814 1026
rect 5796 1170 5814 1188
rect 5796 1188 5814 1206
rect 5796 1206 5814 1224
rect 5796 1224 5814 1242
rect 5796 1242 5814 1260
rect 5796 1260 5814 1278
rect 5796 1278 5814 1296
rect 5796 1296 5814 1314
rect 5796 1314 5814 1332
rect 5796 1332 5814 1350
rect 5796 1350 5814 1368
rect 5796 1368 5814 1386
rect 5796 1386 5814 1404
rect 5796 1404 5814 1422
rect 5796 1422 5814 1440
rect 5796 1440 5814 1458
rect 5796 1458 5814 1476
rect 5796 1476 5814 1494
rect 5796 1494 5814 1512
rect 5796 1512 5814 1530
rect 5796 1530 5814 1548
rect 5796 1548 5814 1566
rect 5796 1566 5814 1584
rect 5796 1584 5814 1602
rect 5796 1602 5814 1620
rect 5796 1620 5814 1638
rect 5796 1638 5814 1656
rect 5796 1656 5814 1674
rect 5796 1674 5814 1692
rect 5796 1692 5814 1710
rect 5796 1710 5814 1728
rect 5796 1728 5814 1746
rect 5796 1746 5814 1764
rect 5796 1764 5814 1782
rect 5796 1782 5814 1800
rect 5796 1800 5814 1818
rect 5796 1818 5814 1836
rect 5796 1836 5814 1854
rect 5796 1854 5814 1872
rect 5796 1872 5814 1890
rect 5796 1890 5814 1908
rect 5796 1908 5814 1926
rect 5796 1926 5814 1944
rect 5796 1944 5814 1962
rect 5796 1962 5814 1980
rect 5796 1980 5814 1998
rect 5796 1998 5814 2016
rect 5796 2016 5814 2034
rect 5796 2034 5814 2052
rect 5796 2052 5814 2070
rect 5796 2070 5814 2088
rect 5796 2088 5814 2106
rect 5796 2106 5814 2124
rect 5796 2124 5814 2142
rect 5796 2142 5814 2160
rect 5796 2160 5814 2178
rect 5796 2178 5814 2196
rect 5796 2196 5814 2214
rect 5796 2214 5814 2232
rect 5796 2232 5814 2250
rect 5796 2250 5814 2268
rect 5796 2268 5814 2286
rect 5796 2286 5814 2304
rect 5796 2304 5814 2322
rect 5796 2322 5814 2340
rect 5796 2340 5814 2358
rect 5796 2358 5814 2376
rect 5796 2376 5814 2394
rect 5796 2394 5814 2412
rect 5796 2412 5814 2430
rect 5796 2430 5814 2448
rect 5796 2448 5814 2466
rect 5796 2466 5814 2484
rect 5796 2484 5814 2502
rect 5796 2502 5814 2520
rect 5796 2520 5814 2538
rect 5796 2538 5814 2556
rect 5796 2556 5814 2574
rect 5796 2574 5814 2592
rect 5796 2592 5814 2610
rect 5796 2610 5814 2628
rect 5796 2628 5814 2646
rect 5796 2646 5814 2664
rect 5796 2880 5814 2898
rect 5796 2898 5814 2916
rect 5796 2916 5814 2934
rect 5796 2934 5814 2952
rect 5796 2952 5814 2970
rect 5796 2970 5814 2988
rect 5796 2988 5814 3006
rect 5796 3006 5814 3024
rect 5796 3024 5814 3042
rect 5796 3042 5814 3060
rect 5796 3060 5814 3078
rect 5796 3078 5814 3096
rect 5796 3096 5814 3114
rect 5796 3114 5814 3132
rect 5796 3132 5814 3150
rect 5796 3150 5814 3168
rect 5796 3168 5814 3186
rect 5796 3186 5814 3204
rect 5796 3204 5814 3222
rect 5796 3222 5814 3240
rect 5796 3240 5814 3258
rect 5796 3258 5814 3276
rect 5796 3276 5814 3294
rect 5796 3294 5814 3312
rect 5796 3312 5814 3330
rect 5796 3330 5814 3348
rect 5796 3348 5814 3366
rect 5796 3366 5814 3384
rect 5796 3384 5814 3402
rect 5796 3402 5814 3420
rect 5796 3420 5814 3438
rect 5796 3438 5814 3456
rect 5796 3456 5814 3474
rect 5796 3474 5814 3492
rect 5796 3492 5814 3510
rect 5796 3510 5814 3528
rect 5796 3528 5814 3546
rect 5796 3546 5814 3564
rect 5796 3564 5814 3582
rect 5796 3582 5814 3600
rect 5796 3600 5814 3618
rect 5796 3618 5814 3636
rect 5796 3636 5814 3654
rect 5796 3654 5814 3672
rect 5796 3672 5814 3690
rect 5796 3690 5814 3708
rect 5796 3708 5814 3726
rect 5796 3726 5814 3744
rect 5796 3744 5814 3762
rect 5796 3762 5814 3780
rect 5796 3780 5814 3798
rect 5796 3798 5814 3816
rect 5796 3816 5814 3834
rect 5796 3834 5814 3852
rect 5796 3852 5814 3870
rect 5796 3870 5814 3888
rect 5796 3888 5814 3906
rect 5796 3906 5814 3924
rect 5796 3924 5814 3942
rect 5796 3942 5814 3960
rect 5796 3960 5814 3978
rect 5796 3978 5814 3996
rect 5796 3996 5814 4014
rect 5796 4014 5814 4032
rect 5796 4032 5814 4050
rect 5796 4050 5814 4068
rect 5796 4068 5814 4086
rect 5796 4086 5814 4104
rect 5796 4104 5814 4122
rect 5796 4122 5814 4140
rect 5796 4140 5814 4158
rect 5796 4158 5814 4176
rect 5796 4176 5814 4194
rect 5796 4194 5814 4212
rect 5796 4212 5814 4230
rect 5796 4230 5814 4248
rect 5796 4248 5814 4266
rect 5796 4266 5814 4284
rect 5796 4284 5814 4302
rect 5796 4302 5814 4320
rect 5796 4320 5814 4338
rect 5796 4338 5814 4356
rect 5796 4356 5814 4374
rect 5796 4374 5814 4392
rect 5796 4392 5814 4410
rect 5796 4410 5814 4428
rect 5796 4428 5814 4446
rect 5796 4446 5814 4464
rect 5796 4464 5814 4482
rect 5796 4482 5814 4500
rect 5796 4500 5814 4518
rect 5796 4518 5814 4536
rect 5796 4536 5814 4554
rect 5796 4554 5814 4572
rect 5796 4572 5814 4590
rect 5796 4590 5814 4608
rect 5796 4608 5814 4626
rect 5796 4626 5814 4644
rect 5796 4644 5814 4662
rect 5796 4662 5814 4680
rect 5796 4680 5814 4698
rect 5796 4698 5814 4716
rect 5796 4716 5814 4734
rect 5796 4734 5814 4752
rect 5796 4752 5814 4770
rect 5796 4770 5814 4788
rect 5796 4788 5814 4806
rect 5796 4806 5814 4824
rect 5796 4824 5814 4842
rect 5796 4842 5814 4860
rect 5796 4860 5814 4878
rect 5796 4878 5814 4896
rect 5796 4896 5814 4914
rect 5796 4914 5814 4932
rect 5796 4932 5814 4950
rect 5796 4950 5814 4968
rect 5796 4968 5814 4986
rect 5796 4986 5814 5004
rect 5796 5004 5814 5022
rect 5796 5022 5814 5040
rect 5796 5040 5814 5058
rect 5796 5058 5814 5076
rect 5796 5076 5814 5094
rect 5796 5094 5814 5112
rect 5796 5112 5814 5130
rect 5796 5130 5814 5148
rect 5796 5148 5814 5166
rect 5796 5166 5814 5184
rect 5796 5436 5814 5454
rect 5796 5454 5814 5472
rect 5796 5472 5814 5490
rect 5796 5490 5814 5508
rect 5796 5508 5814 5526
rect 5796 5526 5814 5544
rect 5796 5544 5814 5562
rect 5796 5562 5814 5580
rect 5796 5580 5814 5598
rect 5796 5598 5814 5616
rect 5796 5616 5814 5634
rect 5796 5634 5814 5652
rect 5796 5652 5814 5670
rect 5796 5670 5814 5688
rect 5796 5688 5814 5706
rect 5796 5706 5814 5724
rect 5796 5724 5814 5742
rect 5796 5742 5814 5760
rect 5796 5760 5814 5778
rect 5796 5778 5814 5796
rect 5796 5796 5814 5814
rect 5796 5814 5814 5832
rect 5796 5832 5814 5850
rect 5796 5850 5814 5868
rect 5796 5868 5814 5886
rect 5796 5886 5814 5904
rect 5796 5904 5814 5922
rect 5796 5922 5814 5940
rect 5796 5940 5814 5958
rect 5796 5958 5814 5976
rect 5796 5976 5814 5994
rect 5796 5994 5814 6012
rect 5796 6012 5814 6030
rect 5796 6030 5814 6048
rect 5796 6048 5814 6066
rect 5796 6066 5814 6084
rect 5796 6084 5814 6102
rect 5796 6102 5814 6120
rect 5796 6120 5814 6138
rect 5796 6138 5814 6156
rect 5796 6156 5814 6174
rect 5796 6174 5814 6192
rect 5796 6192 5814 6210
rect 5796 6210 5814 6228
rect 5796 6228 5814 6246
rect 5796 6246 5814 6264
rect 5796 6264 5814 6282
rect 5796 6282 5814 6300
rect 5796 6300 5814 6318
rect 5796 6318 5814 6336
rect 5796 6336 5814 6354
rect 5796 6354 5814 6372
rect 5796 6372 5814 6390
rect 5796 6390 5814 6408
rect 5796 6408 5814 6426
rect 5796 6426 5814 6444
rect 5796 6444 5814 6462
rect 5796 6462 5814 6480
rect 5796 6480 5814 6498
rect 5796 6498 5814 6516
rect 5796 6516 5814 6534
rect 5796 6534 5814 6552
rect 5796 6552 5814 6570
rect 5796 6570 5814 6588
rect 5796 6588 5814 6606
rect 5796 6606 5814 6624
rect 5796 6624 5814 6642
rect 5796 6642 5814 6660
rect 5796 6660 5814 6678
rect 5796 6678 5814 6696
rect 5796 6696 5814 6714
rect 5796 6714 5814 6732
rect 5796 6732 5814 6750
rect 5796 6750 5814 6768
rect 5796 6768 5814 6786
rect 5796 6786 5814 6804
rect 5796 6804 5814 6822
rect 5796 6822 5814 6840
rect 5796 6840 5814 6858
rect 5796 6858 5814 6876
rect 5796 6876 5814 6894
rect 5796 6894 5814 6912
rect 5796 6912 5814 6930
rect 5796 6930 5814 6948
rect 5796 6948 5814 6966
rect 5796 6966 5814 6984
rect 5796 6984 5814 7002
rect 5796 7002 5814 7020
rect 5796 7020 5814 7038
rect 5796 7038 5814 7056
rect 5796 7056 5814 7074
rect 5796 7074 5814 7092
rect 5796 7092 5814 7110
rect 5796 7110 5814 7128
rect 5796 7128 5814 7146
rect 5796 7146 5814 7164
rect 5796 7164 5814 7182
rect 5796 7182 5814 7200
rect 5796 7200 5814 7218
rect 5796 7218 5814 7236
rect 5796 7236 5814 7254
rect 5796 7254 5814 7272
rect 5796 7272 5814 7290
rect 5796 7290 5814 7308
rect 5796 7308 5814 7326
rect 5796 7326 5814 7344
rect 5796 7344 5814 7362
rect 5796 7362 5814 7380
rect 5796 7380 5814 7398
rect 5796 7398 5814 7416
rect 5796 7416 5814 7434
rect 5796 7434 5814 7452
rect 5796 7452 5814 7470
rect 5796 7470 5814 7488
rect 5796 7488 5814 7506
rect 5796 7506 5814 7524
rect 5796 7524 5814 7542
rect 5796 7542 5814 7560
rect 5796 7560 5814 7578
rect 5796 7578 5814 7596
rect 5796 7596 5814 7614
rect 5796 7614 5814 7632
rect 5796 7632 5814 7650
rect 5796 7650 5814 7668
rect 5796 7668 5814 7686
rect 5796 7686 5814 7704
rect 5796 7704 5814 7722
rect 5796 7722 5814 7740
rect 5796 7740 5814 7758
rect 5796 7758 5814 7776
rect 5796 7776 5814 7794
rect 5796 7794 5814 7812
rect 5796 7812 5814 7830
rect 5796 7830 5814 7848
rect 5796 7848 5814 7866
rect 5796 7866 5814 7884
rect 5796 7884 5814 7902
rect 5796 7902 5814 7920
rect 5796 7920 5814 7938
rect 5796 7938 5814 7956
rect 5796 7956 5814 7974
rect 5796 7974 5814 7992
rect 5796 7992 5814 8010
rect 5796 8010 5814 8028
rect 5796 8028 5814 8046
rect 5796 8046 5814 8064
rect 5796 8064 5814 8082
rect 5796 8082 5814 8100
rect 5796 8100 5814 8118
rect 5796 8118 5814 8136
rect 5796 8136 5814 8154
rect 5796 8154 5814 8172
rect 5796 8172 5814 8190
rect 5796 8190 5814 8208
rect 5796 8208 5814 8226
rect 5796 8226 5814 8244
rect 5796 8244 5814 8262
rect 5796 8262 5814 8280
rect 5796 8280 5814 8298
rect 5796 8298 5814 8316
rect 5796 8316 5814 8334
rect 5796 8334 5814 8352
rect 5796 8352 5814 8370
rect 5796 8370 5814 8388
rect 5796 8388 5814 8406
rect 5796 8406 5814 8424
rect 5796 8424 5814 8442
rect 5796 8442 5814 8460
rect 5796 8460 5814 8478
rect 5796 8478 5814 8496
rect 5796 8496 5814 8514
rect 5796 8514 5814 8532
rect 5796 8532 5814 8550
rect 5796 8550 5814 8568
rect 5796 8568 5814 8586
rect 5796 8586 5814 8604
rect 5796 8604 5814 8622
rect 5796 8622 5814 8640
rect 5796 8640 5814 8658
rect 5796 8658 5814 8676
rect 5796 8676 5814 8694
rect 5796 8694 5814 8712
rect 5796 8712 5814 8730
rect 5796 8730 5814 8748
rect 5796 8748 5814 8766
rect 5796 8766 5814 8784
rect 5796 8784 5814 8802
rect 5796 8802 5814 8820
rect 5796 8820 5814 8838
rect 5796 8838 5814 8856
rect 5796 8856 5814 8874
rect 5796 8874 5814 8892
rect 5796 8892 5814 8910
rect 5796 8910 5814 8928
rect 5796 8928 5814 8946
rect 5796 8946 5814 8964
rect 5814 756 5832 774
rect 5814 774 5832 792
rect 5814 792 5832 810
rect 5814 810 5832 828
rect 5814 828 5832 846
rect 5814 846 5832 864
rect 5814 864 5832 882
rect 5814 882 5832 900
rect 5814 900 5832 918
rect 5814 918 5832 936
rect 5814 936 5832 954
rect 5814 954 5832 972
rect 5814 972 5832 990
rect 5814 990 5832 1008
rect 5814 1008 5832 1026
rect 5814 1026 5832 1044
rect 5814 1188 5832 1206
rect 5814 1206 5832 1224
rect 5814 1224 5832 1242
rect 5814 1242 5832 1260
rect 5814 1260 5832 1278
rect 5814 1278 5832 1296
rect 5814 1296 5832 1314
rect 5814 1314 5832 1332
rect 5814 1332 5832 1350
rect 5814 1350 5832 1368
rect 5814 1368 5832 1386
rect 5814 1386 5832 1404
rect 5814 1404 5832 1422
rect 5814 1422 5832 1440
rect 5814 1440 5832 1458
rect 5814 1458 5832 1476
rect 5814 1476 5832 1494
rect 5814 1494 5832 1512
rect 5814 1512 5832 1530
rect 5814 1530 5832 1548
rect 5814 1548 5832 1566
rect 5814 1566 5832 1584
rect 5814 1584 5832 1602
rect 5814 1602 5832 1620
rect 5814 1620 5832 1638
rect 5814 1638 5832 1656
rect 5814 1656 5832 1674
rect 5814 1674 5832 1692
rect 5814 1692 5832 1710
rect 5814 1710 5832 1728
rect 5814 1728 5832 1746
rect 5814 1746 5832 1764
rect 5814 1764 5832 1782
rect 5814 1782 5832 1800
rect 5814 1800 5832 1818
rect 5814 1818 5832 1836
rect 5814 1836 5832 1854
rect 5814 1854 5832 1872
rect 5814 1872 5832 1890
rect 5814 1890 5832 1908
rect 5814 1908 5832 1926
rect 5814 1926 5832 1944
rect 5814 1944 5832 1962
rect 5814 1962 5832 1980
rect 5814 1980 5832 1998
rect 5814 1998 5832 2016
rect 5814 2016 5832 2034
rect 5814 2034 5832 2052
rect 5814 2052 5832 2070
rect 5814 2070 5832 2088
rect 5814 2088 5832 2106
rect 5814 2106 5832 2124
rect 5814 2124 5832 2142
rect 5814 2142 5832 2160
rect 5814 2160 5832 2178
rect 5814 2178 5832 2196
rect 5814 2196 5832 2214
rect 5814 2214 5832 2232
rect 5814 2232 5832 2250
rect 5814 2250 5832 2268
rect 5814 2268 5832 2286
rect 5814 2286 5832 2304
rect 5814 2304 5832 2322
rect 5814 2322 5832 2340
rect 5814 2340 5832 2358
rect 5814 2358 5832 2376
rect 5814 2376 5832 2394
rect 5814 2394 5832 2412
rect 5814 2412 5832 2430
rect 5814 2430 5832 2448
rect 5814 2448 5832 2466
rect 5814 2466 5832 2484
rect 5814 2484 5832 2502
rect 5814 2502 5832 2520
rect 5814 2520 5832 2538
rect 5814 2538 5832 2556
rect 5814 2556 5832 2574
rect 5814 2574 5832 2592
rect 5814 2592 5832 2610
rect 5814 2610 5832 2628
rect 5814 2628 5832 2646
rect 5814 2646 5832 2664
rect 5814 2898 5832 2916
rect 5814 2916 5832 2934
rect 5814 2934 5832 2952
rect 5814 2952 5832 2970
rect 5814 2970 5832 2988
rect 5814 2988 5832 3006
rect 5814 3006 5832 3024
rect 5814 3024 5832 3042
rect 5814 3042 5832 3060
rect 5814 3060 5832 3078
rect 5814 3078 5832 3096
rect 5814 3096 5832 3114
rect 5814 3114 5832 3132
rect 5814 3132 5832 3150
rect 5814 3150 5832 3168
rect 5814 3168 5832 3186
rect 5814 3186 5832 3204
rect 5814 3204 5832 3222
rect 5814 3222 5832 3240
rect 5814 3240 5832 3258
rect 5814 3258 5832 3276
rect 5814 3276 5832 3294
rect 5814 3294 5832 3312
rect 5814 3312 5832 3330
rect 5814 3330 5832 3348
rect 5814 3348 5832 3366
rect 5814 3366 5832 3384
rect 5814 3384 5832 3402
rect 5814 3402 5832 3420
rect 5814 3420 5832 3438
rect 5814 3438 5832 3456
rect 5814 3456 5832 3474
rect 5814 3474 5832 3492
rect 5814 3492 5832 3510
rect 5814 3510 5832 3528
rect 5814 3528 5832 3546
rect 5814 3546 5832 3564
rect 5814 3564 5832 3582
rect 5814 3582 5832 3600
rect 5814 3600 5832 3618
rect 5814 3618 5832 3636
rect 5814 3636 5832 3654
rect 5814 3654 5832 3672
rect 5814 3672 5832 3690
rect 5814 3690 5832 3708
rect 5814 3708 5832 3726
rect 5814 3726 5832 3744
rect 5814 3744 5832 3762
rect 5814 3762 5832 3780
rect 5814 3780 5832 3798
rect 5814 3798 5832 3816
rect 5814 3816 5832 3834
rect 5814 3834 5832 3852
rect 5814 3852 5832 3870
rect 5814 3870 5832 3888
rect 5814 3888 5832 3906
rect 5814 3906 5832 3924
rect 5814 3924 5832 3942
rect 5814 3942 5832 3960
rect 5814 3960 5832 3978
rect 5814 3978 5832 3996
rect 5814 3996 5832 4014
rect 5814 4014 5832 4032
rect 5814 4032 5832 4050
rect 5814 4050 5832 4068
rect 5814 4068 5832 4086
rect 5814 4086 5832 4104
rect 5814 4104 5832 4122
rect 5814 4122 5832 4140
rect 5814 4140 5832 4158
rect 5814 4158 5832 4176
rect 5814 4176 5832 4194
rect 5814 4194 5832 4212
rect 5814 4212 5832 4230
rect 5814 4230 5832 4248
rect 5814 4248 5832 4266
rect 5814 4266 5832 4284
rect 5814 4284 5832 4302
rect 5814 4302 5832 4320
rect 5814 4320 5832 4338
rect 5814 4338 5832 4356
rect 5814 4356 5832 4374
rect 5814 4374 5832 4392
rect 5814 4392 5832 4410
rect 5814 4410 5832 4428
rect 5814 4428 5832 4446
rect 5814 4446 5832 4464
rect 5814 4464 5832 4482
rect 5814 4482 5832 4500
rect 5814 4500 5832 4518
rect 5814 4518 5832 4536
rect 5814 4536 5832 4554
rect 5814 4554 5832 4572
rect 5814 4572 5832 4590
rect 5814 4590 5832 4608
rect 5814 4608 5832 4626
rect 5814 4626 5832 4644
rect 5814 4644 5832 4662
rect 5814 4662 5832 4680
rect 5814 4680 5832 4698
rect 5814 4698 5832 4716
rect 5814 4716 5832 4734
rect 5814 4734 5832 4752
rect 5814 4752 5832 4770
rect 5814 4770 5832 4788
rect 5814 4788 5832 4806
rect 5814 4806 5832 4824
rect 5814 4824 5832 4842
rect 5814 4842 5832 4860
rect 5814 4860 5832 4878
rect 5814 4878 5832 4896
rect 5814 4896 5832 4914
rect 5814 4914 5832 4932
rect 5814 4932 5832 4950
rect 5814 4950 5832 4968
rect 5814 4968 5832 4986
rect 5814 4986 5832 5004
rect 5814 5004 5832 5022
rect 5814 5022 5832 5040
rect 5814 5040 5832 5058
rect 5814 5058 5832 5076
rect 5814 5076 5832 5094
rect 5814 5094 5832 5112
rect 5814 5112 5832 5130
rect 5814 5130 5832 5148
rect 5814 5148 5832 5166
rect 5814 5166 5832 5184
rect 5814 5184 5832 5202
rect 5814 5454 5832 5472
rect 5814 5472 5832 5490
rect 5814 5490 5832 5508
rect 5814 5508 5832 5526
rect 5814 5526 5832 5544
rect 5814 5544 5832 5562
rect 5814 5562 5832 5580
rect 5814 5580 5832 5598
rect 5814 5598 5832 5616
rect 5814 5616 5832 5634
rect 5814 5634 5832 5652
rect 5814 5652 5832 5670
rect 5814 5670 5832 5688
rect 5814 5688 5832 5706
rect 5814 5706 5832 5724
rect 5814 5724 5832 5742
rect 5814 5742 5832 5760
rect 5814 5760 5832 5778
rect 5814 5778 5832 5796
rect 5814 5796 5832 5814
rect 5814 5814 5832 5832
rect 5814 5832 5832 5850
rect 5814 5850 5832 5868
rect 5814 5868 5832 5886
rect 5814 5886 5832 5904
rect 5814 5904 5832 5922
rect 5814 5922 5832 5940
rect 5814 5940 5832 5958
rect 5814 5958 5832 5976
rect 5814 5976 5832 5994
rect 5814 5994 5832 6012
rect 5814 6012 5832 6030
rect 5814 6030 5832 6048
rect 5814 6048 5832 6066
rect 5814 6066 5832 6084
rect 5814 6084 5832 6102
rect 5814 6102 5832 6120
rect 5814 6120 5832 6138
rect 5814 6138 5832 6156
rect 5814 6156 5832 6174
rect 5814 6174 5832 6192
rect 5814 6192 5832 6210
rect 5814 6210 5832 6228
rect 5814 6228 5832 6246
rect 5814 6246 5832 6264
rect 5814 6264 5832 6282
rect 5814 6282 5832 6300
rect 5814 6300 5832 6318
rect 5814 6318 5832 6336
rect 5814 6336 5832 6354
rect 5814 6354 5832 6372
rect 5814 6372 5832 6390
rect 5814 6390 5832 6408
rect 5814 6408 5832 6426
rect 5814 6426 5832 6444
rect 5814 6444 5832 6462
rect 5814 6462 5832 6480
rect 5814 6480 5832 6498
rect 5814 6498 5832 6516
rect 5814 6516 5832 6534
rect 5814 6534 5832 6552
rect 5814 6552 5832 6570
rect 5814 6570 5832 6588
rect 5814 6588 5832 6606
rect 5814 6606 5832 6624
rect 5814 6624 5832 6642
rect 5814 6642 5832 6660
rect 5814 6660 5832 6678
rect 5814 6678 5832 6696
rect 5814 6696 5832 6714
rect 5814 6714 5832 6732
rect 5814 6732 5832 6750
rect 5814 6750 5832 6768
rect 5814 6768 5832 6786
rect 5814 6786 5832 6804
rect 5814 6804 5832 6822
rect 5814 6822 5832 6840
rect 5814 6840 5832 6858
rect 5814 6858 5832 6876
rect 5814 6876 5832 6894
rect 5814 6894 5832 6912
rect 5814 6912 5832 6930
rect 5814 6930 5832 6948
rect 5814 6948 5832 6966
rect 5814 6966 5832 6984
rect 5814 6984 5832 7002
rect 5814 7002 5832 7020
rect 5814 7020 5832 7038
rect 5814 7038 5832 7056
rect 5814 7056 5832 7074
rect 5814 7074 5832 7092
rect 5814 7092 5832 7110
rect 5814 7110 5832 7128
rect 5814 7128 5832 7146
rect 5814 7146 5832 7164
rect 5814 7164 5832 7182
rect 5814 7182 5832 7200
rect 5814 7200 5832 7218
rect 5814 7218 5832 7236
rect 5814 7236 5832 7254
rect 5814 7254 5832 7272
rect 5814 7272 5832 7290
rect 5814 7290 5832 7308
rect 5814 7308 5832 7326
rect 5814 7326 5832 7344
rect 5814 7344 5832 7362
rect 5814 7362 5832 7380
rect 5814 7380 5832 7398
rect 5814 7398 5832 7416
rect 5814 7416 5832 7434
rect 5814 7434 5832 7452
rect 5814 7452 5832 7470
rect 5814 7470 5832 7488
rect 5814 7488 5832 7506
rect 5814 7506 5832 7524
rect 5814 7524 5832 7542
rect 5814 7542 5832 7560
rect 5814 7560 5832 7578
rect 5814 7578 5832 7596
rect 5814 7596 5832 7614
rect 5814 7614 5832 7632
rect 5814 7632 5832 7650
rect 5814 7650 5832 7668
rect 5814 7668 5832 7686
rect 5814 7686 5832 7704
rect 5814 7704 5832 7722
rect 5814 7722 5832 7740
rect 5814 7740 5832 7758
rect 5814 7758 5832 7776
rect 5814 7776 5832 7794
rect 5814 7794 5832 7812
rect 5814 7812 5832 7830
rect 5814 7830 5832 7848
rect 5814 7848 5832 7866
rect 5814 7866 5832 7884
rect 5814 7884 5832 7902
rect 5814 7902 5832 7920
rect 5814 7920 5832 7938
rect 5814 7938 5832 7956
rect 5814 7956 5832 7974
rect 5814 7974 5832 7992
rect 5814 7992 5832 8010
rect 5814 8010 5832 8028
rect 5814 8028 5832 8046
rect 5814 8046 5832 8064
rect 5814 8064 5832 8082
rect 5814 8082 5832 8100
rect 5814 8100 5832 8118
rect 5814 8118 5832 8136
rect 5814 8136 5832 8154
rect 5814 8154 5832 8172
rect 5814 8172 5832 8190
rect 5814 8190 5832 8208
rect 5814 8208 5832 8226
rect 5814 8226 5832 8244
rect 5814 8244 5832 8262
rect 5814 8262 5832 8280
rect 5814 8280 5832 8298
rect 5814 8298 5832 8316
rect 5814 8316 5832 8334
rect 5814 8334 5832 8352
rect 5814 8352 5832 8370
rect 5814 8370 5832 8388
rect 5814 8388 5832 8406
rect 5814 8406 5832 8424
rect 5814 8424 5832 8442
rect 5814 8442 5832 8460
rect 5814 8460 5832 8478
rect 5814 8478 5832 8496
rect 5814 8496 5832 8514
rect 5814 8514 5832 8532
rect 5814 8532 5832 8550
rect 5814 8550 5832 8568
rect 5814 8568 5832 8586
rect 5814 8586 5832 8604
rect 5814 8604 5832 8622
rect 5814 8622 5832 8640
rect 5814 8640 5832 8658
rect 5814 8658 5832 8676
rect 5814 8676 5832 8694
rect 5814 8694 5832 8712
rect 5814 8712 5832 8730
rect 5814 8730 5832 8748
rect 5814 8748 5832 8766
rect 5814 8766 5832 8784
rect 5814 8784 5832 8802
rect 5814 8802 5832 8820
rect 5814 8820 5832 8838
rect 5814 8838 5832 8856
rect 5814 8856 5832 8874
rect 5814 8874 5832 8892
rect 5814 8892 5832 8910
rect 5814 8910 5832 8928
rect 5814 8928 5832 8946
rect 5814 8946 5832 8964
rect 5814 8964 5832 8982
rect 5832 756 5850 774
rect 5832 774 5850 792
rect 5832 792 5850 810
rect 5832 810 5850 828
rect 5832 828 5850 846
rect 5832 846 5850 864
rect 5832 864 5850 882
rect 5832 882 5850 900
rect 5832 900 5850 918
rect 5832 918 5850 936
rect 5832 936 5850 954
rect 5832 954 5850 972
rect 5832 972 5850 990
rect 5832 990 5850 1008
rect 5832 1008 5850 1026
rect 5832 1026 5850 1044
rect 5832 1188 5850 1206
rect 5832 1206 5850 1224
rect 5832 1224 5850 1242
rect 5832 1242 5850 1260
rect 5832 1260 5850 1278
rect 5832 1278 5850 1296
rect 5832 1296 5850 1314
rect 5832 1314 5850 1332
rect 5832 1332 5850 1350
rect 5832 1350 5850 1368
rect 5832 1368 5850 1386
rect 5832 1386 5850 1404
rect 5832 1404 5850 1422
rect 5832 1422 5850 1440
rect 5832 1440 5850 1458
rect 5832 1458 5850 1476
rect 5832 1476 5850 1494
rect 5832 1494 5850 1512
rect 5832 1512 5850 1530
rect 5832 1530 5850 1548
rect 5832 1548 5850 1566
rect 5832 1566 5850 1584
rect 5832 1584 5850 1602
rect 5832 1602 5850 1620
rect 5832 1620 5850 1638
rect 5832 1638 5850 1656
rect 5832 1656 5850 1674
rect 5832 1674 5850 1692
rect 5832 1692 5850 1710
rect 5832 1710 5850 1728
rect 5832 1728 5850 1746
rect 5832 1746 5850 1764
rect 5832 1764 5850 1782
rect 5832 1782 5850 1800
rect 5832 1800 5850 1818
rect 5832 1818 5850 1836
rect 5832 1836 5850 1854
rect 5832 1854 5850 1872
rect 5832 1872 5850 1890
rect 5832 1890 5850 1908
rect 5832 1908 5850 1926
rect 5832 1926 5850 1944
rect 5832 1944 5850 1962
rect 5832 1962 5850 1980
rect 5832 1980 5850 1998
rect 5832 1998 5850 2016
rect 5832 2016 5850 2034
rect 5832 2034 5850 2052
rect 5832 2052 5850 2070
rect 5832 2070 5850 2088
rect 5832 2088 5850 2106
rect 5832 2106 5850 2124
rect 5832 2124 5850 2142
rect 5832 2142 5850 2160
rect 5832 2160 5850 2178
rect 5832 2178 5850 2196
rect 5832 2196 5850 2214
rect 5832 2214 5850 2232
rect 5832 2232 5850 2250
rect 5832 2250 5850 2268
rect 5832 2268 5850 2286
rect 5832 2286 5850 2304
rect 5832 2304 5850 2322
rect 5832 2322 5850 2340
rect 5832 2340 5850 2358
rect 5832 2358 5850 2376
rect 5832 2376 5850 2394
rect 5832 2394 5850 2412
rect 5832 2412 5850 2430
rect 5832 2430 5850 2448
rect 5832 2448 5850 2466
rect 5832 2466 5850 2484
rect 5832 2484 5850 2502
rect 5832 2502 5850 2520
rect 5832 2520 5850 2538
rect 5832 2538 5850 2556
rect 5832 2556 5850 2574
rect 5832 2574 5850 2592
rect 5832 2592 5850 2610
rect 5832 2610 5850 2628
rect 5832 2628 5850 2646
rect 5832 2646 5850 2664
rect 5832 2664 5850 2682
rect 5832 2898 5850 2916
rect 5832 2916 5850 2934
rect 5832 2934 5850 2952
rect 5832 2952 5850 2970
rect 5832 2970 5850 2988
rect 5832 2988 5850 3006
rect 5832 3006 5850 3024
rect 5832 3024 5850 3042
rect 5832 3042 5850 3060
rect 5832 3060 5850 3078
rect 5832 3078 5850 3096
rect 5832 3096 5850 3114
rect 5832 3114 5850 3132
rect 5832 3132 5850 3150
rect 5832 3150 5850 3168
rect 5832 3168 5850 3186
rect 5832 3186 5850 3204
rect 5832 3204 5850 3222
rect 5832 3222 5850 3240
rect 5832 3240 5850 3258
rect 5832 3258 5850 3276
rect 5832 3276 5850 3294
rect 5832 3294 5850 3312
rect 5832 3312 5850 3330
rect 5832 3330 5850 3348
rect 5832 3348 5850 3366
rect 5832 3366 5850 3384
rect 5832 3384 5850 3402
rect 5832 3402 5850 3420
rect 5832 3420 5850 3438
rect 5832 3438 5850 3456
rect 5832 3456 5850 3474
rect 5832 3474 5850 3492
rect 5832 3492 5850 3510
rect 5832 3510 5850 3528
rect 5832 3528 5850 3546
rect 5832 3546 5850 3564
rect 5832 3564 5850 3582
rect 5832 3582 5850 3600
rect 5832 3600 5850 3618
rect 5832 3618 5850 3636
rect 5832 3636 5850 3654
rect 5832 3654 5850 3672
rect 5832 3672 5850 3690
rect 5832 3690 5850 3708
rect 5832 3708 5850 3726
rect 5832 3726 5850 3744
rect 5832 3744 5850 3762
rect 5832 3762 5850 3780
rect 5832 3780 5850 3798
rect 5832 3798 5850 3816
rect 5832 3816 5850 3834
rect 5832 3834 5850 3852
rect 5832 3852 5850 3870
rect 5832 3870 5850 3888
rect 5832 3888 5850 3906
rect 5832 3906 5850 3924
rect 5832 3924 5850 3942
rect 5832 3942 5850 3960
rect 5832 3960 5850 3978
rect 5832 3978 5850 3996
rect 5832 3996 5850 4014
rect 5832 4014 5850 4032
rect 5832 4032 5850 4050
rect 5832 4050 5850 4068
rect 5832 4068 5850 4086
rect 5832 4086 5850 4104
rect 5832 4104 5850 4122
rect 5832 4122 5850 4140
rect 5832 4140 5850 4158
rect 5832 4158 5850 4176
rect 5832 4176 5850 4194
rect 5832 4194 5850 4212
rect 5832 4212 5850 4230
rect 5832 4230 5850 4248
rect 5832 4248 5850 4266
rect 5832 4266 5850 4284
rect 5832 4284 5850 4302
rect 5832 4302 5850 4320
rect 5832 4320 5850 4338
rect 5832 4338 5850 4356
rect 5832 4356 5850 4374
rect 5832 4374 5850 4392
rect 5832 4392 5850 4410
rect 5832 4410 5850 4428
rect 5832 4428 5850 4446
rect 5832 4446 5850 4464
rect 5832 4464 5850 4482
rect 5832 4482 5850 4500
rect 5832 4500 5850 4518
rect 5832 4518 5850 4536
rect 5832 4536 5850 4554
rect 5832 4554 5850 4572
rect 5832 4572 5850 4590
rect 5832 4590 5850 4608
rect 5832 4608 5850 4626
rect 5832 4626 5850 4644
rect 5832 4644 5850 4662
rect 5832 4662 5850 4680
rect 5832 4680 5850 4698
rect 5832 4698 5850 4716
rect 5832 4716 5850 4734
rect 5832 4734 5850 4752
rect 5832 4752 5850 4770
rect 5832 4770 5850 4788
rect 5832 4788 5850 4806
rect 5832 4806 5850 4824
rect 5832 4824 5850 4842
rect 5832 4842 5850 4860
rect 5832 4860 5850 4878
rect 5832 4878 5850 4896
rect 5832 4896 5850 4914
rect 5832 4914 5850 4932
rect 5832 4932 5850 4950
rect 5832 4950 5850 4968
rect 5832 4968 5850 4986
rect 5832 4986 5850 5004
rect 5832 5004 5850 5022
rect 5832 5022 5850 5040
rect 5832 5040 5850 5058
rect 5832 5058 5850 5076
rect 5832 5076 5850 5094
rect 5832 5094 5850 5112
rect 5832 5112 5850 5130
rect 5832 5130 5850 5148
rect 5832 5148 5850 5166
rect 5832 5166 5850 5184
rect 5832 5184 5850 5202
rect 5832 5202 5850 5220
rect 5832 5472 5850 5490
rect 5832 5490 5850 5508
rect 5832 5508 5850 5526
rect 5832 5526 5850 5544
rect 5832 5544 5850 5562
rect 5832 5562 5850 5580
rect 5832 5580 5850 5598
rect 5832 5598 5850 5616
rect 5832 5616 5850 5634
rect 5832 5634 5850 5652
rect 5832 5652 5850 5670
rect 5832 5670 5850 5688
rect 5832 5688 5850 5706
rect 5832 5706 5850 5724
rect 5832 5724 5850 5742
rect 5832 5742 5850 5760
rect 5832 5760 5850 5778
rect 5832 5778 5850 5796
rect 5832 5796 5850 5814
rect 5832 5814 5850 5832
rect 5832 5832 5850 5850
rect 5832 5850 5850 5868
rect 5832 5868 5850 5886
rect 5832 5886 5850 5904
rect 5832 5904 5850 5922
rect 5832 5922 5850 5940
rect 5832 5940 5850 5958
rect 5832 5958 5850 5976
rect 5832 5976 5850 5994
rect 5832 5994 5850 6012
rect 5832 6012 5850 6030
rect 5832 6030 5850 6048
rect 5832 6048 5850 6066
rect 5832 6066 5850 6084
rect 5832 6084 5850 6102
rect 5832 6102 5850 6120
rect 5832 6120 5850 6138
rect 5832 6138 5850 6156
rect 5832 6156 5850 6174
rect 5832 6174 5850 6192
rect 5832 6192 5850 6210
rect 5832 6210 5850 6228
rect 5832 6228 5850 6246
rect 5832 6246 5850 6264
rect 5832 6264 5850 6282
rect 5832 6282 5850 6300
rect 5832 6300 5850 6318
rect 5832 6318 5850 6336
rect 5832 6336 5850 6354
rect 5832 6354 5850 6372
rect 5832 6372 5850 6390
rect 5832 6390 5850 6408
rect 5832 6408 5850 6426
rect 5832 6426 5850 6444
rect 5832 6444 5850 6462
rect 5832 6462 5850 6480
rect 5832 6480 5850 6498
rect 5832 6498 5850 6516
rect 5832 6516 5850 6534
rect 5832 6534 5850 6552
rect 5832 6552 5850 6570
rect 5832 6570 5850 6588
rect 5832 6588 5850 6606
rect 5832 6606 5850 6624
rect 5832 6624 5850 6642
rect 5832 6642 5850 6660
rect 5832 6660 5850 6678
rect 5832 6678 5850 6696
rect 5832 6696 5850 6714
rect 5832 6714 5850 6732
rect 5832 6732 5850 6750
rect 5832 6750 5850 6768
rect 5832 6768 5850 6786
rect 5832 6786 5850 6804
rect 5832 6804 5850 6822
rect 5832 6822 5850 6840
rect 5832 6840 5850 6858
rect 5832 6858 5850 6876
rect 5832 6876 5850 6894
rect 5832 6894 5850 6912
rect 5832 6912 5850 6930
rect 5832 6930 5850 6948
rect 5832 6948 5850 6966
rect 5832 6966 5850 6984
rect 5832 6984 5850 7002
rect 5832 7002 5850 7020
rect 5832 7020 5850 7038
rect 5832 7038 5850 7056
rect 5832 7056 5850 7074
rect 5832 7074 5850 7092
rect 5832 7092 5850 7110
rect 5832 7110 5850 7128
rect 5832 7128 5850 7146
rect 5832 7146 5850 7164
rect 5832 7164 5850 7182
rect 5832 7182 5850 7200
rect 5832 7200 5850 7218
rect 5832 7218 5850 7236
rect 5832 7236 5850 7254
rect 5832 7254 5850 7272
rect 5832 7272 5850 7290
rect 5832 7290 5850 7308
rect 5832 7308 5850 7326
rect 5832 7326 5850 7344
rect 5832 7344 5850 7362
rect 5832 7362 5850 7380
rect 5832 7380 5850 7398
rect 5832 7398 5850 7416
rect 5832 7416 5850 7434
rect 5832 7434 5850 7452
rect 5832 7452 5850 7470
rect 5832 7470 5850 7488
rect 5832 7488 5850 7506
rect 5832 7506 5850 7524
rect 5832 7524 5850 7542
rect 5832 7542 5850 7560
rect 5832 7560 5850 7578
rect 5832 7578 5850 7596
rect 5832 7596 5850 7614
rect 5832 7614 5850 7632
rect 5832 7632 5850 7650
rect 5832 7650 5850 7668
rect 5832 7668 5850 7686
rect 5832 7686 5850 7704
rect 5832 7704 5850 7722
rect 5832 7722 5850 7740
rect 5832 7740 5850 7758
rect 5832 7758 5850 7776
rect 5832 7776 5850 7794
rect 5832 7794 5850 7812
rect 5832 7812 5850 7830
rect 5832 7830 5850 7848
rect 5832 7848 5850 7866
rect 5832 7866 5850 7884
rect 5832 7884 5850 7902
rect 5832 7902 5850 7920
rect 5832 7920 5850 7938
rect 5832 7938 5850 7956
rect 5832 7956 5850 7974
rect 5832 7974 5850 7992
rect 5832 7992 5850 8010
rect 5832 8010 5850 8028
rect 5832 8028 5850 8046
rect 5832 8046 5850 8064
rect 5832 8064 5850 8082
rect 5832 8082 5850 8100
rect 5832 8100 5850 8118
rect 5832 8118 5850 8136
rect 5832 8136 5850 8154
rect 5832 8154 5850 8172
rect 5832 8172 5850 8190
rect 5832 8190 5850 8208
rect 5832 8208 5850 8226
rect 5832 8226 5850 8244
rect 5832 8244 5850 8262
rect 5832 8262 5850 8280
rect 5832 8280 5850 8298
rect 5832 8298 5850 8316
rect 5832 8316 5850 8334
rect 5832 8334 5850 8352
rect 5832 8352 5850 8370
rect 5832 8370 5850 8388
rect 5832 8388 5850 8406
rect 5832 8406 5850 8424
rect 5832 8424 5850 8442
rect 5832 8442 5850 8460
rect 5832 8460 5850 8478
rect 5832 8478 5850 8496
rect 5832 8496 5850 8514
rect 5832 8514 5850 8532
rect 5832 8532 5850 8550
rect 5832 8550 5850 8568
rect 5832 8568 5850 8586
rect 5832 8586 5850 8604
rect 5832 8604 5850 8622
rect 5832 8622 5850 8640
rect 5832 8640 5850 8658
rect 5832 8658 5850 8676
rect 5832 8676 5850 8694
rect 5832 8694 5850 8712
rect 5832 8712 5850 8730
rect 5832 8730 5850 8748
rect 5832 8748 5850 8766
rect 5832 8766 5850 8784
rect 5832 8784 5850 8802
rect 5832 8802 5850 8820
rect 5832 8820 5850 8838
rect 5832 8838 5850 8856
rect 5832 8856 5850 8874
rect 5832 8874 5850 8892
rect 5832 8892 5850 8910
rect 5832 8910 5850 8928
rect 5832 8928 5850 8946
rect 5832 8946 5850 8964
rect 5832 8964 5850 8982
rect 5832 8982 5850 9000
rect 5832 9000 5850 9018
rect 5850 774 5868 792
rect 5850 792 5868 810
rect 5850 810 5868 828
rect 5850 828 5868 846
rect 5850 846 5868 864
rect 5850 864 5868 882
rect 5850 882 5868 900
rect 5850 900 5868 918
rect 5850 918 5868 936
rect 5850 936 5868 954
rect 5850 954 5868 972
rect 5850 972 5868 990
rect 5850 990 5868 1008
rect 5850 1008 5868 1026
rect 5850 1026 5868 1044
rect 5850 1188 5868 1206
rect 5850 1206 5868 1224
rect 5850 1224 5868 1242
rect 5850 1242 5868 1260
rect 5850 1260 5868 1278
rect 5850 1278 5868 1296
rect 5850 1296 5868 1314
rect 5850 1314 5868 1332
rect 5850 1332 5868 1350
rect 5850 1350 5868 1368
rect 5850 1368 5868 1386
rect 5850 1386 5868 1404
rect 5850 1404 5868 1422
rect 5850 1422 5868 1440
rect 5850 1440 5868 1458
rect 5850 1458 5868 1476
rect 5850 1476 5868 1494
rect 5850 1494 5868 1512
rect 5850 1512 5868 1530
rect 5850 1530 5868 1548
rect 5850 1548 5868 1566
rect 5850 1566 5868 1584
rect 5850 1584 5868 1602
rect 5850 1602 5868 1620
rect 5850 1620 5868 1638
rect 5850 1638 5868 1656
rect 5850 1656 5868 1674
rect 5850 1674 5868 1692
rect 5850 1692 5868 1710
rect 5850 1710 5868 1728
rect 5850 1728 5868 1746
rect 5850 1746 5868 1764
rect 5850 1764 5868 1782
rect 5850 1782 5868 1800
rect 5850 1800 5868 1818
rect 5850 1818 5868 1836
rect 5850 1836 5868 1854
rect 5850 1854 5868 1872
rect 5850 1872 5868 1890
rect 5850 1890 5868 1908
rect 5850 1908 5868 1926
rect 5850 1926 5868 1944
rect 5850 1944 5868 1962
rect 5850 1962 5868 1980
rect 5850 1980 5868 1998
rect 5850 1998 5868 2016
rect 5850 2016 5868 2034
rect 5850 2034 5868 2052
rect 5850 2052 5868 2070
rect 5850 2070 5868 2088
rect 5850 2088 5868 2106
rect 5850 2106 5868 2124
rect 5850 2124 5868 2142
rect 5850 2142 5868 2160
rect 5850 2160 5868 2178
rect 5850 2178 5868 2196
rect 5850 2196 5868 2214
rect 5850 2214 5868 2232
rect 5850 2232 5868 2250
rect 5850 2250 5868 2268
rect 5850 2268 5868 2286
rect 5850 2286 5868 2304
rect 5850 2304 5868 2322
rect 5850 2322 5868 2340
rect 5850 2340 5868 2358
rect 5850 2358 5868 2376
rect 5850 2376 5868 2394
rect 5850 2394 5868 2412
rect 5850 2412 5868 2430
rect 5850 2430 5868 2448
rect 5850 2448 5868 2466
rect 5850 2466 5868 2484
rect 5850 2484 5868 2502
rect 5850 2502 5868 2520
rect 5850 2520 5868 2538
rect 5850 2538 5868 2556
rect 5850 2556 5868 2574
rect 5850 2574 5868 2592
rect 5850 2592 5868 2610
rect 5850 2610 5868 2628
rect 5850 2628 5868 2646
rect 5850 2646 5868 2664
rect 5850 2664 5868 2682
rect 5850 2916 5868 2934
rect 5850 2934 5868 2952
rect 5850 2952 5868 2970
rect 5850 2970 5868 2988
rect 5850 2988 5868 3006
rect 5850 3006 5868 3024
rect 5850 3024 5868 3042
rect 5850 3042 5868 3060
rect 5850 3060 5868 3078
rect 5850 3078 5868 3096
rect 5850 3096 5868 3114
rect 5850 3114 5868 3132
rect 5850 3132 5868 3150
rect 5850 3150 5868 3168
rect 5850 3168 5868 3186
rect 5850 3186 5868 3204
rect 5850 3204 5868 3222
rect 5850 3222 5868 3240
rect 5850 3240 5868 3258
rect 5850 3258 5868 3276
rect 5850 3276 5868 3294
rect 5850 3294 5868 3312
rect 5850 3312 5868 3330
rect 5850 3330 5868 3348
rect 5850 3348 5868 3366
rect 5850 3366 5868 3384
rect 5850 3384 5868 3402
rect 5850 3402 5868 3420
rect 5850 3420 5868 3438
rect 5850 3438 5868 3456
rect 5850 3456 5868 3474
rect 5850 3474 5868 3492
rect 5850 3492 5868 3510
rect 5850 3510 5868 3528
rect 5850 3528 5868 3546
rect 5850 3546 5868 3564
rect 5850 3564 5868 3582
rect 5850 3582 5868 3600
rect 5850 3600 5868 3618
rect 5850 3618 5868 3636
rect 5850 3636 5868 3654
rect 5850 3654 5868 3672
rect 5850 3672 5868 3690
rect 5850 3690 5868 3708
rect 5850 3708 5868 3726
rect 5850 3726 5868 3744
rect 5850 3744 5868 3762
rect 5850 3762 5868 3780
rect 5850 3780 5868 3798
rect 5850 3798 5868 3816
rect 5850 3816 5868 3834
rect 5850 3834 5868 3852
rect 5850 3852 5868 3870
rect 5850 3870 5868 3888
rect 5850 3888 5868 3906
rect 5850 3906 5868 3924
rect 5850 3924 5868 3942
rect 5850 3942 5868 3960
rect 5850 3960 5868 3978
rect 5850 3978 5868 3996
rect 5850 3996 5868 4014
rect 5850 4014 5868 4032
rect 5850 4032 5868 4050
rect 5850 4050 5868 4068
rect 5850 4068 5868 4086
rect 5850 4086 5868 4104
rect 5850 4104 5868 4122
rect 5850 4122 5868 4140
rect 5850 4140 5868 4158
rect 5850 4158 5868 4176
rect 5850 4176 5868 4194
rect 5850 4194 5868 4212
rect 5850 4212 5868 4230
rect 5850 4230 5868 4248
rect 5850 4248 5868 4266
rect 5850 4266 5868 4284
rect 5850 4284 5868 4302
rect 5850 4302 5868 4320
rect 5850 4320 5868 4338
rect 5850 4338 5868 4356
rect 5850 4356 5868 4374
rect 5850 4374 5868 4392
rect 5850 4392 5868 4410
rect 5850 4410 5868 4428
rect 5850 4428 5868 4446
rect 5850 4446 5868 4464
rect 5850 4464 5868 4482
rect 5850 4482 5868 4500
rect 5850 4500 5868 4518
rect 5850 4518 5868 4536
rect 5850 4536 5868 4554
rect 5850 4554 5868 4572
rect 5850 4572 5868 4590
rect 5850 4590 5868 4608
rect 5850 4608 5868 4626
rect 5850 4626 5868 4644
rect 5850 4644 5868 4662
rect 5850 4662 5868 4680
rect 5850 4680 5868 4698
rect 5850 4698 5868 4716
rect 5850 4716 5868 4734
rect 5850 4734 5868 4752
rect 5850 4752 5868 4770
rect 5850 4770 5868 4788
rect 5850 4788 5868 4806
rect 5850 4806 5868 4824
rect 5850 4824 5868 4842
rect 5850 4842 5868 4860
rect 5850 4860 5868 4878
rect 5850 4878 5868 4896
rect 5850 4896 5868 4914
rect 5850 4914 5868 4932
rect 5850 4932 5868 4950
rect 5850 4950 5868 4968
rect 5850 4968 5868 4986
rect 5850 4986 5868 5004
rect 5850 5004 5868 5022
rect 5850 5022 5868 5040
rect 5850 5040 5868 5058
rect 5850 5058 5868 5076
rect 5850 5076 5868 5094
rect 5850 5094 5868 5112
rect 5850 5112 5868 5130
rect 5850 5130 5868 5148
rect 5850 5148 5868 5166
rect 5850 5166 5868 5184
rect 5850 5184 5868 5202
rect 5850 5202 5868 5220
rect 5850 5220 5868 5238
rect 5850 5490 5868 5508
rect 5850 5508 5868 5526
rect 5850 5526 5868 5544
rect 5850 5544 5868 5562
rect 5850 5562 5868 5580
rect 5850 5580 5868 5598
rect 5850 5598 5868 5616
rect 5850 5616 5868 5634
rect 5850 5634 5868 5652
rect 5850 5652 5868 5670
rect 5850 5670 5868 5688
rect 5850 5688 5868 5706
rect 5850 5706 5868 5724
rect 5850 5724 5868 5742
rect 5850 5742 5868 5760
rect 5850 5760 5868 5778
rect 5850 5778 5868 5796
rect 5850 5796 5868 5814
rect 5850 5814 5868 5832
rect 5850 5832 5868 5850
rect 5850 5850 5868 5868
rect 5850 5868 5868 5886
rect 5850 5886 5868 5904
rect 5850 5904 5868 5922
rect 5850 5922 5868 5940
rect 5850 5940 5868 5958
rect 5850 5958 5868 5976
rect 5850 5976 5868 5994
rect 5850 5994 5868 6012
rect 5850 6012 5868 6030
rect 5850 6030 5868 6048
rect 5850 6048 5868 6066
rect 5850 6066 5868 6084
rect 5850 6084 5868 6102
rect 5850 6102 5868 6120
rect 5850 6120 5868 6138
rect 5850 6138 5868 6156
rect 5850 6156 5868 6174
rect 5850 6174 5868 6192
rect 5850 6192 5868 6210
rect 5850 6210 5868 6228
rect 5850 6228 5868 6246
rect 5850 6246 5868 6264
rect 5850 6264 5868 6282
rect 5850 6282 5868 6300
rect 5850 6300 5868 6318
rect 5850 6318 5868 6336
rect 5850 6336 5868 6354
rect 5850 6354 5868 6372
rect 5850 6372 5868 6390
rect 5850 6390 5868 6408
rect 5850 6408 5868 6426
rect 5850 6426 5868 6444
rect 5850 6444 5868 6462
rect 5850 6462 5868 6480
rect 5850 6480 5868 6498
rect 5850 6498 5868 6516
rect 5850 6516 5868 6534
rect 5850 6534 5868 6552
rect 5850 6552 5868 6570
rect 5850 6570 5868 6588
rect 5850 6588 5868 6606
rect 5850 6606 5868 6624
rect 5850 6624 5868 6642
rect 5850 6642 5868 6660
rect 5850 6660 5868 6678
rect 5850 6678 5868 6696
rect 5850 6696 5868 6714
rect 5850 6714 5868 6732
rect 5850 6732 5868 6750
rect 5850 6750 5868 6768
rect 5850 6768 5868 6786
rect 5850 6786 5868 6804
rect 5850 6804 5868 6822
rect 5850 6822 5868 6840
rect 5850 6840 5868 6858
rect 5850 6858 5868 6876
rect 5850 6876 5868 6894
rect 5850 6894 5868 6912
rect 5850 6912 5868 6930
rect 5850 6930 5868 6948
rect 5850 6948 5868 6966
rect 5850 6966 5868 6984
rect 5850 6984 5868 7002
rect 5850 7002 5868 7020
rect 5850 7020 5868 7038
rect 5850 7038 5868 7056
rect 5850 7056 5868 7074
rect 5850 7074 5868 7092
rect 5850 7092 5868 7110
rect 5850 7110 5868 7128
rect 5850 7128 5868 7146
rect 5850 7146 5868 7164
rect 5850 7164 5868 7182
rect 5850 7182 5868 7200
rect 5850 7200 5868 7218
rect 5850 7218 5868 7236
rect 5850 7236 5868 7254
rect 5850 7254 5868 7272
rect 5850 7272 5868 7290
rect 5850 7290 5868 7308
rect 5850 7308 5868 7326
rect 5850 7326 5868 7344
rect 5850 7344 5868 7362
rect 5850 7362 5868 7380
rect 5850 7380 5868 7398
rect 5850 7398 5868 7416
rect 5850 7416 5868 7434
rect 5850 7434 5868 7452
rect 5850 7452 5868 7470
rect 5850 7470 5868 7488
rect 5850 7488 5868 7506
rect 5850 7506 5868 7524
rect 5850 7524 5868 7542
rect 5850 7542 5868 7560
rect 5850 7560 5868 7578
rect 5850 7578 5868 7596
rect 5850 7596 5868 7614
rect 5850 7614 5868 7632
rect 5850 7632 5868 7650
rect 5850 7650 5868 7668
rect 5850 7668 5868 7686
rect 5850 7686 5868 7704
rect 5850 7704 5868 7722
rect 5850 7722 5868 7740
rect 5850 7740 5868 7758
rect 5850 7758 5868 7776
rect 5850 7776 5868 7794
rect 5850 7794 5868 7812
rect 5850 7812 5868 7830
rect 5850 7830 5868 7848
rect 5850 7848 5868 7866
rect 5850 7866 5868 7884
rect 5850 7884 5868 7902
rect 5850 7902 5868 7920
rect 5850 7920 5868 7938
rect 5850 7938 5868 7956
rect 5850 7956 5868 7974
rect 5850 7974 5868 7992
rect 5850 7992 5868 8010
rect 5850 8010 5868 8028
rect 5850 8028 5868 8046
rect 5850 8046 5868 8064
rect 5850 8064 5868 8082
rect 5850 8082 5868 8100
rect 5850 8100 5868 8118
rect 5850 8118 5868 8136
rect 5850 8136 5868 8154
rect 5850 8154 5868 8172
rect 5850 8172 5868 8190
rect 5850 8190 5868 8208
rect 5850 8208 5868 8226
rect 5850 8226 5868 8244
rect 5850 8244 5868 8262
rect 5850 8262 5868 8280
rect 5850 8280 5868 8298
rect 5850 8298 5868 8316
rect 5850 8316 5868 8334
rect 5850 8334 5868 8352
rect 5850 8352 5868 8370
rect 5850 8370 5868 8388
rect 5850 8388 5868 8406
rect 5850 8406 5868 8424
rect 5850 8424 5868 8442
rect 5850 8442 5868 8460
rect 5850 8460 5868 8478
rect 5850 8478 5868 8496
rect 5850 8496 5868 8514
rect 5850 8514 5868 8532
rect 5850 8532 5868 8550
rect 5850 8550 5868 8568
rect 5850 8568 5868 8586
rect 5850 8586 5868 8604
rect 5850 8604 5868 8622
rect 5850 8622 5868 8640
rect 5850 8640 5868 8658
rect 5850 8658 5868 8676
rect 5850 8676 5868 8694
rect 5850 8694 5868 8712
rect 5850 8712 5868 8730
rect 5850 8730 5868 8748
rect 5850 8748 5868 8766
rect 5850 8766 5868 8784
rect 5850 8784 5868 8802
rect 5850 8802 5868 8820
rect 5850 8820 5868 8838
rect 5850 8838 5868 8856
rect 5850 8856 5868 8874
rect 5850 8874 5868 8892
rect 5850 8892 5868 8910
rect 5850 8910 5868 8928
rect 5850 8928 5868 8946
rect 5850 8946 5868 8964
rect 5850 8964 5868 8982
rect 5850 8982 5868 9000
rect 5850 9000 5868 9018
rect 5850 9018 5868 9036
rect 5868 792 5886 810
rect 5868 810 5886 828
rect 5868 828 5886 846
rect 5868 846 5886 864
rect 5868 864 5886 882
rect 5868 882 5886 900
rect 5868 900 5886 918
rect 5868 918 5886 936
rect 5868 936 5886 954
rect 5868 954 5886 972
rect 5868 972 5886 990
rect 5868 990 5886 1008
rect 5868 1008 5886 1026
rect 5868 1026 5886 1044
rect 5868 1044 5886 1062
rect 5868 1206 5886 1224
rect 5868 1224 5886 1242
rect 5868 1242 5886 1260
rect 5868 1260 5886 1278
rect 5868 1278 5886 1296
rect 5868 1296 5886 1314
rect 5868 1314 5886 1332
rect 5868 1332 5886 1350
rect 5868 1350 5886 1368
rect 5868 1368 5886 1386
rect 5868 1386 5886 1404
rect 5868 1404 5886 1422
rect 5868 1422 5886 1440
rect 5868 1440 5886 1458
rect 5868 1458 5886 1476
rect 5868 1476 5886 1494
rect 5868 1494 5886 1512
rect 5868 1512 5886 1530
rect 5868 1530 5886 1548
rect 5868 1548 5886 1566
rect 5868 1566 5886 1584
rect 5868 1584 5886 1602
rect 5868 1602 5886 1620
rect 5868 1620 5886 1638
rect 5868 1638 5886 1656
rect 5868 1656 5886 1674
rect 5868 1674 5886 1692
rect 5868 1692 5886 1710
rect 5868 1710 5886 1728
rect 5868 1728 5886 1746
rect 5868 1746 5886 1764
rect 5868 1764 5886 1782
rect 5868 1782 5886 1800
rect 5868 1800 5886 1818
rect 5868 1818 5886 1836
rect 5868 1836 5886 1854
rect 5868 1854 5886 1872
rect 5868 1872 5886 1890
rect 5868 1890 5886 1908
rect 5868 1908 5886 1926
rect 5868 1926 5886 1944
rect 5868 1944 5886 1962
rect 5868 1962 5886 1980
rect 5868 1980 5886 1998
rect 5868 1998 5886 2016
rect 5868 2016 5886 2034
rect 5868 2034 5886 2052
rect 5868 2052 5886 2070
rect 5868 2070 5886 2088
rect 5868 2088 5886 2106
rect 5868 2106 5886 2124
rect 5868 2124 5886 2142
rect 5868 2142 5886 2160
rect 5868 2160 5886 2178
rect 5868 2178 5886 2196
rect 5868 2196 5886 2214
rect 5868 2214 5886 2232
rect 5868 2232 5886 2250
rect 5868 2250 5886 2268
rect 5868 2268 5886 2286
rect 5868 2286 5886 2304
rect 5868 2304 5886 2322
rect 5868 2322 5886 2340
rect 5868 2340 5886 2358
rect 5868 2358 5886 2376
rect 5868 2376 5886 2394
rect 5868 2394 5886 2412
rect 5868 2412 5886 2430
rect 5868 2430 5886 2448
rect 5868 2448 5886 2466
rect 5868 2466 5886 2484
rect 5868 2484 5886 2502
rect 5868 2502 5886 2520
rect 5868 2520 5886 2538
rect 5868 2538 5886 2556
rect 5868 2556 5886 2574
rect 5868 2574 5886 2592
rect 5868 2592 5886 2610
rect 5868 2610 5886 2628
rect 5868 2628 5886 2646
rect 5868 2646 5886 2664
rect 5868 2664 5886 2682
rect 5868 2682 5886 2700
rect 5868 2916 5886 2934
rect 5868 2934 5886 2952
rect 5868 2952 5886 2970
rect 5868 2970 5886 2988
rect 5868 2988 5886 3006
rect 5868 3006 5886 3024
rect 5868 3024 5886 3042
rect 5868 3042 5886 3060
rect 5868 3060 5886 3078
rect 5868 3078 5886 3096
rect 5868 3096 5886 3114
rect 5868 3114 5886 3132
rect 5868 3132 5886 3150
rect 5868 3150 5886 3168
rect 5868 3168 5886 3186
rect 5868 3186 5886 3204
rect 5868 3204 5886 3222
rect 5868 3222 5886 3240
rect 5868 3240 5886 3258
rect 5868 3258 5886 3276
rect 5868 3276 5886 3294
rect 5868 3294 5886 3312
rect 5868 3312 5886 3330
rect 5868 3330 5886 3348
rect 5868 3348 5886 3366
rect 5868 3366 5886 3384
rect 5868 3384 5886 3402
rect 5868 3402 5886 3420
rect 5868 3420 5886 3438
rect 5868 3438 5886 3456
rect 5868 3456 5886 3474
rect 5868 3474 5886 3492
rect 5868 3492 5886 3510
rect 5868 3510 5886 3528
rect 5868 3528 5886 3546
rect 5868 3546 5886 3564
rect 5868 3564 5886 3582
rect 5868 3582 5886 3600
rect 5868 3600 5886 3618
rect 5868 3618 5886 3636
rect 5868 3636 5886 3654
rect 5868 3654 5886 3672
rect 5868 3672 5886 3690
rect 5868 3690 5886 3708
rect 5868 3708 5886 3726
rect 5868 3726 5886 3744
rect 5868 3744 5886 3762
rect 5868 3762 5886 3780
rect 5868 3780 5886 3798
rect 5868 3798 5886 3816
rect 5868 3816 5886 3834
rect 5868 3834 5886 3852
rect 5868 3852 5886 3870
rect 5868 3870 5886 3888
rect 5868 3888 5886 3906
rect 5868 3906 5886 3924
rect 5868 3924 5886 3942
rect 5868 3942 5886 3960
rect 5868 3960 5886 3978
rect 5868 3978 5886 3996
rect 5868 3996 5886 4014
rect 5868 4014 5886 4032
rect 5868 4032 5886 4050
rect 5868 4050 5886 4068
rect 5868 4068 5886 4086
rect 5868 4086 5886 4104
rect 5868 4104 5886 4122
rect 5868 4122 5886 4140
rect 5868 4140 5886 4158
rect 5868 4158 5886 4176
rect 5868 4176 5886 4194
rect 5868 4194 5886 4212
rect 5868 4212 5886 4230
rect 5868 4230 5886 4248
rect 5868 4248 5886 4266
rect 5868 4266 5886 4284
rect 5868 4284 5886 4302
rect 5868 4302 5886 4320
rect 5868 4320 5886 4338
rect 5868 4338 5886 4356
rect 5868 4356 5886 4374
rect 5868 4374 5886 4392
rect 5868 4392 5886 4410
rect 5868 4410 5886 4428
rect 5868 4428 5886 4446
rect 5868 4446 5886 4464
rect 5868 4464 5886 4482
rect 5868 4482 5886 4500
rect 5868 4500 5886 4518
rect 5868 4518 5886 4536
rect 5868 4536 5886 4554
rect 5868 4554 5886 4572
rect 5868 4572 5886 4590
rect 5868 4590 5886 4608
rect 5868 4608 5886 4626
rect 5868 4626 5886 4644
rect 5868 4644 5886 4662
rect 5868 4662 5886 4680
rect 5868 4680 5886 4698
rect 5868 4698 5886 4716
rect 5868 4716 5886 4734
rect 5868 4734 5886 4752
rect 5868 4752 5886 4770
rect 5868 4770 5886 4788
rect 5868 4788 5886 4806
rect 5868 4806 5886 4824
rect 5868 4824 5886 4842
rect 5868 4842 5886 4860
rect 5868 4860 5886 4878
rect 5868 4878 5886 4896
rect 5868 4896 5886 4914
rect 5868 4914 5886 4932
rect 5868 4932 5886 4950
rect 5868 4950 5886 4968
rect 5868 4968 5886 4986
rect 5868 4986 5886 5004
rect 5868 5004 5886 5022
rect 5868 5022 5886 5040
rect 5868 5040 5886 5058
rect 5868 5058 5886 5076
rect 5868 5076 5886 5094
rect 5868 5094 5886 5112
rect 5868 5112 5886 5130
rect 5868 5130 5886 5148
rect 5868 5148 5886 5166
rect 5868 5166 5886 5184
rect 5868 5184 5886 5202
rect 5868 5202 5886 5220
rect 5868 5220 5886 5238
rect 5868 5238 5886 5256
rect 5868 5508 5886 5526
rect 5868 5526 5886 5544
rect 5868 5544 5886 5562
rect 5868 5562 5886 5580
rect 5868 5580 5886 5598
rect 5868 5598 5886 5616
rect 5868 5616 5886 5634
rect 5868 5634 5886 5652
rect 5868 5652 5886 5670
rect 5868 5670 5886 5688
rect 5868 5688 5886 5706
rect 5868 5706 5886 5724
rect 5868 5724 5886 5742
rect 5868 5742 5886 5760
rect 5868 5760 5886 5778
rect 5868 5778 5886 5796
rect 5868 5796 5886 5814
rect 5868 5814 5886 5832
rect 5868 5832 5886 5850
rect 5868 5850 5886 5868
rect 5868 5868 5886 5886
rect 5868 5886 5886 5904
rect 5868 5904 5886 5922
rect 5868 5922 5886 5940
rect 5868 5940 5886 5958
rect 5868 5958 5886 5976
rect 5868 5976 5886 5994
rect 5868 5994 5886 6012
rect 5868 6012 5886 6030
rect 5868 6030 5886 6048
rect 5868 6048 5886 6066
rect 5868 6066 5886 6084
rect 5868 6084 5886 6102
rect 5868 6102 5886 6120
rect 5868 6120 5886 6138
rect 5868 6138 5886 6156
rect 5868 6156 5886 6174
rect 5868 6174 5886 6192
rect 5868 6192 5886 6210
rect 5868 6210 5886 6228
rect 5868 6228 5886 6246
rect 5868 6246 5886 6264
rect 5868 6264 5886 6282
rect 5868 6282 5886 6300
rect 5868 6300 5886 6318
rect 5868 6318 5886 6336
rect 5868 6336 5886 6354
rect 5868 6354 5886 6372
rect 5868 6372 5886 6390
rect 5868 6390 5886 6408
rect 5868 6408 5886 6426
rect 5868 6426 5886 6444
rect 5868 6444 5886 6462
rect 5868 6462 5886 6480
rect 5868 6480 5886 6498
rect 5868 6498 5886 6516
rect 5868 6516 5886 6534
rect 5868 6534 5886 6552
rect 5868 6552 5886 6570
rect 5868 6570 5886 6588
rect 5868 6588 5886 6606
rect 5868 6606 5886 6624
rect 5868 6624 5886 6642
rect 5868 6642 5886 6660
rect 5868 6660 5886 6678
rect 5868 6678 5886 6696
rect 5868 6696 5886 6714
rect 5868 6714 5886 6732
rect 5868 6732 5886 6750
rect 5868 6750 5886 6768
rect 5868 6768 5886 6786
rect 5868 6786 5886 6804
rect 5868 6804 5886 6822
rect 5868 6822 5886 6840
rect 5868 6840 5886 6858
rect 5868 6858 5886 6876
rect 5868 6876 5886 6894
rect 5868 6894 5886 6912
rect 5868 6912 5886 6930
rect 5868 6930 5886 6948
rect 5868 6948 5886 6966
rect 5868 6966 5886 6984
rect 5868 6984 5886 7002
rect 5868 7002 5886 7020
rect 5868 7020 5886 7038
rect 5868 7038 5886 7056
rect 5868 7056 5886 7074
rect 5868 7074 5886 7092
rect 5868 7092 5886 7110
rect 5868 7110 5886 7128
rect 5868 7128 5886 7146
rect 5868 7146 5886 7164
rect 5868 7164 5886 7182
rect 5868 7182 5886 7200
rect 5868 7200 5886 7218
rect 5868 7218 5886 7236
rect 5868 7236 5886 7254
rect 5868 7254 5886 7272
rect 5868 7272 5886 7290
rect 5868 7290 5886 7308
rect 5868 7308 5886 7326
rect 5868 7326 5886 7344
rect 5868 7344 5886 7362
rect 5868 7362 5886 7380
rect 5868 7380 5886 7398
rect 5868 7398 5886 7416
rect 5868 7416 5886 7434
rect 5868 7434 5886 7452
rect 5868 7452 5886 7470
rect 5868 7470 5886 7488
rect 5868 7488 5886 7506
rect 5868 7506 5886 7524
rect 5868 7524 5886 7542
rect 5868 7542 5886 7560
rect 5868 7560 5886 7578
rect 5868 7578 5886 7596
rect 5868 7596 5886 7614
rect 5868 7614 5886 7632
rect 5868 7632 5886 7650
rect 5868 7650 5886 7668
rect 5868 7668 5886 7686
rect 5868 7686 5886 7704
rect 5868 7704 5886 7722
rect 5868 7722 5886 7740
rect 5868 7740 5886 7758
rect 5868 7758 5886 7776
rect 5868 7776 5886 7794
rect 5868 7794 5886 7812
rect 5868 7812 5886 7830
rect 5868 7830 5886 7848
rect 5868 7848 5886 7866
rect 5868 7866 5886 7884
rect 5868 7884 5886 7902
rect 5868 7902 5886 7920
rect 5868 7920 5886 7938
rect 5868 7938 5886 7956
rect 5868 7956 5886 7974
rect 5868 7974 5886 7992
rect 5868 7992 5886 8010
rect 5868 8010 5886 8028
rect 5868 8028 5886 8046
rect 5868 8046 5886 8064
rect 5868 8064 5886 8082
rect 5868 8082 5886 8100
rect 5868 8100 5886 8118
rect 5868 8118 5886 8136
rect 5868 8136 5886 8154
rect 5868 8154 5886 8172
rect 5868 8172 5886 8190
rect 5868 8190 5886 8208
rect 5868 8208 5886 8226
rect 5868 8226 5886 8244
rect 5868 8244 5886 8262
rect 5868 8262 5886 8280
rect 5868 8280 5886 8298
rect 5868 8298 5886 8316
rect 5868 8316 5886 8334
rect 5868 8334 5886 8352
rect 5868 8352 5886 8370
rect 5868 8370 5886 8388
rect 5868 8388 5886 8406
rect 5868 8406 5886 8424
rect 5868 8424 5886 8442
rect 5868 8442 5886 8460
rect 5868 8460 5886 8478
rect 5868 8478 5886 8496
rect 5868 8496 5886 8514
rect 5868 8514 5886 8532
rect 5868 8532 5886 8550
rect 5868 8550 5886 8568
rect 5868 8568 5886 8586
rect 5868 8586 5886 8604
rect 5868 8604 5886 8622
rect 5868 8622 5886 8640
rect 5868 8640 5886 8658
rect 5868 8658 5886 8676
rect 5868 8676 5886 8694
rect 5868 8694 5886 8712
rect 5868 8712 5886 8730
rect 5868 8730 5886 8748
rect 5868 8748 5886 8766
rect 5868 8766 5886 8784
rect 5868 8784 5886 8802
rect 5868 8802 5886 8820
rect 5868 8820 5886 8838
rect 5868 8838 5886 8856
rect 5868 8856 5886 8874
rect 5868 8874 5886 8892
rect 5868 8892 5886 8910
rect 5868 8910 5886 8928
rect 5868 8928 5886 8946
rect 5868 8946 5886 8964
rect 5868 8964 5886 8982
rect 5868 8982 5886 9000
rect 5868 9000 5886 9018
rect 5868 9018 5886 9036
rect 5868 9036 5886 9054
rect 5886 810 5904 828
rect 5886 828 5904 846
rect 5886 846 5904 864
rect 5886 864 5904 882
rect 5886 882 5904 900
rect 5886 900 5904 918
rect 5886 918 5904 936
rect 5886 936 5904 954
rect 5886 954 5904 972
rect 5886 972 5904 990
rect 5886 990 5904 1008
rect 5886 1008 5904 1026
rect 5886 1026 5904 1044
rect 5886 1044 5904 1062
rect 5886 1206 5904 1224
rect 5886 1224 5904 1242
rect 5886 1242 5904 1260
rect 5886 1260 5904 1278
rect 5886 1278 5904 1296
rect 5886 1296 5904 1314
rect 5886 1314 5904 1332
rect 5886 1332 5904 1350
rect 5886 1350 5904 1368
rect 5886 1368 5904 1386
rect 5886 1386 5904 1404
rect 5886 1404 5904 1422
rect 5886 1422 5904 1440
rect 5886 1440 5904 1458
rect 5886 1458 5904 1476
rect 5886 1476 5904 1494
rect 5886 1494 5904 1512
rect 5886 1512 5904 1530
rect 5886 1530 5904 1548
rect 5886 1548 5904 1566
rect 5886 1566 5904 1584
rect 5886 1584 5904 1602
rect 5886 1602 5904 1620
rect 5886 1620 5904 1638
rect 5886 1638 5904 1656
rect 5886 1656 5904 1674
rect 5886 1674 5904 1692
rect 5886 1692 5904 1710
rect 5886 1710 5904 1728
rect 5886 1728 5904 1746
rect 5886 1746 5904 1764
rect 5886 1764 5904 1782
rect 5886 1782 5904 1800
rect 5886 1800 5904 1818
rect 5886 1818 5904 1836
rect 5886 1836 5904 1854
rect 5886 1854 5904 1872
rect 5886 1872 5904 1890
rect 5886 1890 5904 1908
rect 5886 1908 5904 1926
rect 5886 1926 5904 1944
rect 5886 1944 5904 1962
rect 5886 1962 5904 1980
rect 5886 1980 5904 1998
rect 5886 1998 5904 2016
rect 5886 2016 5904 2034
rect 5886 2034 5904 2052
rect 5886 2052 5904 2070
rect 5886 2070 5904 2088
rect 5886 2088 5904 2106
rect 5886 2106 5904 2124
rect 5886 2124 5904 2142
rect 5886 2142 5904 2160
rect 5886 2160 5904 2178
rect 5886 2178 5904 2196
rect 5886 2196 5904 2214
rect 5886 2214 5904 2232
rect 5886 2232 5904 2250
rect 5886 2250 5904 2268
rect 5886 2268 5904 2286
rect 5886 2286 5904 2304
rect 5886 2304 5904 2322
rect 5886 2322 5904 2340
rect 5886 2340 5904 2358
rect 5886 2358 5904 2376
rect 5886 2376 5904 2394
rect 5886 2394 5904 2412
rect 5886 2412 5904 2430
rect 5886 2430 5904 2448
rect 5886 2448 5904 2466
rect 5886 2466 5904 2484
rect 5886 2484 5904 2502
rect 5886 2502 5904 2520
rect 5886 2520 5904 2538
rect 5886 2538 5904 2556
rect 5886 2556 5904 2574
rect 5886 2574 5904 2592
rect 5886 2592 5904 2610
rect 5886 2610 5904 2628
rect 5886 2628 5904 2646
rect 5886 2646 5904 2664
rect 5886 2664 5904 2682
rect 5886 2682 5904 2700
rect 5886 2934 5904 2952
rect 5886 2952 5904 2970
rect 5886 2970 5904 2988
rect 5886 2988 5904 3006
rect 5886 3006 5904 3024
rect 5886 3024 5904 3042
rect 5886 3042 5904 3060
rect 5886 3060 5904 3078
rect 5886 3078 5904 3096
rect 5886 3096 5904 3114
rect 5886 3114 5904 3132
rect 5886 3132 5904 3150
rect 5886 3150 5904 3168
rect 5886 3168 5904 3186
rect 5886 3186 5904 3204
rect 5886 3204 5904 3222
rect 5886 3222 5904 3240
rect 5886 3240 5904 3258
rect 5886 3258 5904 3276
rect 5886 3276 5904 3294
rect 5886 3294 5904 3312
rect 5886 3312 5904 3330
rect 5886 3330 5904 3348
rect 5886 3348 5904 3366
rect 5886 3366 5904 3384
rect 5886 3384 5904 3402
rect 5886 3402 5904 3420
rect 5886 3420 5904 3438
rect 5886 3438 5904 3456
rect 5886 3456 5904 3474
rect 5886 3474 5904 3492
rect 5886 3492 5904 3510
rect 5886 3510 5904 3528
rect 5886 3528 5904 3546
rect 5886 3546 5904 3564
rect 5886 3564 5904 3582
rect 5886 3582 5904 3600
rect 5886 3600 5904 3618
rect 5886 3618 5904 3636
rect 5886 3636 5904 3654
rect 5886 3654 5904 3672
rect 5886 3672 5904 3690
rect 5886 3690 5904 3708
rect 5886 3708 5904 3726
rect 5886 3726 5904 3744
rect 5886 3744 5904 3762
rect 5886 3762 5904 3780
rect 5886 3780 5904 3798
rect 5886 3798 5904 3816
rect 5886 3816 5904 3834
rect 5886 3834 5904 3852
rect 5886 3852 5904 3870
rect 5886 3870 5904 3888
rect 5886 3888 5904 3906
rect 5886 3906 5904 3924
rect 5886 3924 5904 3942
rect 5886 3942 5904 3960
rect 5886 3960 5904 3978
rect 5886 3978 5904 3996
rect 5886 3996 5904 4014
rect 5886 4014 5904 4032
rect 5886 4032 5904 4050
rect 5886 4050 5904 4068
rect 5886 4068 5904 4086
rect 5886 4086 5904 4104
rect 5886 4104 5904 4122
rect 5886 4122 5904 4140
rect 5886 4140 5904 4158
rect 5886 4158 5904 4176
rect 5886 4176 5904 4194
rect 5886 4194 5904 4212
rect 5886 4212 5904 4230
rect 5886 4230 5904 4248
rect 5886 4248 5904 4266
rect 5886 4266 5904 4284
rect 5886 4284 5904 4302
rect 5886 4302 5904 4320
rect 5886 4320 5904 4338
rect 5886 4338 5904 4356
rect 5886 4356 5904 4374
rect 5886 4374 5904 4392
rect 5886 4392 5904 4410
rect 5886 4410 5904 4428
rect 5886 4428 5904 4446
rect 5886 4446 5904 4464
rect 5886 4464 5904 4482
rect 5886 4482 5904 4500
rect 5886 4500 5904 4518
rect 5886 4518 5904 4536
rect 5886 4536 5904 4554
rect 5886 4554 5904 4572
rect 5886 4572 5904 4590
rect 5886 4590 5904 4608
rect 5886 4608 5904 4626
rect 5886 4626 5904 4644
rect 5886 4644 5904 4662
rect 5886 4662 5904 4680
rect 5886 4680 5904 4698
rect 5886 4698 5904 4716
rect 5886 4716 5904 4734
rect 5886 4734 5904 4752
rect 5886 4752 5904 4770
rect 5886 4770 5904 4788
rect 5886 4788 5904 4806
rect 5886 4806 5904 4824
rect 5886 4824 5904 4842
rect 5886 4842 5904 4860
rect 5886 4860 5904 4878
rect 5886 4878 5904 4896
rect 5886 4896 5904 4914
rect 5886 4914 5904 4932
rect 5886 4932 5904 4950
rect 5886 4950 5904 4968
rect 5886 4968 5904 4986
rect 5886 4986 5904 5004
rect 5886 5004 5904 5022
rect 5886 5022 5904 5040
rect 5886 5040 5904 5058
rect 5886 5058 5904 5076
rect 5886 5076 5904 5094
rect 5886 5094 5904 5112
rect 5886 5112 5904 5130
rect 5886 5130 5904 5148
rect 5886 5148 5904 5166
rect 5886 5166 5904 5184
rect 5886 5184 5904 5202
rect 5886 5202 5904 5220
rect 5886 5220 5904 5238
rect 5886 5238 5904 5256
rect 5886 5256 5904 5274
rect 5886 5526 5904 5544
rect 5886 5544 5904 5562
rect 5886 5562 5904 5580
rect 5886 5580 5904 5598
rect 5886 5598 5904 5616
rect 5886 5616 5904 5634
rect 5886 5634 5904 5652
rect 5886 5652 5904 5670
rect 5886 5670 5904 5688
rect 5886 5688 5904 5706
rect 5886 5706 5904 5724
rect 5886 5724 5904 5742
rect 5886 5742 5904 5760
rect 5886 5760 5904 5778
rect 5886 5778 5904 5796
rect 5886 5796 5904 5814
rect 5886 5814 5904 5832
rect 5886 5832 5904 5850
rect 5886 5850 5904 5868
rect 5886 5868 5904 5886
rect 5886 5886 5904 5904
rect 5886 5904 5904 5922
rect 5886 5922 5904 5940
rect 5886 5940 5904 5958
rect 5886 5958 5904 5976
rect 5886 5976 5904 5994
rect 5886 5994 5904 6012
rect 5886 6012 5904 6030
rect 5886 6030 5904 6048
rect 5886 6048 5904 6066
rect 5886 6066 5904 6084
rect 5886 6084 5904 6102
rect 5886 6102 5904 6120
rect 5886 6120 5904 6138
rect 5886 6138 5904 6156
rect 5886 6156 5904 6174
rect 5886 6174 5904 6192
rect 5886 6192 5904 6210
rect 5886 6210 5904 6228
rect 5886 6228 5904 6246
rect 5886 6246 5904 6264
rect 5886 6264 5904 6282
rect 5886 6282 5904 6300
rect 5886 6300 5904 6318
rect 5886 6318 5904 6336
rect 5886 6336 5904 6354
rect 5886 6354 5904 6372
rect 5886 6372 5904 6390
rect 5886 6390 5904 6408
rect 5886 6408 5904 6426
rect 5886 6426 5904 6444
rect 5886 6444 5904 6462
rect 5886 6462 5904 6480
rect 5886 6480 5904 6498
rect 5886 6498 5904 6516
rect 5886 6516 5904 6534
rect 5886 6534 5904 6552
rect 5886 6552 5904 6570
rect 5886 6570 5904 6588
rect 5886 6588 5904 6606
rect 5886 6606 5904 6624
rect 5886 6624 5904 6642
rect 5886 6642 5904 6660
rect 5886 6660 5904 6678
rect 5886 6678 5904 6696
rect 5886 6696 5904 6714
rect 5886 6714 5904 6732
rect 5886 6732 5904 6750
rect 5886 6750 5904 6768
rect 5886 6768 5904 6786
rect 5886 6786 5904 6804
rect 5886 6804 5904 6822
rect 5886 6822 5904 6840
rect 5886 6840 5904 6858
rect 5886 6858 5904 6876
rect 5886 6876 5904 6894
rect 5886 6894 5904 6912
rect 5886 6912 5904 6930
rect 5886 6930 5904 6948
rect 5886 6948 5904 6966
rect 5886 6966 5904 6984
rect 5886 6984 5904 7002
rect 5886 7002 5904 7020
rect 5886 7020 5904 7038
rect 5886 7038 5904 7056
rect 5886 7056 5904 7074
rect 5886 7074 5904 7092
rect 5886 7092 5904 7110
rect 5886 7110 5904 7128
rect 5886 7128 5904 7146
rect 5886 7146 5904 7164
rect 5886 7164 5904 7182
rect 5886 7182 5904 7200
rect 5886 7200 5904 7218
rect 5886 7218 5904 7236
rect 5886 7236 5904 7254
rect 5886 7254 5904 7272
rect 5886 7272 5904 7290
rect 5886 7290 5904 7308
rect 5886 7308 5904 7326
rect 5886 7326 5904 7344
rect 5886 7344 5904 7362
rect 5886 7362 5904 7380
rect 5886 7380 5904 7398
rect 5886 7398 5904 7416
rect 5886 7416 5904 7434
rect 5886 7434 5904 7452
rect 5886 7452 5904 7470
rect 5886 7470 5904 7488
rect 5886 7488 5904 7506
rect 5886 7506 5904 7524
rect 5886 7524 5904 7542
rect 5886 7542 5904 7560
rect 5886 7560 5904 7578
rect 5886 7578 5904 7596
rect 5886 7596 5904 7614
rect 5886 7614 5904 7632
rect 5886 7632 5904 7650
rect 5886 7650 5904 7668
rect 5886 7668 5904 7686
rect 5886 7686 5904 7704
rect 5886 7704 5904 7722
rect 5886 7722 5904 7740
rect 5886 7740 5904 7758
rect 5886 7758 5904 7776
rect 5886 7776 5904 7794
rect 5886 7794 5904 7812
rect 5886 7812 5904 7830
rect 5886 7830 5904 7848
rect 5886 7848 5904 7866
rect 5886 7866 5904 7884
rect 5886 7884 5904 7902
rect 5886 7902 5904 7920
rect 5886 7920 5904 7938
rect 5886 7938 5904 7956
rect 5886 7956 5904 7974
rect 5886 7974 5904 7992
rect 5886 7992 5904 8010
rect 5886 8010 5904 8028
rect 5886 8028 5904 8046
rect 5886 8046 5904 8064
rect 5886 8064 5904 8082
rect 5886 8082 5904 8100
rect 5886 8100 5904 8118
rect 5886 8118 5904 8136
rect 5886 8136 5904 8154
rect 5886 8154 5904 8172
rect 5886 8172 5904 8190
rect 5886 8190 5904 8208
rect 5886 8208 5904 8226
rect 5886 8226 5904 8244
rect 5886 8244 5904 8262
rect 5886 8262 5904 8280
rect 5886 8280 5904 8298
rect 5886 8298 5904 8316
rect 5886 8316 5904 8334
rect 5886 8334 5904 8352
rect 5886 8352 5904 8370
rect 5886 8370 5904 8388
rect 5886 8388 5904 8406
rect 5886 8406 5904 8424
rect 5886 8424 5904 8442
rect 5886 8442 5904 8460
rect 5886 8460 5904 8478
rect 5886 8478 5904 8496
rect 5886 8496 5904 8514
rect 5886 8514 5904 8532
rect 5886 8532 5904 8550
rect 5886 8550 5904 8568
rect 5886 8568 5904 8586
rect 5886 8586 5904 8604
rect 5886 8604 5904 8622
rect 5886 8622 5904 8640
rect 5886 8640 5904 8658
rect 5886 8658 5904 8676
rect 5886 8676 5904 8694
rect 5886 8694 5904 8712
rect 5886 8712 5904 8730
rect 5886 8730 5904 8748
rect 5886 8748 5904 8766
rect 5886 8766 5904 8784
rect 5886 8784 5904 8802
rect 5886 8802 5904 8820
rect 5886 8820 5904 8838
rect 5886 8838 5904 8856
rect 5886 8856 5904 8874
rect 5886 8874 5904 8892
rect 5886 8892 5904 8910
rect 5886 8910 5904 8928
rect 5886 8928 5904 8946
rect 5886 8946 5904 8964
rect 5886 8964 5904 8982
rect 5886 8982 5904 9000
rect 5886 9000 5904 9018
rect 5886 9018 5904 9036
rect 5886 9036 5904 9054
rect 5886 9054 5904 9072
rect 5886 9072 5904 9090
rect 5904 828 5922 846
rect 5904 846 5922 864
rect 5904 864 5922 882
rect 5904 882 5922 900
rect 5904 900 5922 918
rect 5904 918 5922 936
rect 5904 936 5922 954
rect 5904 954 5922 972
rect 5904 972 5922 990
rect 5904 990 5922 1008
rect 5904 1008 5922 1026
rect 5904 1026 5922 1044
rect 5904 1044 5922 1062
rect 5904 1224 5922 1242
rect 5904 1242 5922 1260
rect 5904 1260 5922 1278
rect 5904 1278 5922 1296
rect 5904 1296 5922 1314
rect 5904 1314 5922 1332
rect 5904 1332 5922 1350
rect 5904 1350 5922 1368
rect 5904 1368 5922 1386
rect 5904 1386 5922 1404
rect 5904 1404 5922 1422
rect 5904 1422 5922 1440
rect 5904 1440 5922 1458
rect 5904 1458 5922 1476
rect 5904 1476 5922 1494
rect 5904 1494 5922 1512
rect 5904 1512 5922 1530
rect 5904 1530 5922 1548
rect 5904 1548 5922 1566
rect 5904 1566 5922 1584
rect 5904 1584 5922 1602
rect 5904 1602 5922 1620
rect 5904 1620 5922 1638
rect 5904 1638 5922 1656
rect 5904 1656 5922 1674
rect 5904 1674 5922 1692
rect 5904 1692 5922 1710
rect 5904 1710 5922 1728
rect 5904 1728 5922 1746
rect 5904 1746 5922 1764
rect 5904 1764 5922 1782
rect 5904 1782 5922 1800
rect 5904 1800 5922 1818
rect 5904 1818 5922 1836
rect 5904 1836 5922 1854
rect 5904 1854 5922 1872
rect 5904 1872 5922 1890
rect 5904 1890 5922 1908
rect 5904 1908 5922 1926
rect 5904 1926 5922 1944
rect 5904 1944 5922 1962
rect 5904 1962 5922 1980
rect 5904 1980 5922 1998
rect 5904 1998 5922 2016
rect 5904 2016 5922 2034
rect 5904 2034 5922 2052
rect 5904 2052 5922 2070
rect 5904 2070 5922 2088
rect 5904 2088 5922 2106
rect 5904 2106 5922 2124
rect 5904 2124 5922 2142
rect 5904 2142 5922 2160
rect 5904 2160 5922 2178
rect 5904 2178 5922 2196
rect 5904 2196 5922 2214
rect 5904 2214 5922 2232
rect 5904 2232 5922 2250
rect 5904 2250 5922 2268
rect 5904 2268 5922 2286
rect 5904 2286 5922 2304
rect 5904 2304 5922 2322
rect 5904 2322 5922 2340
rect 5904 2340 5922 2358
rect 5904 2358 5922 2376
rect 5904 2376 5922 2394
rect 5904 2394 5922 2412
rect 5904 2412 5922 2430
rect 5904 2430 5922 2448
rect 5904 2448 5922 2466
rect 5904 2466 5922 2484
rect 5904 2484 5922 2502
rect 5904 2502 5922 2520
rect 5904 2520 5922 2538
rect 5904 2538 5922 2556
rect 5904 2556 5922 2574
rect 5904 2574 5922 2592
rect 5904 2592 5922 2610
rect 5904 2610 5922 2628
rect 5904 2628 5922 2646
rect 5904 2646 5922 2664
rect 5904 2664 5922 2682
rect 5904 2682 5922 2700
rect 5904 2700 5922 2718
rect 5904 2934 5922 2952
rect 5904 2952 5922 2970
rect 5904 2970 5922 2988
rect 5904 2988 5922 3006
rect 5904 3006 5922 3024
rect 5904 3024 5922 3042
rect 5904 3042 5922 3060
rect 5904 3060 5922 3078
rect 5904 3078 5922 3096
rect 5904 3096 5922 3114
rect 5904 3114 5922 3132
rect 5904 3132 5922 3150
rect 5904 3150 5922 3168
rect 5904 3168 5922 3186
rect 5904 3186 5922 3204
rect 5904 3204 5922 3222
rect 5904 3222 5922 3240
rect 5904 3240 5922 3258
rect 5904 3258 5922 3276
rect 5904 3276 5922 3294
rect 5904 3294 5922 3312
rect 5904 3312 5922 3330
rect 5904 3330 5922 3348
rect 5904 3348 5922 3366
rect 5904 3366 5922 3384
rect 5904 3384 5922 3402
rect 5904 3402 5922 3420
rect 5904 3420 5922 3438
rect 5904 3438 5922 3456
rect 5904 3456 5922 3474
rect 5904 3474 5922 3492
rect 5904 3492 5922 3510
rect 5904 3510 5922 3528
rect 5904 3528 5922 3546
rect 5904 3546 5922 3564
rect 5904 3564 5922 3582
rect 5904 3582 5922 3600
rect 5904 3600 5922 3618
rect 5904 3618 5922 3636
rect 5904 3636 5922 3654
rect 5904 3654 5922 3672
rect 5904 3672 5922 3690
rect 5904 3690 5922 3708
rect 5904 3708 5922 3726
rect 5904 3726 5922 3744
rect 5904 3744 5922 3762
rect 5904 3762 5922 3780
rect 5904 3780 5922 3798
rect 5904 3798 5922 3816
rect 5904 3816 5922 3834
rect 5904 3834 5922 3852
rect 5904 3852 5922 3870
rect 5904 3870 5922 3888
rect 5904 3888 5922 3906
rect 5904 3906 5922 3924
rect 5904 3924 5922 3942
rect 5904 3942 5922 3960
rect 5904 3960 5922 3978
rect 5904 3978 5922 3996
rect 5904 3996 5922 4014
rect 5904 4014 5922 4032
rect 5904 4032 5922 4050
rect 5904 4050 5922 4068
rect 5904 4068 5922 4086
rect 5904 4086 5922 4104
rect 5904 4104 5922 4122
rect 5904 4122 5922 4140
rect 5904 4140 5922 4158
rect 5904 4158 5922 4176
rect 5904 4176 5922 4194
rect 5904 4194 5922 4212
rect 5904 4212 5922 4230
rect 5904 4230 5922 4248
rect 5904 4248 5922 4266
rect 5904 4266 5922 4284
rect 5904 4284 5922 4302
rect 5904 4302 5922 4320
rect 5904 4320 5922 4338
rect 5904 4338 5922 4356
rect 5904 4356 5922 4374
rect 5904 4374 5922 4392
rect 5904 4392 5922 4410
rect 5904 4410 5922 4428
rect 5904 4428 5922 4446
rect 5904 4446 5922 4464
rect 5904 4464 5922 4482
rect 5904 4482 5922 4500
rect 5904 4500 5922 4518
rect 5904 4518 5922 4536
rect 5904 4536 5922 4554
rect 5904 4554 5922 4572
rect 5904 4572 5922 4590
rect 5904 4590 5922 4608
rect 5904 4608 5922 4626
rect 5904 4626 5922 4644
rect 5904 4644 5922 4662
rect 5904 4662 5922 4680
rect 5904 4680 5922 4698
rect 5904 4698 5922 4716
rect 5904 4716 5922 4734
rect 5904 4734 5922 4752
rect 5904 4752 5922 4770
rect 5904 4770 5922 4788
rect 5904 4788 5922 4806
rect 5904 4806 5922 4824
rect 5904 4824 5922 4842
rect 5904 4842 5922 4860
rect 5904 4860 5922 4878
rect 5904 4878 5922 4896
rect 5904 4896 5922 4914
rect 5904 4914 5922 4932
rect 5904 4932 5922 4950
rect 5904 4950 5922 4968
rect 5904 4968 5922 4986
rect 5904 4986 5922 5004
rect 5904 5004 5922 5022
rect 5904 5022 5922 5040
rect 5904 5040 5922 5058
rect 5904 5058 5922 5076
rect 5904 5076 5922 5094
rect 5904 5094 5922 5112
rect 5904 5112 5922 5130
rect 5904 5130 5922 5148
rect 5904 5148 5922 5166
rect 5904 5166 5922 5184
rect 5904 5184 5922 5202
rect 5904 5202 5922 5220
rect 5904 5220 5922 5238
rect 5904 5238 5922 5256
rect 5904 5256 5922 5274
rect 5904 5274 5922 5292
rect 5904 5544 5922 5562
rect 5904 5562 5922 5580
rect 5904 5580 5922 5598
rect 5904 5598 5922 5616
rect 5904 5616 5922 5634
rect 5904 5634 5922 5652
rect 5904 5652 5922 5670
rect 5904 5670 5922 5688
rect 5904 5688 5922 5706
rect 5904 5706 5922 5724
rect 5904 5724 5922 5742
rect 5904 5742 5922 5760
rect 5904 5760 5922 5778
rect 5904 5778 5922 5796
rect 5904 5796 5922 5814
rect 5904 5814 5922 5832
rect 5904 5832 5922 5850
rect 5904 5850 5922 5868
rect 5904 5868 5922 5886
rect 5904 5886 5922 5904
rect 5904 5904 5922 5922
rect 5904 5922 5922 5940
rect 5904 5940 5922 5958
rect 5904 5958 5922 5976
rect 5904 5976 5922 5994
rect 5904 5994 5922 6012
rect 5904 6012 5922 6030
rect 5904 6030 5922 6048
rect 5904 6048 5922 6066
rect 5904 6066 5922 6084
rect 5904 6084 5922 6102
rect 5904 6102 5922 6120
rect 5904 6120 5922 6138
rect 5904 6138 5922 6156
rect 5904 6156 5922 6174
rect 5904 6174 5922 6192
rect 5904 6192 5922 6210
rect 5904 6210 5922 6228
rect 5904 6228 5922 6246
rect 5904 6246 5922 6264
rect 5904 6264 5922 6282
rect 5904 6282 5922 6300
rect 5904 6300 5922 6318
rect 5904 6318 5922 6336
rect 5904 6336 5922 6354
rect 5904 6354 5922 6372
rect 5904 6372 5922 6390
rect 5904 6390 5922 6408
rect 5904 6408 5922 6426
rect 5904 6426 5922 6444
rect 5904 6444 5922 6462
rect 5904 6462 5922 6480
rect 5904 6480 5922 6498
rect 5904 6498 5922 6516
rect 5904 6516 5922 6534
rect 5904 6534 5922 6552
rect 5904 6552 5922 6570
rect 5904 6570 5922 6588
rect 5904 6588 5922 6606
rect 5904 6606 5922 6624
rect 5904 6624 5922 6642
rect 5904 6642 5922 6660
rect 5904 6660 5922 6678
rect 5904 6678 5922 6696
rect 5904 6696 5922 6714
rect 5904 6714 5922 6732
rect 5904 6732 5922 6750
rect 5904 6750 5922 6768
rect 5904 6768 5922 6786
rect 5904 6786 5922 6804
rect 5904 6804 5922 6822
rect 5904 6822 5922 6840
rect 5904 6840 5922 6858
rect 5904 6858 5922 6876
rect 5904 6876 5922 6894
rect 5904 6894 5922 6912
rect 5904 6912 5922 6930
rect 5904 6930 5922 6948
rect 5904 6948 5922 6966
rect 5904 6966 5922 6984
rect 5904 6984 5922 7002
rect 5904 7002 5922 7020
rect 5904 7020 5922 7038
rect 5904 7038 5922 7056
rect 5904 7056 5922 7074
rect 5904 7074 5922 7092
rect 5904 7092 5922 7110
rect 5904 7110 5922 7128
rect 5904 7128 5922 7146
rect 5904 7146 5922 7164
rect 5904 7164 5922 7182
rect 5904 7182 5922 7200
rect 5904 7200 5922 7218
rect 5904 7218 5922 7236
rect 5904 7236 5922 7254
rect 5904 7254 5922 7272
rect 5904 7272 5922 7290
rect 5904 7290 5922 7308
rect 5904 7308 5922 7326
rect 5904 7326 5922 7344
rect 5904 7344 5922 7362
rect 5904 7362 5922 7380
rect 5904 7380 5922 7398
rect 5904 7398 5922 7416
rect 5904 7416 5922 7434
rect 5904 7434 5922 7452
rect 5904 7452 5922 7470
rect 5904 7470 5922 7488
rect 5904 7488 5922 7506
rect 5904 7506 5922 7524
rect 5904 7524 5922 7542
rect 5904 7542 5922 7560
rect 5904 7560 5922 7578
rect 5904 7578 5922 7596
rect 5904 7596 5922 7614
rect 5904 7614 5922 7632
rect 5904 7632 5922 7650
rect 5904 7650 5922 7668
rect 5904 7668 5922 7686
rect 5904 7686 5922 7704
rect 5904 7704 5922 7722
rect 5904 7722 5922 7740
rect 5904 7740 5922 7758
rect 5904 7758 5922 7776
rect 5904 7776 5922 7794
rect 5904 7794 5922 7812
rect 5904 7812 5922 7830
rect 5904 7830 5922 7848
rect 5904 7848 5922 7866
rect 5904 7866 5922 7884
rect 5904 7884 5922 7902
rect 5904 7902 5922 7920
rect 5904 7920 5922 7938
rect 5904 7938 5922 7956
rect 5904 7956 5922 7974
rect 5904 7974 5922 7992
rect 5904 7992 5922 8010
rect 5904 8010 5922 8028
rect 5904 8028 5922 8046
rect 5904 8046 5922 8064
rect 5904 8064 5922 8082
rect 5904 8082 5922 8100
rect 5904 8100 5922 8118
rect 5904 8118 5922 8136
rect 5904 8136 5922 8154
rect 5904 8154 5922 8172
rect 5904 8172 5922 8190
rect 5904 8190 5922 8208
rect 5904 8208 5922 8226
rect 5904 8226 5922 8244
rect 5904 8244 5922 8262
rect 5904 8262 5922 8280
rect 5904 8280 5922 8298
rect 5904 8298 5922 8316
rect 5904 8316 5922 8334
rect 5904 8334 5922 8352
rect 5904 8352 5922 8370
rect 5904 8370 5922 8388
rect 5904 8388 5922 8406
rect 5904 8406 5922 8424
rect 5904 8424 5922 8442
rect 5904 8442 5922 8460
rect 5904 8460 5922 8478
rect 5904 8478 5922 8496
rect 5904 8496 5922 8514
rect 5904 8514 5922 8532
rect 5904 8532 5922 8550
rect 5904 8550 5922 8568
rect 5904 8568 5922 8586
rect 5904 8586 5922 8604
rect 5904 8604 5922 8622
rect 5904 8622 5922 8640
rect 5904 8640 5922 8658
rect 5904 8658 5922 8676
rect 5904 8676 5922 8694
rect 5904 8694 5922 8712
rect 5904 8712 5922 8730
rect 5904 8730 5922 8748
rect 5904 8748 5922 8766
rect 5904 8766 5922 8784
rect 5904 8784 5922 8802
rect 5904 8802 5922 8820
rect 5904 8820 5922 8838
rect 5904 8838 5922 8856
rect 5904 8856 5922 8874
rect 5904 8874 5922 8892
rect 5904 8892 5922 8910
rect 5904 8910 5922 8928
rect 5904 8928 5922 8946
rect 5904 8946 5922 8964
rect 5904 8964 5922 8982
rect 5904 8982 5922 9000
rect 5904 9000 5922 9018
rect 5904 9018 5922 9036
rect 5904 9036 5922 9054
rect 5904 9054 5922 9072
rect 5904 9072 5922 9090
rect 5904 9090 5922 9108
rect 5922 846 5940 864
rect 5922 864 5940 882
rect 5922 882 5940 900
rect 5922 900 5940 918
rect 5922 918 5940 936
rect 5922 936 5940 954
rect 5922 954 5940 972
rect 5922 972 5940 990
rect 5922 990 5940 1008
rect 5922 1008 5940 1026
rect 5922 1026 5940 1044
rect 5922 1044 5940 1062
rect 5922 1062 5940 1080
rect 5922 1224 5940 1242
rect 5922 1242 5940 1260
rect 5922 1260 5940 1278
rect 5922 1278 5940 1296
rect 5922 1296 5940 1314
rect 5922 1314 5940 1332
rect 5922 1332 5940 1350
rect 5922 1350 5940 1368
rect 5922 1368 5940 1386
rect 5922 1386 5940 1404
rect 5922 1404 5940 1422
rect 5922 1422 5940 1440
rect 5922 1440 5940 1458
rect 5922 1458 5940 1476
rect 5922 1476 5940 1494
rect 5922 1494 5940 1512
rect 5922 1512 5940 1530
rect 5922 1530 5940 1548
rect 5922 1548 5940 1566
rect 5922 1566 5940 1584
rect 5922 1584 5940 1602
rect 5922 1602 5940 1620
rect 5922 1620 5940 1638
rect 5922 1638 5940 1656
rect 5922 1656 5940 1674
rect 5922 1674 5940 1692
rect 5922 1692 5940 1710
rect 5922 1710 5940 1728
rect 5922 1728 5940 1746
rect 5922 1746 5940 1764
rect 5922 1764 5940 1782
rect 5922 1782 5940 1800
rect 5922 1800 5940 1818
rect 5922 1818 5940 1836
rect 5922 1836 5940 1854
rect 5922 1854 5940 1872
rect 5922 1872 5940 1890
rect 5922 1890 5940 1908
rect 5922 1908 5940 1926
rect 5922 1926 5940 1944
rect 5922 1944 5940 1962
rect 5922 1962 5940 1980
rect 5922 1980 5940 1998
rect 5922 1998 5940 2016
rect 5922 2016 5940 2034
rect 5922 2034 5940 2052
rect 5922 2052 5940 2070
rect 5922 2070 5940 2088
rect 5922 2088 5940 2106
rect 5922 2106 5940 2124
rect 5922 2124 5940 2142
rect 5922 2142 5940 2160
rect 5922 2160 5940 2178
rect 5922 2178 5940 2196
rect 5922 2196 5940 2214
rect 5922 2214 5940 2232
rect 5922 2232 5940 2250
rect 5922 2250 5940 2268
rect 5922 2268 5940 2286
rect 5922 2286 5940 2304
rect 5922 2304 5940 2322
rect 5922 2322 5940 2340
rect 5922 2340 5940 2358
rect 5922 2358 5940 2376
rect 5922 2376 5940 2394
rect 5922 2394 5940 2412
rect 5922 2412 5940 2430
rect 5922 2430 5940 2448
rect 5922 2448 5940 2466
rect 5922 2466 5940 2484
rect 5922 2484 5940 2502
rect 5922 2502 5940 2520
rect 5922 2520 5940 2538
rect 5922 2538 5940 2556
rect 5922 2556 5940 2574
rect 5922 2574 5940 2592
rect 5922 2592 5940 2610
rect 5922 2610 5940 2628
rect 5922 2628 5940 2646
rect 5922 2646 5940 2664
rect 5922 2664 5940 2682
rect 5922 2682 5940 2700
rect 5922 2700 5940 2718
rect 5922 2952 5940 2970
rect 5922 2970 5940 2988
rect 5922 2988 5940 3006
rect 5922 3006 5940 3024
rect 5922 3024 5940 3042
rect 5922 3042 5940 3060
rect 5922 3060 5940 3078
rect 5922 3078 5940 3096
rect 5922 3096 5940 3114
rect 5922 3114 5940 3132
rect 5922 3132 5940 3150
rect 5922 3150 5940 3168
rect 5922 3168 5940 3186
rect 5922 3186 5940 3204
rect 5922 3204 5940 3222
rect 5922 3222 5940 3240
rect 5922 3240 5940 3258
rect 5922 3258 5940 3276
rect 5922 3276 5940 3294
rect 5922 3294 5940 3312
rect 5922 3312 5940 3330
rect 5922 3330 5940 3348
rect 5922 3348 5940 3366
rect 5922 3366 5940 3384
rect 5922 3384 5940 3402
rect 5922 3402 5940 3420
rect 5922 3420 5940 3438
rect 5922 3438 5940 3456
rect 5922 3456 5940 3474
rect 5922 3474 5940 3492
rect 5922 3492 5940 3510
rect 5922 3510 5940 3528
rect 5922 3528 5940 3546
rect 5922 3546 5940 3564
rect 5922 3564 5940 3582
rect 5922 3582 5940 3600
rect 5922 3600 5940 3618
rect 5922 3618 5940 3636
rect 5922 3636 5940 3654
rect 5922 3654 5940 3672
rect 5922 3672 5940 3690
rect 5922 3690 5940 3708
rect 5922 3708 5940 3726
rect 5922 3726 5940 3744
rect 5922 3744 5940 3762
rect 5922 3762 5940 3780
rect 5922 3780 5940 3798
rect 5922 3798 5940 3816
rect 5922 3816 5940 3834
rect 5922 3834 5940 3852
rect 5922 3852 5940 3870
rect 5922 3870 5940 3888
rect 5922 3888 5940 3906
rect 5922 3906 5940 3924
rect 5922 3924 5940 3942
rect 5922 3942 5940 3960
rect 5922 3960 5940 3978
rect 5922 3978 5940 3996
rect 5922 3996 5940 4014
rect 5922 4014 5940 4032
rect 5922 4032 5940 4050
rect 5922 4050 5940 4068
rect 5922 4068 5940 4086
rect 5922 4086 5940 4104
rect 5922 4104 5940 4122
rect 5922 4122 5940 4140
rect 5922 4140 5940 4158
rect 5922 4158 5940 4176
rect 5922 4176 5940 4194
rect 5922 4194 5940 4212
rect 5922 4212 5940 4230
rect 5922 4230 5940 4248
rect 5922 4248 5940 4266
rect 5922 4266 5940 4284
rect 5922 4284 5940 4302
rect 5922 4302 5940 4320
rect 5922 4320 5940 4338
rect 5922 4338 5940 4356
rect 5922 4356 5940 4374
rect 5922 4374 5940 4392
rect 5922 4392 5940 4410
rect 5922 4410 5940 4428
rect 5922 4428 5940 4446
rect 5922 4446 5940 4464
rect 5922 4464 5940 4482
rect 5922 4482 5940 4500
rect 5922 4500 5940 4518
rect 5922 4518 5940 4536
rect 5922 4536 5940 4554
rect 5922 4554 5940 4572
rect 5922 4572 5940 4590
rect 5922 4590 5940 4608
rect 5922 4608 5940 4626
rect 5922 4626 5940 4644
rect 5922 4644 5940 4662
rect 5922 4662 5940 4680
rect 5922 4680 5940 4698
rect 5922 4698 5940 4716
rect 5922 4716 5940 4734
rect 5922 4734 5940 4752
rect 5922 4752 5940 4770
rect 5922 4770 5940 4788
rect 5922 4788 5940 4806
rect 5922 4806 5940 4824
rect 5922 4824 5940 4842
rect 5922 4842 5940 4860
rect 5922 4860 5940 4878
rect 5922 4878 5940 4896
rect 5922 4896 5940 4914
rect 5922 4914 5940 4932
rect 5922 4932 5940 4950
rect 5922 4950 5940 4968
rect 5922 4968 5940 4986
rect 5922 4986 5940 5004
rect 5922 5004 5940 5022
rect 5922 5022 5940 5040
rect 5922 5040 5940 5058
rect 5922 5058 5940 5076
rect 5922 5076 5940 5094
rect 5922 5094 5940 5112
rect 5922 5112 5940 5130
rect 5922 5130 5940 5148
rect 5922 5148 5940 5166
rect 5922 5166 5940 5184
rect 5922 5184 5940 5202
rect 5922 5202 5940 5220
rect 5922 5220 5940 5238
rect 5922 5238 5940 5256
rect 5922 5256 5940 5274
rect 5922 5274 5940 5292
rect 5922 5292 5940 5310
rect 5922 5562 5940 5580
rect 5922 5580 5940 5598
rect 5922 5598 5940 5616
rect 5922 5616 5940 5634
rect 5922 5634 5940 5652
rect 5922 5652 5940 5670
rect 5922 5670 5940 5688
rect 5922 5688 5940 5706
rect 5922 5706 5940 5724
rect 5922 5724 5940 5742
rect 5922 5742 5940 5760
rect 5922 5760 5940 5778
rect 5922 5778 5940 5796
rect 5922 5796 5940 5814
rect 5922 5814 5940 5832
rect 5922 5832 5940 5850
rect 5922 5850 5940 5868
rect 5922 5868 5940 5886
rect 5922 5886 5940 5904
rect 5922 5904 5940 5922
rect 5922 5922 5940 5940
rect 5922 5940 5940 5958
rect 5922 5958 5940 5976
rect 5922 5976 5940 5994
rect 5922 5994 5940 6012
rect 5922 6012 5940 6030
rect 5922 6030 5940 6048
rect 5922 6048 5940 6066
rect 5922 6066 5940 6084
rect 5922 6084 5940 6102
rect 5922 6102 5940 6120
rect 5922 6120 5940 6138
rect 5922 6138 5940 6156
rect 5922 6156 5940 6174
rect 5922 6174 5940 6192
rect 5922 6192 5940 6210
rect 5922 6210 5940 6228
rect 5922 6228 5940 6246
rect 5922 6246 5940 6264
rect 5922 6264 5940 6282
rect 5922 6282 5940 6300
rect 5922 6300 5940 6318
rect 5922 6318 5940 6336
rect 5922 6336 5940 6354
rect 5922 6354 5940 6372
rect 5922 6372 5940 6390
rect 5922 6390 5940 6408
rect 5922 6408 5940 6426
rect 5922 6426 5940 6444
rect 5922 6444 5940 6462
rect 5922 6462 5940 6480
rect 5922 6480 5940 6498
rect 5922 6498 5940 6516
rect 5922 6516 5940 6534
rect 5922 6534 5940 6552
rect 5922 6552 5940 6570
rect 5922 6570 5940 6588
rect 5922 6588 5940 6606
rect 5922 6606 5940 6624
rect 5922 6624 5940 6642
rect 5922 6642 5940 6660
rect 5922 6660 5940 6678
rect 5922 6678 5940 6696
rect 5922 6696 5940 6714
rect 5922 6714 5940 6732
rect 5922 6732 5940 6750
rect 5922 6750 5940 6768
rect 5922 6768 5940 6786
rect 5922 6786 5940 6804
rect 5922 6804 5940 6822
rect 5922 6822 5940 6840
rect 5922 6840 5940 6858
rect 5922 6858 5940 6876
rect 5922 6876 5940 6894
rect 5922 6894 5940 6912
rect 5922 6912 5940 6930
rect 5922 6930 5940 6948
rect 5922 6948 5940 6966
rect 5922 6966 5940 6984
rect 5922 6984 5940 7002
rect 5922 7002 5940 7020
rect 5922 7020 5940 7038
rect 5922 7038 5940 7056
rect 5922 7056 5940 7074
rect 5922 7074 5940 7092
rect 5922 7092 5940 7110
rect 5922 7110 5940 7128
rect 5922 7128 5940 7146
rect 5922 7146 5940 7164
rect 5922 7164 5940 7182
rect 5922 7182 5940 7200
rect 5922 7200 5940 7218
rect 5922 7218 5940 7236
rect 5922 7236 5940 7254
rect 5922 7254 5940 7272
rect 5922 7272 5940 7290
rect 5922 7290 5940 7308
rect 5922 7308 5940 7326
rect 5922 7326 5940 7344
rect 5922 7344 5940 7362
rect 5922 7362 5940 7380
rect 5922 7380 5940 7398
rect 5922 7398 5940 7416
rect 5922 7416 5940 7434
rect 5922 7434 5940 7452
rect 5922 7452 5940 7470
rect 5922 7470 5940 7488
rect 5922 7488 5940 7506
rect 5922 7506 5940 7524
rect 5922 7524 5940 7542
rect 5922 7542 5940 7560
rect 5922 7560 5940 7578
rect 5922 7578 5940 7596
rect 5922 7596 5940 7614
rect 5922 7614 5940 7632
rect 5922 7632 5940 7650
rect 5922 7650 5940 7668
rect 5922 7668 5940 7686
rect 5922 7686 5940 7704
rect 5922 7704 5940 7722
rect 5922 7722 5940 7740
rect 5922 7740 5940 7758
rect 5922 7758 5940 7776
rect 5922 7776 5940 7794
rect 5922 7794 5940 7812
rect 5922 7812 5940 7830
rect 5922 7830 5940 7848
rect 5922 7848 5940 7866
rect 5922 7866 5940 7884
rect 5922 7884 5940 7902
rect 5922 7902 5940 7920
rect 5922 7920 5940 7938
rect 5922 7938 5940 7956
rect 5922 7956 5940 7974
rect 5922 7974 5940 7992
rect 5922 7992 5940 8010
rect 5922 8010 5940 8028
rect 5922 8028 5940 8046
rect 5922 8046 5940 8064
rect 5922 8064 5940 8082
rect 5922 8082 5940 8100
rect 5922 8100 5940 8118
rect 5922 8118 5940 8136
rect 5922 8136 5940 8154
rect 5922 8154 5940 8172
rect 5922 8172 5940 8190
rect 5922 8190 5940 8208
rect 5922 8208 5940 8226
rect 5922 8226 5940 8244
rect 5922 8244 5940 8262
rect 5922 8262 5940 8280
rect 5922 8280 5940 8298
rect 5922 8298 5940 8316
rect 5922 8316 5940 8334
rect 5922 8334 5940 8352
rect 5922 8352 5940 8370
rect 5922 8370 5940 8388
rect 5922 8388 5940 8406
rect 5922 8406 5940 8424
rect 5922 8424 5940 8442
rect 5922 8442 5940 8460
rect 5922 8460 5940 8478
rect 5922 8478 5940 8496
rect 5922 8496 5940 8514
rect 5922 8514 5940 8532
rect 5922 8532 5940 8550
rect 5922 8550 5940 8568
rect 5922 8568 5940 8586
rect 5922 8586 5940 8604
rect 5922 8604 5940 8622
rect 5922 8622 5940 8640
rect 5922 8640 5940 8658
rect 5922 8658 5940 8676
rect 5922 8676 5940 8694
rect 5922 8694 5940 8712
rect 5922 8712 5940 8730
rect 5922 8730 5940 8748
rect 5922 8748 5940 8766
rect 5922 8766 5940 8784
rect 5922 8784 5940 8802
rect 5922 8802 5940 8820
rect 5922 8820 5940 8838
rect 5922 8838 5940 8856
rect 5922 8856 5940 8874
rect 5922 8874 5940 8892
rect 5922 8892 5940 8910
rect 5922 8910 5940 8928
rect 5922 8928 5940 8946
rect 5922 8946 5940 8964
rect 5922 8964 5940 8982
rect 5922 8982 5940 9000
rect 5922 9000 5940 9018
rect 5922 9018 5940 9036
rect 5922 9036 5940 9054
rect 5922 9054 5940 9072
rect 5922 9072 5940 9090
rect 5922 9090 5940 9108
rect 5922 9108 5940 9126
rect 5940 864 5958 882
rect 5940 882 5958 900
rect 5940 900 5958 918
rect 5940 918 5958 936
rect 5940 936 5958 954
rect 5940 954 5958 972
rect 5940 972 5958 990
rect 5940 990 5958 1008
rect 5940 1008 5958 1026
rect 5940 1026 5958 1044
rect 5940 1044 5958 1062
rect 5940 1062 5958 1080
rect 5940 1224 5958 1242
rect 5940 1242 5958 1260
rect 5940 1260 5958 1278
rect 5940 1278 5958 1296
rect 5940 1296 5958 1314
rect 5940 1314 5958 1332
rect 5940 1332 5958 1350
rect 5940 1350 5958 1368
rect 5940 1368 5958 1386
rect 5940 1386 5958 1404
rect 5940 1404 5958 1422
rect 5940 1422 5958 1440
rect 5940 1440 5958 1458
rect 5940 1458 5958 1476
rect 5940 1476 5958 1494
rect 5940 1494 5958 1512
rect 5940 1512 5958 1530
rect 5940 1530 5958 1548
rect 5940 1548 5958 1566
rect 5940 1566 5958 1584
rect 5940 1584 5958 1602
rect 5940 1602 5958 1620
rect 5940 1620 5958 1638
rect 5940 1638 5958 1656
rect 5940 1656 5958 1674
rect 5940 1674 5958 1692
rect 5940 1692 5958 1710
rect 5940 1710 5958 1728
rect 5940 1728 5958 1746
rect 5940 1746 5958 1764
rect 5940 1764 5958 1782
rect 5940 1782 5958 1800
rect 5940 1800 5958 1818
rect 5940 1818 5958 1836
rect 5940 1836 5958 1854
rect 5940 1854 5958 1872
rect 5940 1872 5958 1890
rect 5940 1890 5958 1908
rect 5940 1908 5958 1926
rect 5940 1926 5958 1944
rect 5940 1944 5958 1962
rect 5940 1962 5958 1980
rect 5940 1980 5958 1998
rect 5940 1998 5958 2016
rect 5940 2016 5958 2034
rect 5940 2034 5958 2052
rect 5940 2052 5958 2070
rect 5940 2070 5958 2088
rect 5940 2088 5958 2106
rect 5940 2106 5958 2124
rect 5940 2124 5958 2142
rect 5940 2142 5958 2160
rect 5940 2160 5958 2178
rect 5940 2178 5958 2196
rect 5940 2196 5958 2214
rect 5940 2214 5958 2232
rect 5940 2232 5958 2250
rect 5940 2250 5958 2268
rect 5940 2268 5958 2286
rect 5940 2286 5958 2304
rect 5940 2304 5958 2322
rect 5940 2322 5958 2340
rect 5940 2340 5958 2358
rect 5940 2358 5958 2376
rect 5940 2376 5958 2394
rect 5940 2394 5958 2412
rect 5940 2412 5958 2430
rect 5940 2430 5958 2448
rect 5940 2448 5958 2466
rect 5940 2466 5958 2484
rect 5940 2484 5958 2502
rect 5940 2502 5958 2520
rect 5940 2520 5958 2538
rect 5940 2538 5958 2556
rect 5940 2556 5958 2574
rect 5940 2574 5958 2592
rect 5940 2592 5958 2610
rect 5940 2610 5958 2628
rect 5940 2628 5958 2646
rect 5940 2646 5958 2664
rect 5940 2664 5958 2682
rect 5940 2682 5958 2700
rect 5940 2700 5958 2718
rect 5940 2952 5958 2970
rect 5940 2970 5958 2988
rect 5940 2988 5958 3006
rect 5940 3006 5958 3024
rect 5940 3024 5958 3042
rect 5940 3042 5958 3060
rect 5940 3060 5958 3078
rect 5940 3078 5958 3096
rect 5940 3096 5958 3114
rect 5940 3114 5958 3132
rect 5940 3132 5958 3150
rect 5940 3150 5958 3168
rect 5940 3168 5958 3186
rect 5940 3186 5958 3204
rect 5940 3204 5958 3222
rect 5940 3222 5958 3240
rect 5940 3240 5958 3258
rect 5940 3258 5958 3276
rect 5940 3276 5958 3294
rect 5940 3294 5958 3312
rect 5940 3312 5958 3330
rect 5940 3330 5958 3348
rect 5940 3348 5958 3366
rect 5940 3366 5958 3384
rect 5940 3384 5958 3402
rect 5940 3402 5958 3420
rect 5940 3420 5958 3438
rect 5940 3438 5958 3456
rect 5940 3456 5958 3474
rect 5940 3474 5958 3492
rect 5940 3492 5958 3510
rect 5940 3510 5958 3528
rect 5940 3528 5958 3546
rect 5940 3546 5958 3564
rect 5940 3564 5958 3582
rect 5940 3582 5958 3600
rect 5940 3600 5958 3618
rect 5940 3618 5958 3636
rect 5940 3636 5958 3654
rect 5940 3654 5958 3672
rect 5940 3672 5958 3690
rect 5940 3690 5958 3708
rect 5940 3708 5958 3726
rect 5940 3726 5958 3744
rect 5940 3744 5958 3762
rect 5940 3762 5958 3780
rect 5940 3780 5958 3798
rect 5940 3798 5958 3816
rect 5940 3816 5958 3834
rect 5940 3834 5958 3852
rect 5940 3852 5958 3870
rect 5940 3870 5958 3888
rect 5940 3888 5958 3906
rect 5940 3906 5958 3924
rect 5940 3924 5958 3942
rect 5940 3942 5958 3960
rect 5940 3960 5958 3978
rect 5940 3978 5958 3996
rect 5940 3996 5958 4014
rect 5940 4014 5958 4032
rect 5940 4032 5958 4050
rect 5940 4050 5958 4068
rect 5940 4068 5958 4086
rect 5940 4086 5958 4104
rect 5940 4104 5958 4122
rect 5940 4122 5958 4140
rect 5940 4140 5958 4158
rect 5940 4158 5958 4176
rect 5940 4176 5958 4194
rect 5940 4194 5958 4212
rect 5940 4212 5958 4230
rect 5940 4230 5958 4248
rect 5940 4248 5958 4266
rect 5940 4266 5958 4284
rect 5940 4284 5958 4302
rect 5940 4302 5958 4320
rect 5940 4320 5958 4338
rect 5940 4338 5958 4356
rect 5940 4356 5958 4374
rect 5940 4374 5958 4392
rect 5940 4392 5958 4410
rect 5940 4410 5958 4428
rect 5940 4428 5958 4446
rect 5940 4446 5958 4464
rect 5940 4464 5958 4482
rect 5940 4482 5958 4500
rect 5940 4500 5958 4518
rect 5940 4518 5958 4536
rect 5940 4536 5958 4554
rect 5940 4554 5958 4572
rect 5940 4572 5958 4590
rect 5940 4590 5958 4608
rect 5940 4608 5958 4626
rect 5940 4626 5958 4644
rect 5940 4644 5958 4662
rect 5940 4662 5958 4680
rect 5940 4680 5958 4698
rect 5940 4698 5958 4716
rect 5940 4716 5958 4734
rect 5940 4734 5958 4752
rect 5940 4752 5958 4770
rect 5940 4770 5958 4788
rect 5940 4788 5958 4806
rect 5940 4806 5958 4824
rect 5940 4824 5958 4842
rect 5940 4842 5958 4860
rect 5940 4860 5958 4878
rect 5940 4878 5958 4896
rect 5940 4896 5958 4914
rect 5940 4914 5958 4932
rect 5940 4932 5958 4950
rect 5940 4950 5958 4968
rect 5940 4968 5958 4986
rect 5940 4986 5958 5004
rect 5940 5004 5958 5022
rect 5940 5022 5958 5040
rect 5940 5040 5958 5058
rect 5940 5058 5958 5076
rect 5940 5076 5958 5094
rect 5940 5094 5958 5112
rect 5940 5112 5958 5130
rect 5940 5130 5958 5148
rect 5940 5148 5958 5166
rect 5940 5166 5958 5184
rect 5940 5184 5958 5202
rect 5940 5202 5958 5220
rect 5940 5220 5958 5238
rect 5940 5238 5958 5256
rect 5940 5256 5958 5274
rect 5940 5274 5958 5292
rect 5940 5292 5958 5310
rect 5940 5310 5958 5328
rect 5940 5580 5958 5598
rect 5940 5598 5958 5616
rect 5940 5616 5958 5634
rect 5940 5634 5958 5652
rect 5940 5652 5958 5670
rect 5940 5670 5958 5688
rect 5940 5688 5958 5706
rect 5940 5706 5958 5724
rect 5940 5724 5958 5742
rect 5940 5742 5958 5760
rect 5940 5760 5958 5778
rect 5940 5778 5958 5796
rect 5940 5796 5958 5814
rect 5940 5814 5958 5832
rect 5940 5832 5958 5850
rect 5940 5850 5958 5868
rect 5940 5868 5958 5886
rect 5940 5886 5958 5904
rect 5940 5904 5958 5922
rect 5940 5922 5958 5940
rect 5940 5940 5958 5958
rect 5940 5958 5958 5976
rect 5940 5976 5958 5994
rect 5940 5994 5958 6012
rect 5940 6012 5958 6030
rect 5940 6030 5958 6048
rect 5940 6048 5958 6066
rect 5940 6066 5958 6084
rect 5940 6084 5958 6102
rect 5940 6102 5958 6120
rect 5940 6120 5958 6138
rect 5940 6138 5958 6156
rect 5940 6156 5958 6174
rect 5940 6174 5958 6192
rect 5940 6192 5958 6210
rect 5940 6210 5958 6228
rect 5940 6228 5958 6246
rect 5940 6246 5958 6264
rect 5940 6264 5958 6282
rect 5940 6282 5958 6300
rect 5940 6300 5958 6318
rect 5940 6318 5958 6336
rect 5940 6336 5958 6354
rect 5940 6354 5958 6372
rect 5940 6372 5958 6390
rect 5940 6390 5958 6408
rect 5940 6408 5958 6426
rect 5940 6426 5958 6444
rect 5940 6444 5958 6462
rect 5940 6462 5958 6480
rect 5940 6480 5958 6498
rect 5940 6498 5958 6516
rect 5940 6516 5958 6534
rect 5940 6534 5958 6552
rect 5940 6552 5958 6570
rect 5940 6570 5958 6588
rect 5940 6588 5958 6606
rect 5940 6606 5958 6624
rect 5940 6624 5958 6642
rect 5940 6642 5958 6660
rect 5940 6660 5958 6678
rect 5940 6678 5958 6696
rect 5940 6696 5958 6714
rect 5940 6714 5958 6732
rect 5940 6732 5958 6750
rect 5940 6750 5958 6768
rect 5940 6768 5958 6786
rect 5940 6786 5958 6804
rect 5940 6804 5958 6822
rect 5940 6822 5958 6840
rect 5940 6840 5958 6858
rect 5940 6858 5958 6876
rect 5940 6876 5958 6894
rect 5940 6894 5958 6912
rect 5940 6912 5958 6930
rect 5940 6930 5958 6948
rect 5940 6948 5958 6966
rect 5940 6966 5958 6984
rect 5940 6984 5958 7002
rect 5940 7002 5958 7020
rect 5940 7020 5958 7038
rect 5940 7038 5958 7056
rect 5940 7056 5958 7074
rect 5940 7074 5958 7092
rect 5940 7092 5958 7110
rect 5940 7110 5958 7128
rect 5940 7128 5958 7146
rect 5940 7146 5958 7164
rect 5940 7164 5958 7182
rect 5940 7182 5958 7200
rect 5940 7200 5958 7218
rect 5940 7218 5958 7236
rect 5940 7236 5958 7254
rect 5940 7254 5958 7272
rect 5940 7272 5958 7290
rect 5940 7290 5958 7308
rect 5940 7308 5958 7326
rect 5940 7326 5958 7344
rect 5940 7344 5958 7362
rect 5940 7362 5958 7380
rect 5940 7380 5958 7398
rect 5940 7398 5958 7416
rect 5940 7416 5958 7434
rect 5940 7434 5958 7452
rect 5940 7452 5958 7470
rect 5940 7470 5958 7488
rect 5940 7488 5958 7506
rect 5940 7506 5958 7524
rect 5940 7524 5958 7542
rect 5940 7542 5958 7560
rect 5940 7560 5958 7578
rect 5940 7578 5958 7596
rect 5940 7596 5958 7614
rect 5940 7614 5958 7632
rect 5940 7632 5958 7650
rect 5940 7650 5958 7668
rect 5940 7668 5958 7686
rect 5940 7686 5958 7704
rect 5940 7704 5958 7722
rect 5940 7722 5958 7740
rect 5940 7740 5958 7758
rect 5940 7758 5958 7776
rect 5940 7776 5958 7794
rect 5940 7794 5958 7812
rect 5940 7812 5958 7830
rect 5940 7830 5958 7848
rect 5940 7848 5958 7866
rect 5940 7866 5958 7884
rect 5940 7884 5958 7902
rect 5940 7902 5958 7920
rect 5940 7920 5958 7938
rect 5940 7938 5958 7956
rect 5940 7956 5958 7974
rect 5940 7974 5958 7992
rect 5940 7992 5958 8010
rect 5940 8010 5958 8028
rect 5940 8028 5958 8046
rect 5940 8046 5958 8064
rect 5940 8064 5958 8082
rect 5940 8082 5958 8100
rect 5940 8100 5958 8118
rect 5940 8118 5958 8136
rect 5940 8136 5958 8154
rect 5940 8154 5958 8172
rect 5940 8172 5958 8190
rect 5940 8190 5958 8208
rect 5940 8208 5958 8226
rect 5940 8226 5958 8244
rect 5940 8244 5958 8262
rect 5940 8262 5958 8280
rect 5940 8280 5958 8298
rect 5940 8298 5958 8316
rect 5940 8316 5958 8334
rect 5940 8334 5958 8352
rect 5940 8352 5958 8370
rect 5940 8370 5958 8388
rect 5940 8388 5958 8406
rect 5940 8406 5958 8424
rect 5940 8424 5958 8442
rect 5940 8442 5958 8460
rect 5940 8460 5958 8478
rect 5940 8478 5958 8496
rect 5940 8496 5958 8514
rect 5940 8514 5958 8532
rect 5940 8532 5958 8550
rect 5940 8550 5958 8568
rect 5940 8568 5958 8586
rect 5940 8586 5958 8604
rect 5940 8604 5958 8622
rect 5940 8622 5958 8640
rect 5940 8640 5958 8658
rect 5940 8658 5958 8676
rect 5940 8676 5958 8694
rect 5940 8694 5958 8712
rect 5940 8712 5958 8730
rect 5940 8730 5958 8748
rect 5940 8748 5958 8766
rect 5940 8766 5958 8784
rect 5940 8784 5958 8802
rect 5940 8802 5958 8820
rect 5940 8820 5958 8838
rect 5940 8838 5958 8856
rect 5940 8856 5958 8874
rect 5940 8874 5958 8892
rect 5940 8892 5958 8910
rect 5940 8910 5958 8928
rect 5940 8928 5958 8946
rect 5940 8946 5958 8964
rect 5940 8964 5958 8982
rect 5940 8982 5958 9000
rect 5940 9000 5958 9018
rect 5940 9018 5958 9036
rect 5940 9036 5958 9054
rect 5940 9054 5958 9072
rect 5940 9072 5958 9090
rect 5940 9090 5958 9108
rect 5940 9108 5958 9126
rect 5940 9126 5958 9144
rect 5958 882 5976 900
rect 5958 900 5976 918
rect 5958 918 5976 936
rect 5958 936 5976 954
rect 5958 954 5976 972
rect 5958 972 5976 990
rect 5958 990 5976 1008
rect 5958 1008 5976 1026
rect 5958 1026 5976 1044
rect 5958 1044 5976 1062
rect 5958 1062 5976 1080
rect 5958 1080 5976 1098
rect 5958 1242 5976 1260
rect 5958 1260 5976 1278
rect 5958 1278 5976 1296
rect 5958 1296 5976 1314
rect 5958 1314 5976 1332
rect 5958 1332 5976 1350
rect 5958 1350 5976 1368
rect 5958 1368 5976 1386
rect 5958 1386 5976 1404
rect 5958 1404 5976 1422
rect 5958 1422 5976 1440
rect 5958 1440 5976 1458
rect 5958 1458 5976 1476
rect 5958 1476 5976 1494
rect 5958 1494 5976 1512
rect 5958 1512 5976 1530
rect 5958 1530 5976 1548
rect 5958 1548 5976 1566
rect 5958 1566 5976 1584
rect 5958 1584 5976 1602
rect 5958 1602 5976 1620
rect 5958 1620 5976 1638
rect 5958 1638 5976 1656
rect 5958 1656 5976 1674
rect 5958 1674 5976 1692
rect 5958 1692 5976 1710
rect 5958 1710 5976 1728
rect 5958 1728 5976 1746
rect 5958 1746 5976 1764
rect 5958 1764 5976 1782
rect 5958 1782 5976 1800
rect 5958 1800 5976 1818
rect 5958 1818 5976 1836
rect 5958 1836 5976 1854
rect 5958 1854 5976 1872
rect 5958 1872 5976 1890
rect 5958 1890 5976 1908
rect 5958 1908 5976 1926
rect 5958 1926 5976 1944
rect 5958 1944 5976 1962
rect 5958 1962 5976 1980
rect 5958 1980 5976 1998
rect 5958 1998 5976 2016
rect 5958 2016 5976 2034
rect 5958 2034 5976 2052
rect 5958 2052 5976 2070
rect 5958 2070 5976 2088
rect 5958 2088 5976 2106
rect 5958 2106 5976 2124
rect 5958 2124 5976 2142
rect 5958 2142 5976 2160
rect 5958 2160 5976 2178
rect 5958 2178 5976 2196
rect 5958 2196 5976 2214
rect 5958 2214 5976 2232
rect 5958 2232 5976 2250
rect 5958 2250 5976 2268
rect 5958 2268 5976 2286
rect 5958 2286 5976 2304
rect 5958 2304 5976 2322
rect 5958 2322 5976 2340
rect 5958 2340 5976 2358
rect 5958 2358 5976 2376
rect 5958 2376 5976 2394
rect 5958 2394 5976 2412
rect 5958 2412 5976 2430
rect 5958 2430 5976 2448
rect 5958 2448 5976 2466
rect 5958 2466 5976 2484
rect 5958 2484 5976 2502
rect 5958 2502 5976 2520
rect 5958 2520 5976 2538
rect 5958 2538 5976 2556
rect 5958 2556 5976 2574
rect 5958 2574 5976 2592
rect 5958 2592 5976 2610
rect 5958 2610 5976 2628
rect 5958 2628 5976 2646
rect 5958 2646 5976 2664
rect 5958 2664 5976 2682
rect 5958 2682 5976 2700
rect 5958 2700 5976 2718
rect 5958 2718 5976 2736
rect 5958 2970 5976 2988
rect 5958 2988 5976 3006
rect 5958 3006 5976 3024
rect 5958 3024 5976 3042
rect 5958 3042 5976 3060
rect 5958 3060 5976 3078
rect 5958 3078 5976 3096
rect 5958 3096 5976 3114
rect 5958 3114 5976 3132
rect 5958 3132 5976 3150
rect 5958 3150 5976 3168
rect 5958 3168 5976 3186
rect 5958 3186 5976 3204
rect 5958 3204 5976 3222
rect 5958 3222 5976 3240
rect 5958 3240 5976 3258
rect 5958 3258 5976 3276
rect 5958 3276 5976 3294
rect 5958 3294 5976 3312
rect 5958 3312 5976 3330
rect 5958 3330 5976 3348
rect 5958 3348 5976 3366
rect 5958 3366 5976 3384
rect 5958 3384 5976 3402
rect 5958 3402 5976 3420
rect 5958 3420 5976 3438
rect 5958 3438 5976 3456
rect 5958 3456 5976 3474
rect 5958 3474 5976 3492
rect 5958 3492 5976 3510
rect 5958 3510 5976 3528
rect 5958 3528 5976 3546
rect 5958 3546 5976 3564
rect 5958 3564 5976 3582
rect 5958 3582 5976 3600
rect 5958 3600 5976 3618
rect 5958 3618 5976 3636
rect 5958 3636 5976 3654
rect 5958 3654 5976 3672
rect 5958 3672 5976 3690
rect 5958 3690 5976 3708
rect 5958 3708 5976 3726
rect 5958 3726 5976 3744
rect 5958 3744 5976 3762
rect 5958 3762 5976 3780
rect 5958 3780 5976 3798
rect 5958 3798 5976 3816
rect 5958 3816 5976 3834
rect 5958 3834 5976 3852
rect 5958 3852 5976 3870
rect 5958 3870 5976 3888
rect 5958 3888 5976 3906
rect 5958 3906 5976 3924
rect 5958 3924 5976 3942
rect 5958 3942 5976 3960
rect 5958 3960 5976 3978
rect 5958 3978 5976 3996
rect 5958 3996 5976 4014
rect 5958 4014 5976 4032
rect 5958 4032 5976 4050
rect 5958 4050 5976 4068
rect 5958 4068 5976 4086
rect 5958 4086 5976 4104
rect 5958 4104 5976 4122
rect 5958 4122 5976 4140
rect 5958 4140 5976 4158
rect 5958 4158 5976 4176
rect 5958 4176 5976 4194
rect 5958 4194 5976 4212
rect 5958 4212 5976 4230
rect 5958 4230 5976 4248
rect 5958 4248 5976 4266
rect 5958 4266 5976 4284
rect 5958 4284 5976 4302
rect 5958 4302 5976 4320
rect 5958 4320 5976 4338
rect 5958 4338 5976 4356
rect 5958 4356 5976 4374
rect 5958 4374 5976 4392
rect 5958 4392 5976 4410
rect 5958 4410 5976 4428
rect 5958 4428 5976 4446
rect 5958 4446 5976 4464
rect 5958 4464 5976 4482
rect 5958 4482 5976 4500
rect 5958 4500 5976 4518
rect 5958 4518 5976 4536
rect 5958 4536 5976 4554
rect 5958 4554 5976 4572
rect 5958 4572 5976 4590
rect 5958 4590 5976 4608
rect 5958 4608 5976 4626
rect 5958 4626 5976 4644
rect 5958 4644 5976 4662
rect 5958 4662 5976 4680
rect 5958 4680 5976 4698
rect 5958 4698 5976 4716
rect 5958 4716 5976 4734
rect 5958 4734 5976 4752
rect 5958 4752 5976 4770
rect 5958 4770 5976 4788
rect 5958 4788 5976 4806
rect 5958 4806 5976 4824
rect 5958 4824 5976 4842
rect 5958 4842 5976 4860
rect 5958 4860 5976 4878
rect 5958 4878 5976 4896
rect 5958 4896 5976 4914
rect 5958 4914 5976 4932
rect 5958 4932 5976 4950
rect 5958 4950 5976 4968
rect 5958 4968 5976 4986
rect 5958 4986 5976 5004
rect 5958 5004 5976 5022
rect 5958 5022 5976 5040
rect 5958 5040 5976 5058
rect 5958 5058 5976 5076
rect 5958 5076 5976 5094
rect 5958 5094 5976 5112
rect 5958 5112 5976 5130
rect 5958 5130 5976 5148
rect 5958 5148 5976 5166
rect 5958 5166 5976 5184
rect 5958 5184 5976 5202
rect 5958 5202 5976 5220
rect 5958 5220 5976 5238
rect 5958 5238 5976 5256
rect 5958 5256 5976 5274
rect 5958 5274 5976 5292
rect 5958 5292 5976 5310
rect 5958 5310 5976 5328
rect 5958 5328 5976 5346
rect 5958 5598 5976 5616
rect 5958 5616 5976 5634
rect 5958 5634 5976 5652
rect 5958 5652 5976 5670
rect 5958 5670 5976 5688
rect 5958 5688 5976 5706
rect 5958 5706 5976 5724
rect 5958 5724 5976 5742
rect 5958 5742 5976 5760
rect 5958 5760 5976 5778
rect 5958 5778 5976 5796
rect 5958 5796 5976 5814
rect 5958 5814 5976 5832
rect 5958 5832 5976 5850
rect 5958 5850 5976 5868
rect 5958 5868 5976 5886
rect 5958 5886 5976 5904
rect 5958 5904 5976 5922
rect 5958 5922 5976 5940
rect 5958 5940 5976 5958
rect 5958 5958 5976 5976
rect 5958 5976 5976 5994
rect 5958 5994 5976 6012
rect 5958 6012 5976 6030
rect 5958 6030 5976 6048
rect 5958 6048 5976 6066
rect 5958 6066 5976 6084
rect 5958 6084 5976 6102
rect 5958 6102 5976 6120
rect 5958 6120 5976 6138
rect 5958 6138 5976 6156
rect 5958 6156 5976 6174
rect 5958 6174 5976 6192
rect 5958 6192 5976 6210
rect 5958 6210 5976 6228
rect 5958 6228 5976 6246
rect 5958 6246 5976 6264
rect 5958 6264 5976 6282
rect 5958 6282 5976 6300
rect 5958 6300 5976 6318
rect 5958 6318 5976 6336
rect 5958 6336 5976 6354
rect 5958 6354 5976 6372
rect 5958 6372 5976 6390
rect 5958 6390 5976 6408
rect 5958 6408 5976 6426
rect 5958 6426 5976 6444
rect 5958 6444 5976 6462
rect 5958 6462 5976 6480
rect 5958 6480 5976 6498
rect 5958 6498 5976 6516
rect 5958 6516 5976 6534
rect 5958 6534 5976 6552
rect 5958 6552 5976 6570
rect 5958 6570 5976 6588
rect 5958 6588 5976 6606
rect 5958 6606 5976 6624
rect 5958 6624 5976 6642
rect 5958 6642 5976 6660
rect 5958 6660 5976 6678
rect 5958 6678 5976 6696
rect 5958 6696 5976 6714
rect 5958 6714 5976 6732
rect 5958 6732 5976 6750
rect 5958 6750 5976 6768
rect 5958 6768 5976 6786
rect 5958 6786 5976 6804
rect 5958 6804 5976 6822
rect 5958 6822 5976 6840
rect 5958 6840 5976 6858
rect 5958 6858 5976 6876
rect 5958 6876 5976 6894
rect 5958 6894 5976 6912
rect 5958 6912 5976 6930
rect 5958 6930 5976 6948
rect 5958 6948 5976 6966
rect 5958 6966 5976 6984
rect 5958 6984 5976 7002
rect 5958 7002 5976 7020
rect 5958 7020 5976 7038
rect 5958 7038 5976 7056
rect 5958 7056 5976 7074
rect 5958 7074 5976 7092
rect 5958 7092 5976 7110
rect 5958 7110 5976 7128
rect 5958 7128 5976 7146
rect 5958 7146 5976 7164
rect 5958 7164 5976 7182
rect 5958 7182 5976 7200
rect 5958 7200 5976 7218
rect 5958 7218 5976 7236
rect 5958 7236 5976 7254
rect 5958 7254 5976 7272
rect 5958 7272 5976 7290
rect 5958 7290 5976 7308
rect 5958 7308 5976 7326
rect 5958 7326 5976 7344
rect 5958 7344 5976 7362
rect 5958 7362 5976 7380
rect 5958 7380 5976 7398
rect 5958 7398 5976 7416
rect 5958 7416 5976 7434
rect 5958 7434 5976 7452
rect 5958 7452 5976 7470
rect 5958 7470 5976 7488
rect 5958 7488 5976 7506
rect 5958 7506 5976 7524
rect 5958 7524 5976 7542
rect 5958 7542 5976 7560
rect 5958 7560 5976 7578
rect 5958 7578 5976 7596
rect 5958 7596 5976 7614
rect 5958 7614 5976 7632
rect 5958 7632 5976 7650
rect 5958 7650 5976 7668
rect 5958 7668 5976 7686
rect 5958 7686 5976 7704
rect 5958 7704 5976 7722
rect 5958 7722 5976 7740
rect 5958 7740 5976 7758
rect 5958 7758 5976 7776
rect 5958 7776 5976 7794
rect 5958 7794 5976 7812
rect 5958 7812 5976 7830
rect 5958 7830 5976 7848
rect 5958 7848 5976 7866
rect 5958 7866 5976 7884
rect 5958 7884 5976 7902
rect 5958 7902 5976 7920
rect 5958 7920 5976 7938
rect 5958 7938 5976 7956
rect 5958 7956 5976 7974
rect 5958 7974 5976 7992
rect 5958 7992 5976 8010
rect 5958 8010 5976 8028
rect 5958 8028 5976 8046
rect 5958 8046 5976 8064
rect 5958 8064 5976 8082
rect 5958 8082 5976 8100
rect 5958 8100 5976 8118
rect 5958 8118 5976 8136
rect 5958 8136 5976 8154
rect 5958 8154 5976 8172
rect 5958 8172 5976 8190
rect 5958 8190 5976 8208
rect 5958 8208 5976 8226
rect 5958 8226 5976 8244
rect 5958 8244 5976 8262
rect 5958 8262 5976 8280
rect 5958 8280 5976 8298
rect 5958 8298 5976 8316
rect 5958 8316 5976 8334
rect 5958 8334 5976 8352
rect 5958 8352 5976 8370
rect 5958 8370 5976 8388
rect 5958 8388 5976 8406
rect 5958 8406 5976 8424
rect 5958 8424 5976 8442
rect 5958 8442 5976 8460
rect 5958 8460 5976 8478
rect 5958 8478 5976 8496
rect 5958 8496 5976 8514
rect 5958 8514 5976 8532
rect 5958 8532 5976 8550
rect 5958 8550 5976 8568
rect 5958 8568 5976 8586
rect 5958 8586 5976 8604
rect 5958 8604 5976 8622
rect 5958 8622 5976 8640
rect 5958 8640 5976 8658
rect 5958 8658 5976 8676
rect 5958 8676 5976 8694
rect 5958 8694 5976 8712
rect 5958 8712 5976 8730
rect 5958 8730 5976 8748
rect 5958 8748 5976 8766
rect 5958 8766 5976 8784
rect 5958 8784 5976 8802
rect 5958 8802 5976 8820
rect 5958 8820 5976 8838
rect 5958 8838 5976 8856
rect 5958 8856 5976 8874
rect 5958 8874 5976 8892
rect 5958 8892 5976 8910
rect 5958 8910 5976 8928
rect 5958 8928 5976 8946
rect 5958 8946 5976 8964
rect 5958 8964 5976 8982
rect 5958 8982 5976 9000
rect 5958 9000 5976 9018
rect 5958 9018 5976 9036
rect 5958 9036 5976 9054
rect 5958 9054 5976 9072
rect 5958 9072 5976 9090
rect 5958 9090 5976 9108
rect 5958 9108 5976 9126
rect 5958 9126 5976 9144
rect 5958 9144 5976 9162
rect 5958 9162 5976 9180
rect 5976 882 5994 900
rect 5976 900 5994 918
rect 5976 918 5994 936
rect 5976 936 5994 954
rect 5976 954 5994 972
rect 5976 972 5994 990
rect 5976 990 5994 1008
rect 5976 1008 5994 1026
rect 5976 1026 5994 1044
rect 5976 1044 5994 1062
rect 5976 1062 5994 1080
rect 5976 1080 5994 1098
rect 5976 1242 5994 1260
rect 5976 1260 5994 1278
rect 5976 1278 5994 1296
rect 5976 1296 5994 1314
rect 5976 1314 5994 1332
rect 5976 1332 5994 1350
rect 5976 1350 5994 1368
rect 5976 1368 5994 1386
rect 5976 1386 5994 1404
rect 5976 1404 5994 1422
rect 5976 1422 5994 1440
rect 5976 1440 5994 1458
rect 5976 1458 5994 1476
rect 5976 1476 5994 1494
rect 5976 1494 5994 1512
rect 5976 1512 5994 1530
rect 5976 1530 5994 1548
rect 5976 1548 5994 1566
rect 5976 1566 5994 1584
rect 5976 1584 5994 1602
rect 5976 1602 5994 1620
rect 5976 1620 5994 1638
rect 5976 1638 5994 1656
rect 5976 1656 5994 1674
rect 5976 1674 5994 1692
rect 5976 1692 5994 1710
rect 5976 1710 5994 1728
rect 5976 1728 5994 1746
rect 5976 1746 5994 1764
rect 5976 1764 5994 1782
rect 5976 1782 5994 1800
rect 5976 1800 5994 1818
rect 5976 1818 5994 1836
rect 5976 1836 5994 1854
rect 5976 1854 5994 1872
rect 5976 1872 5994 1890
rect 5976 1890 5994 1908
rect 5976 1908 5994 1926
rect 5976 1926 5994 1944
rect 5976 1944 5994 1962
rect 5976 1962 5994 1980
rect 5976 1980 5994 1998
rect 5976 1998 5994 2016
rect 5976 2016 5994 2034
rect 5976 2034 5994 2052
rect 5976 2052 5994 2070
rect 5976 2070 5994 2088
rect 5976 2088 5994 2106
rect 5976 2106 5994 2124
rect 5976 2124 5994 2142
rect 5976 2142 5994 2160
rect 5976 2160 5994 2178
rect 5976 2178 5994 2196
rect 5976 2196 5994 2214
rect 5976 2214 5994 2232
rect 5976 2232 5994 2250
rect 5976 2250 5994 2268
rect 5976 2268 5994 2286
rect 5976 2286 5994 2304
rect 5976 2304 5994 2322
rect 5976 2322 5994 2340
rect 5976 2340 5994 2358
rect 5976 2358 5994 2376
rect 5976 2376 5994 2394
rect 5976 2394 5994 2412
rect 5976 2412 5994 2430
rect 5976 2430 5994 2448
rect 5976 2448 5994 2466
rect 5976 2466 5994 2484
rect 5976 2484 5994 2502
rect 5976 2502 5994 2520
rect 5976 2520 5994 2538
rect 5976 2538 5994 2556
rect 5976 2556 5994 2574
rect 5976 2574 5994 2592
rect 5976 2592 5994 2610
rect 5976 2610 5994 2628
rect 5976 2628 5994 2646
rect 5976 2646 5994 2664
rect 5976 2664 5994 2682
rect 5976 2682 5994 2700
rect 5976 2700 5994 2718
rect 5976 2718 5994 2736
rect 5976 2970 5994 2988
rect 5976 2988 5994 3006
rect 5976 3006 5994 3024
rect 5976 3024 5994 3042
rect 5976 3042 5994 3060
rect 5976 3060 5994 3078
rect 5976 3078 5994 3096
rect 5976 3096 5994 3114
rect 5976 3114 5994 3132
rect 5976 3132 5994 3150
rect 5976 3150 5994 3168
rect 5976 3168 5994 3186
rect 5976 3186 5994 3204
rect 5976 3204 5994 3222
rect 5976 3222 5994 3240
rect 5976 3240 5994 3258
rect 5976 3258 5994 3276
rect 5976 3276 5994 3294
rect 5976 3294 5994 3312
rect 5976 3312 5994 3330
rect 5976 3330 5994 3348
rect 5976 3348 5994 3366
rect 5976 3366 5994 3384
rect 5976 3384 5994 3402
rect 5976 3402 5994 3420
rect 5976 3420 5994 3438
rect 5976 3438 5994 3456
rect 5976 3456 5994 3474
rect 5976 3474 5994 3492
rect 5976 3492 5994 3510
rect 5976 3510 5994 3528
rect 5976 3528 5994 3546
rect 5976 3546 5994 3564
rect 5976 3564 5994 3582
rect 5976 3582 5994 3600
rect 5976 3600 5994 3618
rect 5976 3618 5994 3636
rect 5976 3636 5994 3654
rect 5976 3654 5994 3672
rect 5976 3672 5994 3690
rect 5976 3690 5994 3708
rect 5976 3708 5994 3726
rect 5976 3726 5994 3744
rect 5976 3744 5994 3762
rect 5976 3762 5994 3780
rect 5976 3780 5994 3798
rect 5976 3798 5994 3816
rect 5976 3816 5994 3834
rect 5976 3834 5994 3852
rect 5976 3852 5994 3870
rect 5976 3870 5994 3888
rect 5976 3888 5994 3906
rect 5976 3906 5994 3924
rect 5976 3924 5994 3942
rect 5976 3942 5994 3960
rect 5976 3960 5994 3978
rect 5976 3978 5994 3996
rect 5976 3996 5994 4014
rect 5976 4014 5994 4032
rect 5976 4032 5994 4050
rect 5976 4050 5994 4068
rect 5976 4068 5994 4086
rect 5976 4086 5994 4104
rect 5976 4104 5994 4122
rect 5976 4122 5994 4140
rect 5976 4140 5994 4158
rect 5976 4158 5994 4176
rect 5976 4176 5994 4194
rect 5976 4194 5994 4212
rect 5976 4212 5994 4230
rect 5976 4230 5994 4248
rect 5976 4248 5994 4266
rect 5976 4266 5994 4284
rect 5976 4284 5994 4302
rect 5976 4302 5994 4320
rect 5976 4320 5994 4338
rect 5976 4338 5994 4356
rect 5976 4356 5994 4374
rect 5976 4374 5994 4392
rect 5976 4392 5994 4410
rect 5976 4410 5994 4428
rect 5976 4428 5994 4446
rect 5976 4446 5994 4464
rect 5976 4464 5994 4482
rect 5976 4482 5994 4500
rect 5976 4500 5994 4518
rect 5976 4518 5994 4536
rect 5976 4536 5994 4554
rect 5976 4554 5994 4572
rect 5976 4572 5994 4590
rect 5976 4590 5994 4608
rect 5976 4608 5994 4626
rect 5976 4626 5994 4644
rect 5976 4644 5994 4662
rect 5976 4662 5994 4680
rect 5976 4680 5994 4698
rect 5976 4698 5994 4716
rect 5976 4716 5994 4734
rect 5976 4734 5994 4752
rect 5976 4752 5994 4770
rect 5976 4770 5994 4788
rect 5976 4788 5994 4806
rect 5976 4806 5994 4824
rect 5976 4824 5994 4842
rect 5976 4842 5994 4860
rect 5976 4860 5994 4878
rect 5976 4878 5994 4896
rect 5976 4896 5994 4914
rect 5976 4914 5994 4932
rect 5976 4932 5994 4950
rect 5976 4950 5994 4968
rect 5976 4968 5994 4986
rect 5976 4986 5994 5004
rect 5976 5004 5994 5022
rect 5976 5022 5994 5040
rect 5976 5040 5994 5058
rect 5976 5058 5994 5076
rect 5976 5076 5994 5094
rect 5976 5094 5994 5112
rect 5976 5112 5994 5130
rect 5976 5130 5994 5148
rect 5976 5148 5994 5166
rect 5976 5166 5994 5184
rect 5976 5184 5994 5202
rect 5976 5202 5994 5220
rect 5976 5220 5994 5238
rect 5976 5238 5994 5256
rect 5976 5256 5994 5274
rect 5976 5274 5994 5292
rect 5976 5292 5994 5310
rect 5976 5310 5994 5328
rect 5976 5328 5994 5346
rect 5976 5346 5994 5364
rect 5976 5616 5994 5634
rect 5976 5634 5994 5652
rect 5976 5652 5994 5670
rect 5976 5670 5994 5688
rect 5976 5688 5994 5706
rect 5976 5706 5994 5724
rect 5976 5724 5994 5742
rect 5976 5742 5994 5760
rect 5976 5760 5994 5778
rect 5976 5778 5994 5796
rect 5976 5796 5994 5814
rect 5976 5814 5994 5832
rect 5976 5832 5994 5850
rect 5976 5850 5994 5868
rect 5976 5868 5994 5886
rect 5976 5886 5994 5904
rect 5976 5904 5994 5922
rect 5976 5922 5994 5940
rect 5976 5940 5994 5958
rect 5976 5958 5994 5976
rect 5976 5976 5994 5994
rect 5976 5994 5994 6012
rect 5976 6012 5994 6030
rect 5976 6030 5994 6048
rect 5976 6048 5994 6066
rect 5976 6066 5994 6084
rect 5976 6084 5994 6102
rect 5976 6102 5994 6120
rect 5976 6120 5994 6138
rect 5976 6138 5994 6156
rect 5976 6156 5994 6174
rect 5976 6174 5994 6192
rect 5976 6192 5994 6210
rect 5976 6210 5994 6228
rect 5976 6228 5994 6246
rect 5976 6246 5994 6264
rect 5976 6264 5994 6282
rect 5976 6282 5994 6300
rect 5976 6300 5994 6318
rect 5976 6318 5994 6336
rect 5976 6336 5994 6354
rect 5976 6354 5994 6372
rect 5976 6372 5994 6390
rect 5976 6390 5994 6408
rect 5976 6408 5994 6426
rect 5976 6426 5994 6444
rect 5976 6444 5994 6462
rect 5976 6462 5994 6480
rect 5976 6480 5994 6498
rect 5976 6498 5994 6516
rect 5976 6516 5994 6534
rect 5976 6534 5994 6552
rect 5976 6552 5994 6570
rect 5976 6570 5994 6588
rect 5976 6588 5994 6606
rect 5976 6606 5994 6624
rect 5976 6624 5994 6642
rect 5976 6642 5994 6660
rect 5976 6660 5994 6678
rect 5976 6678 5994 6696
rect 5976 6696 5994 6714
rect 5976 6714 5994 6732
rect 5976 6732 5994 6750
rect 5976 6750 5994 6768
rect 5976 6768 5994 6786
rect 5976 6786 5994 6804
rect 5976 6804 5994 6822
rect 5976 6822 5994 6840
rect 5976 6840 5994 6858
rect 5976 6858 5994 6876
rect 5976 6876 5994 6894
rect 5976 6894 5994 6912
rect 5976 6912 5994 6930
rect 5976 6930 5994 6948
rect 5976 6948 5994 6966
rect 5976 6966 5994 6984
rect 5976 6984 5994 7002
rect 5976 7002 5994 7020
rect 5976 7020 5994 7038
rect 5976 7038 5994 7056
rect 5976 7056 5994 7074
rect 5976 7074 5994 7092
rect 5976 7092 5994 7110
rect 5976 7110 5994 7128
rect 5976 7128 5994 7146
rect 5976 7146 5994 7164
rect 5976 7164 5994 7182
rect 5976 7182 5994 7200
rect 5976 7200 5994 7218
rect 5976 7218 5994 7236
rect 5976 7236 5994 7254
rect 5976 7254 5994 7272
rect 5976 7272 5994 7290
rect 5976 7290 5994 7308
rect 5976 7308 5994 7326
rect 5976 7326 5994 7344
rect 5976 7344 5994 7362
rect 5976 7362 5994 7380
rect 5976 7380 5994 7398
rect 5976 7398 5994 7416
rect 5976 7416 5994 7434
rect 5976 7434 5994 7452
rect 5976 7452 5994 7470
rect 5976 7470 5994 7488
rect 5976 7488 5994 7506
rect 5976 7506 5994 7524
rect 5976 7524 5994 7542
rect 5976 7542 5994 7560
rect 5976 7560 5994 7578
rect 5976 7578 5994 7596
rect 5976 7596 5994 7614
rect 5976 7614 5994 7632
rect 5976 7632 5994 7650
rect 5976 7650 5994 7668
rect 5976 7668 5994 7686
rect 5976 7686 5994 7704
rect 5976 7704 5994 7722
rect 5976 7722 5994 7740
rect 5976 7740 5994 7758
rect 5976 7758 5994 7776
rect 5976 7776 5994 7794
rect 5976 7794 5994 7812
rect 5976 7812 5994 7830
rect 5976 7830 5994 7848
rect 5976 7848 5994 7866
rect 5976 7866 5994 7884
rect 5976 7884 5994 7902
rect 5976 7902 5994 7920
rect 5976 7920 5994 7938
rect 5976 7938 5994 7956
rect 5976 7956 5994 7974
rect 5976 7974 5994 7992
rect 5976 7992 5994 8010
rect 5976 8010 5994 8028
rect 5976 8028 5994 8046
rect 5976 8046 5994 8064
rect 5976 8064 5994 8082
rect 5976 8082 5994 8100
rect 5976 8100 5994 8118
rect 5976 8118 5994 8136
rect 5976 8136 5994 8154
rect 5976 8154 5994 8172
rect 5976 8172 5994 8190
rect 5976 8190 5994 8208
rect 5976 8208 5994 8226
rect 5976 8226 5994 8244
rect 5976 8244 5994 8262
rect 5976 8262 5994 8280
rect 5976 8280 5994 8298
rect 5976 8298 5994 8316
rect 5976 8316 5994 8334
rect 5976 8334 5994 8352
rect 5976 8352 5994 8370
rect 5976 8370 5994 8388
rect 5976 8388 5994 8406
rect 5976 8406 5994 8424
rect 5976 8424 5994 8442
rect 5976 8442 5994 8460
rect 5976 8460 5994 8478
rect 5976 8478 5994 8496
rect 5976 8496 5994 8514
rect 5976 8514 5994 8532
rect 5976 8532 5994 8550
rect 5976 8550 5994 8568
rect 5976 8568 5994 8586
rect 5976 8586 5994 8604
rect 5976 8604 5994 8622
rect 5976 8622 5994 8640
rect 5976 8640 5994 8658
rect 5976 8658 5994 8676
rect 5976 8676 5994 8694
rect 5976 8694 5994 8712
rect 5976 8712 5994 8730
rect 5976 8730 5994 8748
rect 5976 8748 5994 8766
rect 5976 8766 5994 8784
rect 5976 8784 5994 8802
rect 5976 8802 5994 8820
rect 5976 8820 5994 8838
rect 5976 8838 5994 8856
rect 5976 8856 5994 8874
rect 5976 8874 5994 8892
rect 5976 8892 5994 8910
rect 5976 8910 5994 8928
rect 5976 8928 5994 8946
rect 5976 8946 5994 8964
rect 5976 8964 5994 8982
rect 5976 8982 5994 9000
rect 5976 9000 5994 9018
rect 5976 9018 5994 9036
rect 5976 9036 5994 9054
rect 5976 9054 5994 9072
rect 5976 9072 5994 9090
rect 5976 9090 5994 9108
rect 5976 9108 5994 9126
rect 5976 9126 5994 9144
rect 5976 9144 5994 9162
rect 5976 9162 5994 9180
rect 5976 9180 5994 9198
rect 5994 900 6012 918
rect 5994 918 6012 936
rect 5994 936 6012 954
rect 5994 954 6012 972
rect 5994 972 6012 990
rect 5994 990 6012 1008
rect 5994 1008 6012 1026
rect 5994 1026 6012 1044
rect 5994 1044 6012 1062
rect 5994 1062 6012 1080
rect 5994 1080 6012 1098
rect 5994 1260 6012 1278
rect 5994 1278 6012 1296
rect 5994 1296 6012 1314
rect 5994 1314 6012 1332
rect 5994 1332 6012 1350
rect 5994 1350 6012 1368
rect 5994 1368 6012 1386
rect 5994 1386 6012 1404
rect 5994 1404 6012 1422
rect 5994 1422 6012 1440
rect 5994 1440 6012 1458
rect 5994 1458 6012 1476
rect 5994 1476 6012 1494
rect 5994 1494 6012 1512
rect 5994 1512 6012 1530
rect 5994 1530 6012 1548
rect 5994 1548 6012 1566
rect 5994 1566 6012 1584
rect 5994 1584 6012 1602
rect 5994 1602 6012 1620
rect 5994 1620 6012 1638
rect 5994 1638 6012 1656
rect 5994 1656 6012 1674
rect 5994 1674 6012 1692
rect 5994 1692 6012 1710
rect 5994 1710 6012 1728
rect 5994 1728 6012 1746
rect 5994 1746 6012 1764
rect 5994 1764 6012 1782
rect 5994 1782 6012 1800
rect 5994 1800 6012 1818
rect 5994 1818 6012 1836
rect 5994 1836 6012 1854
rect 5994 1854 6012 1872
rect 5994 1872 6012 1890
rect 5994 1890 6012 1908
rect 5994 1908 6012 1926
rect 5994 1926 6012 1944
rect 5994 1944 6012 1962
rect 5994 1962 6012 1980
rect 5994 1980 6012 1998
rect 5994 1998 6012 2016
rect 5994 2016 6012 2034
rect 5994 2034 6012 2052
rect 5994 2052 6012 2070
rect 5994 2070 6012 2088
rect 5994 2088 6012 2106
rect 5994 2106 6012 2124
rect 5994 2124 6012 2142
rect 5994 2142 6012 2160
rect 5994 2160 6012 2178
rect 5994 2178 6012 2196
rect 5994 2196 6012 2214
rect 5994 2214 6012 2232
rect 5994 2232 6012 2250
rect 5994 2250 6012 2268
rect 5994 2268 6012 2286
rect 5994 2286 6012 2304
rect 5994 2304 6012 2322
rect 5994 2322 6012 2340
rect 5994 2340 6012 2358
rect 5994 2358 6012 2376
rect 5994 2376 6012 2394
rect 5994 2394 6012 2412
rect 5994 2412 6012 2430
rect 5994 2430 6012 2448
rect 5994 2448 6012 2466
rect 5994 2466 6012 2484
rect 5994 2484 6012 2502
rect 5994 2502 6012 2520
rect 5994 2520 6012 2538
rect 5994 2538 6012 2556
rect 5994 2556 6012 2574
rect 5994 2574 6012 2592
rect 5994 2592 6012 2610
rect 5994 2610 6012 2628
rect 5994 2628 6012 2646
rect 5994 2646 6012 2664
rect 5994 2664 6012 2682
rect 5994 2682 6012 2700
rect 5994 2700 6012 2718
rect 5994 2718 6012 2736
rect 5994 2736 6012 2754
rect 5994 2988 6012 3006
rect 5994 3006 6012 3024
rect 5994 3024 6012 3042
rect 5994 3042 6012 3060
rect 5994 3060 6012 3078
rect 5994 3078 6012 3096
rect 5994 3096 6012 3114
rect 5994 3114 6012 3132
rect 5994 3132 6012 3150
rect 5994 3150 6012 3168
rect 5994 3168 6012 3186
rect 5994 3186 6012 3204
rect 5994 3204 6012 3222
rect 5994 3222 6012 3240
rect 5994 3240 6012 3258
rect 5994 3258 6012 3276
rect 5994 3276 6012 3294
rect 5994 3294 6012 3312
rect 5994 3312 6012 3330
rect 5994 3330 6012 3348
rect 5994 3348 6012 3366
rect 5994 3366 6012 3384
rect 5994 3384 6012 3402
rect 5994 3402 6012 3420
rect 5994 3420 6012 3438
rect 5994 3438 6012 3456
rect 5994 3456 6012 3474
rect 5994 3474 6012 3492
rect 5994 3492 6012 3510
rect 5994 3510 6012 3528
rect 5994 3528 6012 3546
rect 5994 3546 6012 3564
rect 5994 3564 6012 3582
rect 5994 3582 6012 3600
rect 5994 3600 6012 3618
rect 5994 3618 6012 3636
rect 5994 3636 6012 3654
rect 5994 3654 6012 3672
rect 5994 3672 6012 3690
rect 5994 3690 6012 3708
rect 5994 3708 6012 3726
rect 5994 3726 6012 3744
rect 5994 3744 6012 3762
rect 5994 3762 6012 3780
rect 5994 3780 6012 3798
rect 5994 3798 6012 3816
rect 5994 3816 6012 3834
rect 5994 3834 6012 3852
rect 5994 3852 6012 3870
rect 5994 3870 6012 3888
rect 5994 3888 6012 3906
rect 5994 3906 6012 3924
rect 5994 3924 6012 3942
rect 5994 3942 6012 3960
rect 5994 3960 6012 3978
rect 5994 3978 6012 3996
rect 5994 3996 6012 4014
rect 5994 4014 6012 4032
rect 5994 4032 6012 4050
rect 5994 4050 6012 4068
rect 5994 4068 6012 4086
rect 5994 4086 6012 4104
rect 5994 4104 6012 4122
rect 5994 4122 6012 4140
rect 5994 4140 6012 4158
rect 5994 4158 6012 4176
rect 5994 4176 6012 4194
rect 5994 4194 6012 4212
rect 5994 4212 6012 4230
rect 5994 4230 6012 4248
rect 5994 4248 6012 4266
rect 5994 4266 6012 4284
rect 5994 4284 6012 4302
rect 5994 4302 6012 4320
rect 5994 4320 6012 4338
rect 5994 4338 6012 4356
rect 5994 4356 6012 4374
rect 5994 4374 6012 4392
rect 5994 4392 6012 4410
rect 5994 4410 6012 4428
rect 5994 4428 6012 4446
rect 5994 4446 6012 4464
rect 5994 4464 6012 4482
rect 5994 4482 6012 4500
rect 5994 4500 6012 4518
rect 5994 4518 6012 4536
rect 5994 4536 6012 4554
rect 5994 4554 6012 4572
rect 5994 4572 6012 4590
rect 5994 4590 6012 4608
rect 5994 4608 6012 4626
rect 5994 4626 6012 4644
rect 5994 4644 6012 4662
rect 5994 4662 6012 4680
rect 5994 4680 6012 4698
rect 5994 4698 6012 4716
rect 5994 4716 6012 4734
rect 5994 4734 6012 4752
rect 5994 4752 6012 4770
rect 5994 4770 6012 4788
rect 5994 4788 6012 4806
rect 5994 4806 6012 4824
rect 5994 4824 6012 4842
rect 5994 4842 6012 4860
rect 5994 4860 6012 4878
rect 5994 4878 6012 4896
rect 5994 4896 6012 4914
rect 5994 4914 6012 4932
rect 5994 4932 6012 4950
rect 5994 4950 6012 4968
rect 5994 4968 6012 4986
rect 5994 4986 6012 5004
rect 5994 5004 6012 5022
rect 5994 5022 6012 5040
rect 5994 5040 6012 5058
rect 5994 5058 6012 5076
rect 5994 5076 6012 5094
rect 5994 5094 6012 5112
rect 5994 5112 6012 5130
rect 5994 5130 6012 5148
rect 5994 5148 6012 5166
rect 5994 5166 6012 5184
rect 5994 5184 6012 5202
rect 5994 5202 6012 5220
rect 5994 5220 6012 5238
rect 5994 5238 6012 5256
rect 5994 5256 6012 5274
rect 5994 5274 6012 5292
rect 5994 5292 6012 5310
rect 5994 5310 6012 5328
rect 5994 5328 6012 5346
rect 5994 5346 6012 5364
rect 5994 5364 6012 5382
rect 5994 5634 6012 5652
rect 5994 5652 6012 5670
rect 5994 5670 6012 5688
rect 5994 5688 6012 5706
rect 5994 5706 6012 5724
rect 5994 5724 6012 5742
rect 5994 5742 6012 5760
rect 5994 5760 6012 5778
rect 5994 5778 6012 5796
rect 5994 5796 6012 5814
rect 5994 5814 6012 5832
rect 5994 5832 6012 5850
rect 5994 5850 6012 5868
rect 5994 5868 6012 5886
rect 5994 5886 6012 5904
rect 5994 5904 6012 5922
rect 5994 5922 6012 5940
rect 5994 5940 6012 5958
rect 5994 5958 6012 5976
rect 5994 5976 6012 5994
rect 5994 5994 6012 6012
rect 5994 6012 6012 6030
rect 5994 6030 6012 6048
rect 5994 6048 6012 6066
rect 5994 6066 6012 6084
rect 5994 6084 6012 6102
rect 5994 6102 6012 6120
rect 5994 6120 6012 6138
rect 5994 6138 6012 6156
rect 5994 6156 6012 6174
rect 5994 6174 6012 6192
rect 5994 6192 6012 6210
rect 5994 6210 6012 6228
rect 5994 6228 6012 6246
rect 5994 6246 6012 6264
rect 5994 6264 6012 6282
rect 5994 6282 6012 6300
rect 5994 6300 6012 6318
rect 5994 6318 6012 6336
rect 5994 6336 6012 6354
rect 5994 6354 6012 6372
rect 5994 6372 6012 6390
rect 5994 6390 6012 6408
rect 5994 6408 6012 6426
rect 5994 6426 6012 6444
rect 5994 6444 6012 6462
rect 5994 6462 6012 6480
rect 5994 6480 6012 6498
rect 5994 6498 6012 6516
rect 5994 6516 6012 6534
rect 5994 6534 6012 6552
rect 5994 6552 6012 6570
rect 5994 6570 6012 6588
rect 5994 6588 6012 6606
rect 5994 6606 6012 6624
rect 5994 6624 6012 6642
rect 5994 6642 6012 6660
rect 5994 6660 6012 6678
rect 5994 6678 6012 6696
rect 5994 6696 6012 6714
rect 5994 6714 6012 6732
rect 5994 6732 6012 6750
rect 5994 6750 6012 6768
rect 5994 6768 6012 6786
rect 5994 6786 6012 6804
rect 5994 6804 6012 6822
rect 5994 6822 6012 6840
rect 5994 6840 6012 6858
rect 5994 6858 6012 6876
rect 5994 6876 6012 6894
rect 5994 6894 6012 6912
rect 5994 6912 6012 6930
rect 5994 6930 6012 6948
rect 5994 6948 6012 6966
rect 5994 6966 6012 6984
rect 5994 6984 6012 7002
rect 5994 7002 6012 7020
rect 5994 7020 6012 7038
rect 5994 7038 6012 7056
rect 5994 7056 6012 7074
rect 5994 7074 6012 7092
rect 5994 7092 6012 7110
rect 5994 7110 6012 7128
rect 5994 7128 6012 7146
rect 5994 7146 6012 7164
rect 5994 7164 6012 7182
rect 5994 7182 6012 7200
rect 5994 7200 6012 7218
rect 5994 7218 6012 7236
rect 5994 7236 6012 7254
rect 5994 7254 6012 7272
rect 5994 7272 6012 7290
rect 5994 7290 6012 7308
rect 5994 7308 6012 7326
rect 5994 7326 6012 7344
rect 5994 7344 6012 7362
rect 5994 7362 6012 7380
rect 5994 7380 6012 7398
rect 5994 7398 6012 7416
rect 5994 7416 6012 7434
rect 5994 7434 6012 7452
rect 5994 7452 6012 7470
rect 5994 7470 6012 7488
rect 5994 7488 6012 7506
rect 5994 7506 6012 7524
rect 5994 7524 6012 7542
rect 5994 7542 6012 7560
rect 5994 7560 6012 7578
rect 5994 7578 6012 7596
rect 5994 7596 6012 7614
rect 5994 7614 6012 7632
rect 5994 7632 6012 7650
rect 5994 7650 6012 7668
rect 5994 7668 6012 7686
rect 5994 7686 6012 7704
rect 5994 7704 6012 7722
rect 5994 7722 6012 7740
rect 5994 7740 6012 7758
rect 5994 7758 6012 7776
rect 5994 7776 6012 7794
rect 5994 7794 6012 7812
rect 5994 7812 6012 7830
rect 5994 7830 6012 7848
rect 5994 7848 6012 7866
rect 5994 7866 6012 7884
rect 5994 7884 6012 7902
rect 5994 7902 6012 7920
rect 5994 7920 6012 7938
rect 5994 7938 6012 7956
rect 5994 7956 6012 7974
rect 5994 7974 6012 7992
rect 5994 7992 6012 8010
rect 5994 8010 6012 8028
rect 5994 8028 6012 8046
rect 5994 8046 6012 8064
rect 5994 8064 6012 8082
rect 5994 8082 6012 8100
rect 5994 8100 6012 8118
rect 5994 8118 6012 8136
rect 5994 8136 6012 8154
rect 5994 8154 6012 8172
rect 5994 8172 6012 8190
rect 5994 8190 6012 8208
rect 5994 8208 6012 8226
rect 5994 8226 6012 8244
rect 5994 8244 6012 8262
rect 5994 8262 6012 8280
rect 5994 8280 6012 8298
rect 5994 8298 6012 8316
rect 5994 8316 6012 8334
rect 5994 8334 6012 8352
rect 5994 8352 6012 8370
rect 5994 8370 6012 8388
rect 5994 8388 6012 8406
rect 5994 8406 6012 8424
rect 5994 8424 6012 8442
rect 5994 8442 6012 8460
rect 5994 8460 6012 8478
rect 5994 8478 6012 8496
rect 5994 8496 6012 8514
rect 5994 8514 6012 8532
rect 5994 8532 6012 8550
rect 5994 8550 6012 8568
rect 5994 8568 6012 8586
rect 5994 8586 6012 8604
rect 5994 8604 6012 8622
rect 5994 8622 6012 8640
rect 5994 8640 6012 8658
rect 5994 8658 6012 8676
rect 5994 8676 6012 8694
rect 5994 8694 6012 8712
rect 5994 8712 6012 8730
rect 5994 8730 6012 8748
rect 5994 8748 6012 8766
rect 5994 8766 6012 8784
rect 5994 8784 6012 8802
rect 5994 8802 6012 8820
rect 5994 8820 6012 8838
rect 5994 8838 6012 8856
rect 5994 8856 6012 8874
rect 5994 8874 6012 8892
rect 5994 8892 6012 8910
rect 5994 8910 6012 8928
rect 5994 8928 6012 8946
rect 5994 8946 6012 8964
rect 5994 8964 6012 8982
rect 5994 8982 6012 9000
rect 5994 9000 6012 9018
rect 5994 9018 6012 9036
rect 5994 9036 6012 9054
rect 5994 9054 6012 9072
rect 5994 9072 6012 9090
rect 5994 9090 6012 9108
rect 5994 9108 6012 9126
rect 5994 9126 6012 9144
rect 5994 9144 6012 9162
rect 5994 9162 6012 9180
rect 5994 9180 6012 9198
rect 5994 9198 6012 9216
rect 6012 918 6030 936
rect 6012 936 6030 954
rect 6012 954 6030 972
rect 6012 972 6030 990
rect 6012 990 6030 1008
rect 6012 1008 6030 1026
rect 6012 1026 6030 1044
rect 6012 1044 6030 1062
rect 6012 1062 6030 1080
rect 6012 1080 6030 1098
rect 6012 1098 6030 1116
rect 6012 1260 6030 1278
rect 6012 1278 6030 1296
rect 6012 1296 6030 1314
rect 6012 1314 6030 1332
rect 6012 1332 6030 1350
rect 6012 1350 6030 1368
rect 6012 1368 6030 1386
rect 6012 1386 6030 1404
rect 6012 1404 6030 1422
rect 6012 1422 6030 1440
rect 6012 1440 6030 1458
rect 6012 1458 6030 1476
rect 6012 1476 6030 1494
rect 6012 1494 6030 1512
rect 6012 1512 6030 1530
rect 6012 1530 6030 1548
rect 6012 1548 6030 1566
rect 6012 1566 6030 1584
rect 6012 1584 6030 1602
rect 6012 1602 6030 1620
rect 6012 1620 6030 1638
rect 6012 1638 6030 1656
rect 6012 1656 6030 1674
rect 6012 1674 6030 1692
rect 6012 1692 6030 1710
rect 6012 1710 6030 1728
rect 6012 1728 6030 1746
rect 6012 1746 6030 1764
rect 6012 1764 6030 1782
rect 6012 1782 6030 1800
rect 6012 1800 6030 1818
rect 6012 1818 6030 1836
rect 6012 1836 6030 1854
rect 6012 1854 6030 1872
rect 6012 1872 6030 1890
rect 6012 1890 6030 1908
rect 6012 1908 6030 1926
rect 6012 1926 6030 1944
rect 6012 1944 6030 1962
rect 6012 1962 6030 1980
rect 6012 1980 6030 1998
rect 6012 1998 6030 2016
rect 6012 2016 6030 2034
rect 6012 2034 6030 2052
rect 6012 2052 6030 2070
rect 6012 2070 6030 2088
rect 6012 2088 6030 2106
rect 6012 2106 6030 2124
rect 6012 2124 6030 2142
rect 6012 2142 6030 2160
rect 6012 2160 6030 2178
rect 6012 2178 6030 2196
rect 6012 2196 6030 2214
rect 6012 2214 6030 2232
rect 6012 2232 6030 2250
rect 6012 2250 6030 2268
rect 6012 2268 6030 2286
rect 6012 2286 6030 2304
rect 6012 2304 6030 2322
rect 6012 2322 6030 2340
rect 6012 2340 6030 2358
rect 6012 2358 6030 2376
rect 6012 2376 6030 2394
rect 6012 2394 6030 2412
rect 6012 2412 6030 2430
rect 6012 2430 6030 2448
rect 6012 2448 6030 2466
rect 6012 2466 6030 2484
rect 6012 2484 6030 2502
rect 6012 2502 6030 2520
rect 6012 2520 6030 2538
rect 6012 2538 6030 2556
rect 6012 2556 6030 2574
rect 6012 2574 6030 2592
rect 6012 2592 6030 2610
rect 6012 2610 6030 2628
rect 6012 2628 6030 2646
rect 6012 2646 6030 2664
rect 6012 2664 6030 2682
rect 6012 2682 6030 2700
rect 6012 2700 6030 2718
rect 6012 2718 6030 2736
rect 6012 2736 6030 2754
rect 6012 2988 6030 3006
rect 6012 3006 6030 3024
rect 6012 3024 6030 3042
rect 6012 3042 6030 3060
rect 6012 3060 6030 3078
rect 6012 3078 6030 3096
rect 6012 3096 6030 3114
rect 6012 3114 6030 3132
rect 6012 3132 6030 3150
rect 6012 3150 6030 3168
rect 6012 3168 6030 3186
rect 6012 3186 6030 3204
rect 6012 3204 6030 3222
rect 6012 3222 6030 3240
rect 6012 3240 6030 3258
rect 6012 3258 6030 3276
rect 6012 3276 6030 3294
rect 6012 3294 6030 3312
rect 6012 3312 6030 3330
rect 6012 3330 6030 3348
rect 6012 3348 6030 3366
rect 6012 3366 6030 3384
rect 6012 3384 6030 3402
rect 6012 3402 6030 3420
rect 6012 3420 6030 3438
rect 6012 3438 6030 3456
rect 6012 3456 6030 3474
rect 6012 3474 6030 3492
rect 6012 3492 6030 3510
rect 6012 3510 6030 3528
rect 6012 3528 6030 3546
rect 6012 3546 6030 3564
rect 6012 3564 6030 3582
rect 6012 3582 6030 3600
rect 6012 3600 6030 3618
rect 6012 3618 6030 3636
rect 6012 3636 6030 3654
rect 6012 3654 6030 3672
rect 6012 3672 6030 3690
rect 6012 3690 6030 3708
rect 6012 3708 6030 3726
rect 6012 3726 6030 3744
rect 6012 3744 6030 3762
rect 6012 3762 6030 3780
rect 6012 3780 6030 3798
rect 6012 3798 6030 3816
rect 6012 3816 6030 3834
rect 6012 3834 6030 3852
rect 6012 3852 6030 3870
rect 6012 3870 6030 3888
rect 6012 3888 6030 3906
rect 6012 3906 6030 3924
rect 6012 3924 6030 3942
rect 6012 3942 6030 3960
rect 6012 3960 6030 3978
rect 6012 3978 6030 3996
rect 6012 3996 6030 4014
rect 6012 4014 6030 4032
rect 6012 4032 6030 4050
rect 6012 4050 6030 4068
rect 6012 4068 6030 4086
rect 6012 4086 6030 4104
rect 6012 4104 6030 4122
rect 6012 4122 6030 4140
rect 6012 4140 6030 4158
rect 6012 4158 6030 4176
rect 6012 4176 6030 4194
rect 6012 4194 6030 4212
rect 6012 4212 6030 4230
rect 6012 4230 6030 4248
rect 6012 4248 6030 4266
rect 6012 4266 6030 4284
rect 6012 4284 6030 4302
rect 6012 4302 6030 4320
rect 6012 4320 6030 4338
rect 6012 4338 6030 4356
rect 6012 4356 6030 4374
rect 6012 4374 6030 4392
rect 6012 4392 6030 4410
rect 6012 4410 6030 4428
rect 6012 4428 6030 4446
rect 6012 4446 6030 4464
rect 6012 4464 6030 4482
rect 6012 4482 6030 4500
rect 6012 4500 6030 4518
rect 6012 4518 6030 4536
rect 6012 4536 6030 4554
rect 6012 4554 6030 4572
rect 6012 4572 6030 4590
rect 6012 4590 6030 4608
rect 6012 4608 6030 4626
rect 6012 4626 6030 4644
rect 6012 4644 6030 4662
rect 6012 4662 6030 4680
rect 6012 4680 6030 4698
rect 6012 4698 6030 4716
rect 6012 4716 6030 4734
rect 6012 4734 6030 4752
rect 6012 4752 6030 4770
rect 6012 4770 6030 4788
rect 6012 4788 6030 4806
rect 6012 4806 6030 4824
rect 6012 4824 6030 4842
rect 6012 4842 6030 4860
rect 6012 4860 6030 4878
rect 6012 4878 6030 4896
rect 6012 4896 6030 4914
rect 6012 4914 6030 4932
rect 6012 4932 6030 4950
rect 6012 4950 6030 4968
rect 6012 4968 6030 4986
rect 6012 4986 6030 5004
rect 6012 5004 6030 5022
rect 6012 5022 6030 5040
rect 6012 5040 6030 5058
rect 6012 5058 6030 5076
rect 6012 5076 6030 5094
rect 6012 5094 6030 5112
rect 6012 5112 6030 5130
rect 6012 5130 6030 5148
rect 6012 5148 6030 5166
rect 6012 5166 6030 5184
rect 6012 5184 6030 5202
rect 6012 5202 6030 5220
rect 6012 5220 6030 5238
rect 6012 5238 6030 5256
rect 6012 5256 6030 5274
rect 6012 5274 6030 5292
rect 6012 5292 6030 5310
rect 6012 5310 6030 5328
rect 6012 5328 6030 5346
rect 6012 5346 6030 5364
rect 6012 5364 6030 5382
rect 6012 5382 6030 5400
rect 6012 5652 6030 5670
rect 6012 5670 6030 5688
rect 6012 5688 6030 5706
rect 6012 5706 6030 5724
rect 6012 5724 6030 5742
rect 6012 5742 6030 5760
rect 6012 5760 6030 5778
rect 6012 5778 6030 5796
rect 6012 5796 6030 5814
rect 6012 5814 6030 5832
rect 6012 5832 6030 5850
rect 6012 5850 6030 5868
rect 6012 5868 6030 5886
rect 6012 5886 6030 5904
rect 6012 5904 6030 5922
rect 6012 5922 6030 5940
rect 6012 5940 6030 5958
rect 6012 5958 6030 5976
rect 6012 5976 6030 5994
rect 6012 5994 6030 6012
rect 6012 6012 6030 6030
rect 6012 6030 6030 6048
rect 6012 6048 6030 6066
rect 6012 6066 6030 6084
rect 6012 6084 6030 6102
rect 6012 6102 6030 6120
rect 6012 6120 6030 6138
rect 6012 6138 6030 6156
rect 6012 6156 6030 6174
rect 6012 6174 6030 6192
rect 6012 6192 6030 6210
rect 6012 6210 6030 6228
rect 6012 6228 6030 6246
rect 6012 6246 6030 6264
rect 6012 6264 6030 6282
rect 6012 6282 6030 6300
rect 6012 6300 6030 6318
rect 6012 6318 6030 6336
rect 6012 6336 6030 6354
rect 6012 6354 6030 6372
rect 6012 6372 6030 6390
rect 6012 6390 6030 6408
rect 6012 6408 6030 6426
rect 6012 6426 6030 6444
rect 6012 6444 6030 6462
rect 6012 6462 6030 6480
rect 6012 6480 6030 6498
rect 6012 6498 6030 6516
rect 6012 6516 6030 6534
rect 6012 6534 6030 6552
rect 6012 6552 6030 6570
rect 6012 6570 6030 6588
rect 6012 6588 6030 6606
rect 6012 6606 6030 6624
rect 6012 6624 6030 6642
rect 6012 6642 6030 6660
rect 6012 6660 6030 6678
rect 6012 6678 6030 6696
rect 6012 6696 6030 6714
rect 6012 6714 6030 6732
rect 6012 6732 6030 6750
rect 6012 6750 6030 6768
rect 6012 6768 6030 6786
rect 6012 6786 6030 6804
rect 6012 6804 6030 6822
rect 6012 6822 6030 6840
rect 6012 6840 6030 6858
rect 6012 6858 6030 6876
rect 6012 6876 6030 6894
rect 6012 6894 6030 6912
rect 6012 6912 6030 6930
rect 6012 6930 6030 6948
rect 6012 6948 6030 6966
rect 6012 6966 6030 6984
rect 6012 6984 6030 7002
rect 6012 7002 6030 7020
rect 6012 7020 6030 7038
rect 6012 7038 6030 7056
rect 6012 7056 6030 7074
rect 6012 7074 6030 7092
rect 6012 7092 6030 7110
rect 6012 7110 6030 7128
rect 6012 7128 6030 7146
rect 6012 7146 6030 7164
rect 6012 7164 6030 7182
rect 6012 7182 6030 7200
rect 6012 7200 6030 7218
rect 6012 7218 6030 7236
rect 6012 7236 6030 7254
rect 6012 7254 6030 7272
rect 6012 7272 6030 7290
rect 6012 7290 6030 7308
rect 6012 7308 6030 7326
rect 6012 7326 6030 7344
rect 6012 7344 6030 7362
rect 6012 7362 6030 7380
rect 6012 7380 6030 7398
rect 6012 7398 6030 7416
rect 6012 7416 6030 7434
rect 6012 7434 6030 7452
rect 6012 7452 6030 7470
rect 6012 7470 6030 7488
rect 6012 7488 6030 7506
rect 6012 7506 6030 7524
rect 6012 7524 6030 7542
rect 6012 7542 6030 7560
rect 6012 7560 6030 7578
rect 6012 7578 6030 7596
rect 6012 7596 6030 7614
rect 6012 7614 6030 7632
rect 6012 7632 6030 7650
rect 6012 7650 6030 7668
rect 6012 7668 6030 7686
rect 6012 7686 6030 7704
rect 6012 7704 6030 7722
rect 6012 7722 6030 7740
rect 6012 7740 6030 7758
rect 6012 7758 6030 7776
rect 6012 7776 6030 7794
rect 6012 7794 6030 7812
rect 6012 7812 6030 7830
rect 6012 7830 6030 7848
rect 6012 7848 6030 7866
rect 6012 7866 6030 7884
rect 6012 7884 6030 7902
rect 6012 7902 6030 7920
rect 6012 7920 6030 7938
rect 6012 7938 6030 7956
rect 6012 7956 6030 7974
rect 6012 7974 6030 7992
rect 6012 7992 6030 8010
rect 6012 8010 6030 8028
rect 6012 8028 6030 8046
rect 6012 8046 6030 8064
rect 6012 8064 6030 8082
rect 6012 8082 6030 8100
rect 6012 8100 6030 8118
rect 6012 8118 6030 8136
rect 6012 8136 6030 8154
rect 6012 8154 6030 8172
rect 6012 8172 6030 8190
rect 6012 8190 6030 8208
rect 6012 8208 6030 8226
rect 6012 8226 6030 8244
rect 6012 8244 6030 8262
rect 6012 8262 6030 8280
rect 6012 8280 6030 8298
rect 6012 8298 6030 8316
rect 6012 8316 6030 8334
rect 6012 8334 6030 8352
rect 6012 8352 6030 8370
rect 6012 8370 6030 8388
rect 6012 8388 6030 8406
rect 6012 8406 6030 8424
rect 6012 8424 6030 8442
rect 6012 8442 6030 8460
rect 6012 8460 6030 8478
rect 6012 8478 6030 8496
rect 6012 8496 6030 8514
rect 6012 8514 6030 8532
rect 6012 8532 6030 8550
rect 6012 8550 6030 8568
rect 6012 8568 6030 8586
rect 6012 8586 6030 8604
rect 6012 8604 6030 8622
rect 6012 8622 6030 8640
rect 6012 8640 6030 8658
rect 6012 8658 6030 8676
rect 6012 8676 6030 8694
rect 6012 8694 6030 8712
rect 6012 8712 6030 8730
rect 6012 8730 6030 8748
rect 6012 8748 6030 8766
rect 6012 8766 6030 8784
rect 6012 8784 6030 8802
rect 6012 8802 6030 8820
rect 6012 8820 6030 8838
rect 6012 8838 6030 8856
rect 6012 8856 6030 8874
rect 6012 8874 6030 8892
rect 6012 8892 6030 8910
rect 6012 8910 6030 8928
rect 6012 8928 6030 8946
rect 6012 8946 6030 8964
rect 6012 8964 6030 8982
rect 6012 8982 6030 9000
rect 6012 9000 6030 9018
rect 6012 9018 6030 9036
rect 6012 9036 6030 9054
rect 6012 9054 6030 9072
rect 6012 9072 6030 9090
rect 6012 9090 6030 9108
rect 6012 9108 6030 9126
rect 6012 9126 6030 9144
rect 6012 9144 6030 9162
rect 6012 9162 6030 9180
rect 6012 9180 6030 9198
rect 6012 9198 6030 9216
rect 6012 9216 6030 9234
rect 6012 9234 6030 9252
rect 6030 936 6048 954
rect 6030 954 6048 972
rect 6030 972 6048 990
rect 6030 990 6048 1008
rect 6030 1008 6048 1026
rect 6030 1026 6048 1044
rect 6030 1044 6048 1062
rect 6030 1062 6048 1080
rect 6030 1080 6048 1098
rect 6030 1098 6048 1116
rect 6030 1260 6048 1278
rect 6030 1278 6048 1296
rect 6030 1296 6048 1314
rect 6030 1314 6048 1332
rect 6030 1332 6048 1350
rect 6030 1350 6048 1368
rect 6030 1368 6048 1386
rect 6030 1386 6048 1404
rect 6030 1404 6048 1422
rect 6030 1422 6048 1440
rect 6030 1440 6048 1458
rect 6030 1458 6048 1476
rect 6030 1476 6048 1494
rect 6030 1494 6048 1512
rect 6030 1512 6048 1530
rect 6030 1530 6048 1548
rect 6030 1548 6048 1566
rect 6030 1566 6048 1584
rect 6030 1584 6048 1602
rect 6030 1602 6048 1620
rect 6030 1620 6048 1638
rect 6030 1638 6048 1656
rect 6030 1656 6048 1674
rect 6030 1674 6048 1692
rect 6030 1692 6048 1710
rect 6030 1710 6048 1728
rect 6030 1728 6048 1746
rect 6030 1746 6048 1764
rect 6030 1764 6048 1782
rect 6030 1782 6048 1800
rect 6030 1800 6048 1818
rect 6030 1818 6048 1836
rect 6030 1836 6048 1854
rect 6030 1854 6048 1872
rect 6030 1872 6048 1890
rect 6030 1890 6048 1908
rect 6030 1908 6048 1926
rect 6030 1926 6048 1944
rect 6030 1944 6048 1962
rect 6030 1962 6048 1980
rect 6030 1980 6048 1998
rect 6030 1998 6048 2016
rect 6030 2016 6048 2034
rect 6030 2034 6048 2052
rect 6030 2052 6048 2070
rect 6030 2070 6048 2088
rect 6030 2088 6048 2106
rect 6030 2106 6048 2124
rect 6030 2124 6048 2142
rect 6030 2142 6048 2160
rect 6030 2160 6048 2178
rect 6030 2178 6048 2196
rect 6030 2196 6048 2214
rect 6030 2214 6048 2232
rect 6030 2232 6048 2250
rect 6030 2250 6048 2268
rect 6030 2268 6048 2286
rect 6030 2286 6048 2304
rect 6030 2304 6048 2322
rect 6030 2322 6048 2340
rect 6030 2340 6048 2358
rect 6030 2358 6048 2376
rect 6030 2376 6048 2394
rect 6030 2394 6048 2412
rect 6030 2412 6048 2430
rect 6030 2430 6048 2448
rect 6030 2448 6048 2466
rect 6030 2466 6048 2484
rect 6030 2484 6048 2502
rect 6030 2502 6048 2520
rect 6030 2520 6048 2538
rect 6030 2538 6048 2556
rect 6030 2556 6048 2574
rect 6030 2574 6048 2592
rect 6030 2592 6048 2610
rect 6030 2610 6048 2628
rect 6030 2628 6048 2646
rect 6030 2646 6048 2664
rect 6030 2664 6048 2682
rect 6030 2682 6048 2700
rect 6030 2700 6048 2718
rect 6030 2718 6048 2736
rect 6030 2736 6048 2754
rect 6030 3006 6048 3024
rect 6030 3024 6048 3042
rect 6030 3042 6048 3060
rect 6030 3060 6048 3078
rect 6030 3078 6048 3096
rect 6030 3096 6048 3114
rect 6030 3114 6048 3132
rect 6030 3132 6048 3150
rect 6030 3150 6048 3168
rect 6030 3168 6048 3186
rect 6030 3186 6048 3204
rect 6030 3204 6048 3222
rect 6030 3222 6048 3240
rect 6030 3240 6048 3258
rect 6030 3258 6048 3276
rect 6030 3276 6048 3294
rect 6030 3294 6048 3312
rect 6030 3312 6048 3330
rect 6030 3330 6048 3348
rect 6030 3348 6048 3366
rect 6030 3366 6048 3384
rect 6030 3384 6048 3402
rect 6030 3402 6048 3420
rect 6030 3420 6048 3438
rect 6030 3438 6048 3456
rect 6030 3456 6048 3474
rect 6030 3474 6048 3492
rect 6030 3492 6048 3510
rect 6030 3510 6048 3528
rect 6030 3528 6048 3546
rect 6030 3546 6048 3564
rect 6030 3564 6048 3582
rect 6030 3582 6048 3600
rect 6030 3600 6048 3618
rect 6030 3618 6048 3636
rect 6030 3636 6048 3654
rect 6030 3654 6048 3672
rect 6030 3672 6048 3690
rect 6030 3690 6048 3708
rect 6030 3708 6048 3726
rect 6030 3726 6048 3744
rect 6030 3744 6048 3762
rect 6030 3762 6048 3780
rect 6030 3780 6048 3798
rect 6030 3798 6048 3816
rect 6030 3816 6048 3834
rect 6030 3834 6048 3852
rect 6030 3852 6048 3870
rect 6030 3870 6048 3888
rect 6030 3888 6048 3906
rect 6030 3906 6048 3924
rect 6030 3924 6048 3942
rect 6030 3942 6048 3960
rect 6030 3960 6048 3978
rect 6030 3978 6048 3996
rect 6030 3996 6048 4014
rect 6030 4014 6048 4032
rect 6030 4032 6048 4050
rect 6030 4050 6048 4068
rect 6030 4068 6048 4086
rect 6030 4086 6048 4104
rect 6030 4104 6048 4122
rect 6030 4122 6048 4140
rect 6030 4140 6048 4158
rect 6030 4158 6048 4176
rect 6030 4176 6048 4194
rect 6030 4194 6048 4212
rect 6030 4212 6048 4230
rect 6030 4230 6048 4248
rect 6030 4248 6048 4266
rect 6030 4266 6048 4284
rect 6030 4284 6048 4302
rect 6030 4302 6048 4320
rect 6030 4320 6048 4338
rect 6030 4338 6048 4356
rect 6030 4356 6048 4374
rect 6030 4374 6048 4392
rect 6030 4392 6048 4410
rect 6030 4410 6048 4428
rect 6030 4428 6048 4446
rect 6030 4446 6048 4464
rect 6030 4464 6048 4482
rect 6030 4482 6048 4500
rect 6030 4500 6048 4518
rect 6030 4518 6048 4536
rect 6030 4536 6048 4554
rect 6030 4554 6048 4572
rect 6030 4572 6048 4590
rect 6030 4590 6048 4608
rect 6030 4608 6048 4626
rect 6030 4626 6048 4644
rect 6030 4644 6048 4662
rect 6030 4662 6048 4680
rect 6030 4680 6048 4698
rect 6030 4698 6048 4716
rect 6030 4716 6048 4734
rect 6030 4734 6048 4752
rect 6030 4752 6048 4770
rect 6030 4770 6048 4788
rect 6030 4788 6048 4806
rect 6030 4806 6048 4824
rect 6030 4824 6048 4842
rect 6030 4842 6048 4860
rect 6030 4860 6048 4878
rect 6030 4878 6048 4896
rect 6030 4896 6048 4914
rect 6030 4914 6048 4932
rect 6030 4932 6048 4950
rect 6030 4950 6048 4968
rect 6030 4968 6048 4986
rect 6030 4986 6048 5004
rect 6030 5004 6048 5022
rect 6030 5022 6048 5040
rect 6030 5040 6048 5058
rect 6030 5058 6048 5076
rect 6030 5076 6048 5094
rect 6030 5094 6048 5112
rect 6030 5112 6048 5130
rect 6030 5130 6048 5148
rect 6030 5148 6048 5166
rect 6030 5166 6048 5184
rect 6030 5184 6048 5202
rect 6030 5202 6048 5220
rect 6030 5220 6048 5238
rect 6030 5238 6048 5256
rect 6030 5256 6048 5274
rect 6030 5274 6048 5292
rect 6030 5292 6048 5310
rect 6030 5310 6048 5328
rect 6030 5328 6048 5346
rect 6030 5346 6048 5364
rect 6030 5364 6048 5382
rect 6030 5382 6048 5400
rect 6030 5400 6048 5418
rect 6030 5670 6048 5688
rect 6030 5688 6048 5706
rect 6030 5706 6048 5724
rect 6030 5724 6048 5742
rect 6030 5742 6048 5760
rect 6030 5760 6048 5778
rect 6030 5778 6048 5796
rect 6030 5796 6048 5814
rect 6030 5814 6048 5832
rect 6030 5832 6048 5850
rect 6030 5850 6048 5868
rect 6030 5868 6048 5886
rect 6030 5886 6048 5904
rect 6030 5904 6048 5922
rect 6030 5922 6048 5940
rect 6030 5940 6048 5958
rect 6030 5958 6048 5976
rect 6030 5976 6048 5994
rect 6030 5994 6048 6012
rect 6030 6012 6048 6030
rect 6030 6030 6048 6048
rect 6030 6048 6048 6066
rect 6030 6066 6048 6084
rect 6030 6084 6048 6102
rect 6030 6102 6048 6120
rect 6030 6120 6048 6138
rect 6030 6138 6048 6156
rect 6030 6156 6048 6174
rect 6030 6174 6048 6192
rect 6030 6192 6048 6210
rect 6030 6210 6048 6228
rect 6030 6228 6048 6246
rect 6030 6246 6048 6264
rect 6030 6264 6048 6282
rect 6030 6282 6048 6300
rect 6030 6300 6048 6318
rect 6030 6318 6048 6336
rect 6030 6336 6048 6354
rect 6030 6354 6048 6372
rect 6030 6372 6048 6390
rect 6030 6390 6048 6408
rect 6030 6408 6048 6426
rect 6030 6426 6048 6444
rect 6030 6444 6048 6462
rect 6030 6462 6048 6480
rect 6030 6480 6048 6498
rect 6030 6498 6048 6516
rect 6030 6516 6048 6534
rect 6030 6534 6048 6552
rect 6030 6552 6048 6570
rect 6030 6570 6048 6588
rect 6030 6588 6048 6606
rect 6030 6606 6048 6624
rect 6030 6624 6048 6642
rect 6030 6642 6048 6660
rect 6030 6660 6048 6678
rect 6030 6678 6048 6696
rect 6030 6696 6048 6714
rect 6030 6714 6048 6732
rect 6030 6732 6048 6750
rect 6030 6750 6048 6768
rect 6030 6768 6048 6786
rect 6030 6786 6048 6804
rect 6030 6804 6048 6822
rect 6030 6822 6048 6840
rect 6030 6840 6048 6858
rect 6030 6858 6048 6876
rect 6030 6876 6048 6894
rect 6030 6894 6048 6912
rect 6030 6912 6048 6930
rect 6030 6930 6048 6948
rect 6030 6948 6048 6966
rect 6030 6966 6048 6984
rect 6030 6984 6048 7002
rect 6030 7002 6048 7020
rect 6030 7020 6048 7038
rect 6030 7038 6048 7056
rect 6030 7056 6048 7074
rect 6030 7074 6048 7092
rect 6030 7092 6048 7110
rect 6030 7110 6048 7128
rect 6030 7128 6048 7146
rect 6030 7146 6048 7164
rect 6030 7164 6048 7182
rect 6030 7182 6048 7200
rect 6030 7200 6048 7218
rect 6030 7218 6048 7236
rect 6030 7236 6048 7254
rect 6030 7254 6048 7272
rect 6030 7272 6048 7290
rect 6030 7290 6048 7308
rect 6030 7308 6048 7326
rect 6030 7326 6048 7344
rect 6030 7344 6048 7362
rect 6030 7362 6048 7380
rect 6030 7380 6048 7398
rect 6030 7398 6048 7416
rect 6030 7416 6048 7434
rect 6030 7434 6048 7452
rect 6030 7452 6048 7470
rect 6030 7470 6048 7488
rect 6030 7488 6048 7506
rect 6030 7506 6048 7524
rect 6030 7524 6048 7542
rect 6030 7542 6048 7560
rect 6030 7560 6048 7578
rect 6030 7578 6048 7596
rect 6030 7596 6048 7614
rect 6030 7614 6048 7632
rect 6030 7632 6048 7650
rect 6030 7650 6048 7668
rect 6030 7668 6048 7686
rect 6030 7686 6048 7704
rect 6030 7704 6048 7722
rect 6030 7722 6048 7740
rect 6030 7740 6048 7758
rect 6030 7758 6048 7776
rect 6030 7776 6048 7794
rect 6030 7794 6048 7812
rect 6030 7812 6048 7830
rect 6030 7830 6048 7848
rect 6030 7848 6048 7866
rect 6030 7866 6048 7884
rect 6030 7884 6048 7902
rect 6030 7902 6048 7920
rect 6030 7920 6048 7938
rect 6030 7938 6048 7956
rect 6030 7956 6048 7974
rect 6030 7974 6048 7992
rect 6030 7992 6048 8010
rect 6030 8010 6048 8028
rect 6030 8028 6048 8046
rect 6030 8046 6048 8064
rect 6030 8064 6048 8082
rect 6030 8082 6048 8100
rect 6030 8100 6048 8118
rect 6030 8118 6048 8136
rect 6030 8136 6048 8154
rect 6030 8154 6048 8172
rect 6030 8172 6048 8190
rect 6030 8190 6048 8208
rect 6030 8208 6048 8226
rect 6030 8226 6048 8244
rect 6030 8244 6048 8262
rect 6030 8262 6048 8280
rect 6030 8280 6048 8298
rect 6030 8298 6048 8316
rect 6030 8316 6048 8334
rect 6030 8334 6048 8352
rect 6030 8352 6048 8370
rect 6030 8370 6048 8388
rect 6030 8388 6048 8406
rect 6030 8406 6048 8424
rect 6030 8424 6048 8442
rect 6030 8442 6048 8460
rect 6030 8460 6048 8478
rect 6030 8478 6048 8496
rect 6030 8496 6048 8514
rect 6030 8514 6048 8532
rect 6030 8532 6048 8550
rect 6030 8550 6048 8568
rect 6030 8568 6048 8586
rect 6030 8586 6048 8604
rect 6030 8604 6048 8622
rect 6030 8622 6048 8640
rect 6030 8640 6048 8658
rect 6030 8658 6048 8676
rect 6030 8676 6048 8694
rect 6030 8694 6048 8712
rect 6030 8712 6048 8730
rect 6030 8730 6048 8748
rect 6030 8748 6048 8766
rect 6030 8766 6048 8784
rect 6030 8784 6048 8802
rect 6030 8802 6048 8820
rect 6030 8820 6048 8838
rect 6030 8838 6048 8856
rect 6030 8856 6048 8874
rect 6030 8874 6048 8892
rect 6030 8892 6048 8910
rect 6030 8910 6048 8928
rect 6030 8928 6048 8946
rect 6030 8946 6048 8964
rect 6030 8964 6048 8982
rect 6030 8982 6048 9000
rect 6030 9000 6048 9018
rect 6030 9018 6048 9036
rect 6030 9036 6048 9054
rect 6030 9054 6048 9072
rect 6030 9072 6048 9090
rect 6030 9090 6048 9108
rect 6030 9108 6048 9126
rect 6030 9126 6048 9144
rect 6030 9144 6048 9162
rect 6030 9162 6048 9180
rect 6030 9180 6048 9198
rect 6030 9198 6048 9216
rect 6030 9216 6048 9234
rect 6030 9234 6048 9252
rect 6030 9252 6048 9270
rect 6048 954 6066 972
rect 6048 972 6066 990
rect 6048 990 6066 1008
rect 6048 1008 6066 1026
rect 6048 1026 6066 1044
rect 6048 1044 6066 1062
rect 6048 1062 6066 1080
rect 6048 1080 6066 1098
rect 6048 1098 6066 1116
rect 6048 1278 6066 1296
rect 6048 1296 6066 1314
rect 6048 1314 6066 1332
rect 6048 1332 6066 1350
rect 6048 1350 6066 1368
rect 6048 1368 6066 1386
rect 6048 1386 6066 1404
rect 6048 1404 6066 1422
rect 6048 1422 6066 1440
rect 6048 1440 6066 1458
rect 6048 1458 6066 1476
rect 6048 1476 6066 1494
rect 6048 1494 6066 1512
rect 6048 1512 6066 1530
rect 6048 1530 6066 1548
rect 6048 1548 6066 1566
rect 6048 1566 6066 1584
rect 6048 1584 6066 1602
rect 6048 1602 6066 1620
rect 6048 1620 6066 1638
rect 6048 1638 6066 1656
rect 6048 1656 6066 1674
rect 6048 1674 6066 1692
rect 6048 1692 6066 1710
rect 6048 1710 6066 1728
rect 6048 1728 6066 1746
rect 6048 1746 6066 1764
rect 6048 1764 6066 1782
rect 6048 1782 6066 1800
rect 6048 1800 6066 1818
rect 6048 1818 6066 1836
rect 6048 1836 6066 1854
rect 6048 1854 6066 1872
rect 6048 1872 6066 1890
rect 6048 1890 6066 1908
rect 6048 1908 6066 1926
rect 6048 1926 6066 1944
rect 6048 1944 6066 1962
rect 6048 1962 6066 1980
rect 6048 1980 6066 1998
rect 6048 1998 6066 2016
rect 6048 2016 6066 2034
rect 6048 2034 6066 2052
rect 6048 2052 6066 2070
rect 6048 2070 6066 2088
rect 6048 2088 6066 2106
rect 6048 2106 6066 2124
rect 6048 2124 6066 2142
rect 6048 2142 6066 2160
rect 6048 2160 6066 2178
rect 6048 2178 6066 2196
rect 6048 2196 6066 2214
rect 6048 2214 6066 2232
rect 6048 2232 6066 2250
rect 6048 2250 6066 2268
rect 6048 2268 6066 2286
rect 6048 2286 6066 2304
rect 6048 2304 6066 2322
rect 6048 2322 6066 2340
rect 6048 2340 6066 2358
rect 6048 2358 6066 2376
rect 6048 2376 6066 2394
rect 6048 2394 6066 2412
rect 6048 2412 6066 2430
rect 6048 2430 6066 2448
rect 6048 2448 6066 2466
rect 6048 2466 6066 2484
rect 6048 2484 6066 2502
rect 6048 2502 6066 2520
rect 6048 2520 6066 2538
rect 6048 2538 6066 2556
rect 6048 2556 6066 2574
rect 6048 2574 6066 2592
rect 6048 2592 6066 2610
rect 6048 2610 6066 2628
rect 6048 2628 6066 2646
rect 6048 2646 6066 2664
rect 6048 2664 6066 2682
rect 6048 2682 6066 2700
rect 6048 2700 6066 2718
rect 6048 2718 6066 2736
rect 6048 2736 6066 2754
rect 6048 2754 6066 2772
rect 6048 3006 6066 3024
rect 6048 3024 6066 3042
rect 6048 3042 6066 3060
rect 6048 3060 6066 3078
rect 6048 3078 6066 3096
rect 6048 3096 6066 3114
rect 6048 3114 6066 3132
rect 6048 3132 6066 3150
rect 6048 3150 6066 3168
rect 6048 3168 6066 3186
rect 6048 3186 6066 3204
rect 6048 3204 6066 3222
rect 6048 3222 6066 3240
rect 6048 3240 6066 3258
rect 6048 3258 6066 3276
rect 6048 3276 6066 3294
rect 6048 3294 6066 3312
rect 6048 3312 6066 3330
rect 6048 3330 6066 3348
rect 6048 3348 6066 3366
rect 6048 3366 6066 3384
rect 6048 3384 6066 3402
rect 6048 3402 6066 3420
rect 6048 3420 6066 3438
rect 6048 3438 6066 3456
rect 6048 3456 6066 3474
rect 6048 3474 6066 3492
rect 6048 3492 6066 3510
rect 6048 3510 6066 3528
rect 6048 3528 6066 3546
rect 6048 3546 6066 3564
rect 6048 3564 6066 3582
rect 6048 3582 6066 3600
rect 6048 3600 6066 3618
rect 6048 3618 6066 3636
rect 6048 3636 6066 3654
rect 6048 3654 6066 3672
rect 6048 3672 6066 3690
rect 6048 3690 6066 3708
rect 6048 3708 6066 3726
rect 6048 3726 6066 3744
rect 6048 3744 6066 3762
rect 6048 3762 6066 3780
rect 6048 3780 6066 3798
rect 6048 3798 6066 3816
rect 6048 3816 6066 3834
rect 6048 3834 6066 3852
rect 6048 3852 6066 3870
rect 6048 3870 6066 3888
rect 6048 3888 6066 3906
rect 6048 3906 6066 3924
rect 6048 3924 6066 3942
rect 6048 3942 6066 3960
rect 6048 3960 6066 3978
rect 6048 3978 6066 3996
rect 6048 3996 6066 4014
rect 6048 4014 6066 4032
rect 6048 4032 6066 4050
rect 6048 4050 6066 4068
rect 6048 4068 6066 4086
rect 6048 4086 6066 4104
rect 6048 4104 6066 4122
rect 6048 4122 6066 4140
rect 6048 4140 6066 4158
rect 6048 4158 6066 4176
rect 6048 4176 6066 4194
rect 6048 4194 6066 4212
rect 6048 4212 6066 4230
rect 6048 4230 6066 4248
rect 6048 4248 6066 4266
rect 6048 4266 6066 4284
rect 6048 4284 6066 4302
rect 6048 4302 6066 4320
rect 6048 4320 6066 4338
rect 6048 4338 6066 4356
rect 6048 4356 6066 4374
rect 6048 4374 6066 4392
rect 6048 4392 6066 4410
rect 6048 4410 6066 4428
rect 6048 4428 6066 4446
rect 6048 4446 6066 4464
rect 6048 4464 6066 4482
rect 6048 4482 6066 4500
rect 6048 4500 6066 4518
rect 6048 4518 6066 4536
rect 6048 4536 6066 4554
rect 6048 4554 6066 4572
rect 6048 4572 6066 4590
rect 6048 4590 6066 4608
rect 6048 4608 6066 4626
rect 6048 4626 6066 4644
rect 6048 4644 6066 4662
rect 6048 4662 6066 4680
rect 6048 4680 6066 4698
rect 6048 4698 6066 4716
rect 6048 4716 6066 4734
rect 6048 4734 6066 4752
rect 6048 4752 6066 4770
rect 6048 4770 6066 4788
rect 6048 4788 6066 4806
rect 6048 4806 6066 4824
rect 6048 4824 6066 4842
rect 6048 4842 6066 4860
rect 6048 4860 6066 4878
rect 6048 4878 6066 4896
rect 6048 4896 6066 4914
rect 6048 4914 6066 4932
rect 6048 4932 6066 4950
rect 6048 4950 6066 4968
rect 6048 4968 6066 4986
rect 6048 4986 6066 5004
rect 6048 5004 6066 5022
rect 6048 5022 6066 5040
rect 6048 5040 6066 5058
rect 6048 5058 6066 5076
rect 6048 5076 6066 5094
rect 6048 5094 6066 5112
rect 6048 5112 6066 5130
rect 6048 5130 6066 5148
rect 6048 5148 6066 5166
rect 6048 5166 6066 5184
rect 6048 5184 6066 5202
rect 6048 5202 6066 5220
rect 6048 5220 6066 5238
rect 6048 5238 6066 5256
rect 6048 5256 6066 5274
rect 6048 5274 6066 5292
rect 6048 5292 6066 5310
rect 6048 5310 6066 5328
rect 6048 5328 6066 5346
rect 6048 5346 6066 5364
rect 6048 5364 6066 5382
rect 6048 5382 6066 5400
rect 6048 5400 6066 5418
rect 6048 5418 6066 5436
rect 6048 5688 6066 5706
rect 6048 5706 6066 5724
rect 6048 5724 6066 5742
rect 6048 5742 6066 5760
rect 6048 5760 6066 5778
rect 6048 5778 6066 5796
rect 6048 5796 6066 5814
rect 6048 5814 6066 5832
rect 6048 5832 6066 5850
rect 6048 5850 6066 5868
rect 6048 5868 6066 5886
rect 6048 5886 6066 5904
rect 6048 5904 6066 5922
rect 6048 5922 6066 5940
rect 6048 5940 6066 5958
rect 6048 5958 6066 5976
rect 6048 5976 6066 5994
rect 6048 5994 6066 6012
rect 6048 6012 6066 6030
rect 6048 6030 6066 6048
rect 6048 6048 6066 6066
rect 6048 6066 6066 6084
rect 6048 6084 6066 6102
rect 6048 6102 6066 6120
rect 6048 6120 6066 6138
rect 6048 6138 6066 6156
rect 6048 6156 6066 6174
rect 6048 6174 6066 6192
rect 6048 6192 6066 6210
rect 6048 6210 6066 6228
rect 6048 6228 6066 6246
rect 6048 6246 6066 6264
rect 6048 6264 6066 6282
rect 6048 6282 6066 6300
rect 6048 6300 6066 6318
rect 6048 6318 6066 6336
rect 6048 6336 6066 6354
rect 6048 6354 6066 6372
rect 6048 6372 6066 6390
rect 6048 6390 6066 6408
rect 6048 6408 6066 6426
rect 6048 6426 6066 6444
rect 6048 6444 6066 6462
rect 6048 6462 6066 6480
rect 6048 6480 6066 6498
rect 6048 6498 6066 6516
rect 6048 6516 6066 6534
rect 6048 6534 6066 6552
rect 6048 6552 6066 6570
rect 6048 6570 6066 6588
rect 6048 6588 6066 6606
rect 6048 6606 6066 6624
rect 6048 6624 6066 6642
rect 6048 6642 6066 6660
rect 6048 6660 6066 6678
rect 6048 6678 6066 6696
rect 6048 6696 6066 6714
rect 6048 6714 6066 6732
rect 6048 6732 6066 6750
rect 6048 6750 6066 6768
rect 6048 6768 6066 6786
rect 6048 6786 6066 6804
rect 6048 6804 6066 6822
rect 6048 6822 6066 6840
rect 6048 6840 6066 6858
rect 6048 6858 6066 6876
rect 6048 6876 6066 6894
rect 6048 6894 6066 6912
rect 6048 6912 6066 6930
rect 6048 6930 6066 6948
rect 6048 6948 6066 6966
rect 6048 6966 6066 6984
rect 6048 6984 6066 7002
rect 6048 7002 6066 7020
rect 6048 7020 6066 7038
rect 6048 7038 6066 7056
rect 6048 7056 6066 7074
rect 6048 7074 6066 7092
rect 6048 7092 6066 7110
rect 6048 7110 6066 7128
rect 6048 7128 6066 7146
rect 6048 7146 6066 7164
rect 6048 7164 6066 7182
rect 6048 7182 6066 7200
rect 6048 7200 6066 7218
rect 6048 7218 6066 7236
rect 6048 7236 6066 7254
rect 6048 7254 6066 7272
rect 6048 7272 6066 7290
rect 6048 7290 6066 7308
rect 6048 7308 6066 7326
rect 6048 7326 6066 7344
rect 6048 7344 6066 7362
rect 6048 7362 6066 7380
rect 6048 7380 6066 7398
rect 6048 7398 6066 7416
rect 6048 7416 6066 7434
rect 6048 7434 6066 7452
rect 6048 7452 6066 7470
rect 6048 7470 6066 7488
rect 6048 7488 6066 7506
rect 6048 7506 6066 7524
rect 6048 7524 6066 7542
rect 6048 7542 6066 7560
rect 6048 7560 6066 7578
rect 6048 7578 6066 7596
rect 6048 7596 6066 7614
rect 6048 7614 6066 7632
rect 6048 7632 6066 7650
rect 6048 7650 6066 7668
rect 6048 7668 6066 7686
rect 6048 7686 6066 7704
rect 6048 7704 6066 7722
rect 6048 7722 6066 7740
rect 6048 7740 6066 7758
rect 6048 7758 6066 7776
rect 6048 7776 6066 7794
rect 6048 7794 6066 7812
rect 6048 7812 6066 7830
rect 6048 7830 6066 7848
rect 6048 7848 6066 7866
rect 6048 7866 6066 7884
rect 6048 7884 6066 7902
rect 6048 7902 6066 7920
rect 6048 7920 6066 7938
rect 6048 7938 6066 7956
rect 6048 7956 6066 7974
rect 6048 7974 6066 7992
rect 6048 7992 6066 8010
rect 6048 8010 6066 8028
rect 6048 8028 6066 8046
rect 6048 8046 6066 8064
rect 6048 8064 6066 8082
rect 6048 8082 6066 8100
rect 6048 8100 6066 8118
rect 6048 8118 6066 8136
rect 6048 8136 6066 8154
rect 6048 8154 6066 8172
rect 6048 8172 6066 8190
rect 6048 8190 6066 8208
rect 6048 8208 6066 8226
rect 6048 8226 6066 8244
rect 6048 8244 6066 8262
rect 6048 8262 6066 8280
rect 6048 8280 6066 8298
rect 6048 8298 6066 8316
rect 6048 8316 6066 8334
rect 6048 8334 6066 8352
rect 6048 8352 6066 8370
rect 6048 8370 6066 8388
rect 6048 8388 6066 8406
rect 6048 8406 6066 8424
rect 6048 8424 6066 8442
rect 6048 8442 6066 8460
rect 6048 8460 6066 8478
rect 6048 8478 6066 8496
rect 6048 8496 6066 8514
rect 6048 8514 6066 8532
rect 6048 8532 6066 8550
rect 6048 8550 6066 8568
rect 6048 8568 6066 8586
rect 6048 8586 6066 8604
rect 6048 8604 6066 8622
rect 6048 8622 6066 8640
rect 6048 8640 6066 8658
rect 6048 8658 6066 8676
rect 6048 8676 6066 8694
rect 6048 8694 6066 8712
rect 6048 8712 6066 8730
rect 6048 8730 6066 8748
rect 6048 8748 6066 8766
rect 6048 8766 6066 8784
rect 6048 8784 6066 8802
rect 6048 8802 6066 8820
rect 6048 8820 6066 8838
rect 6048 8838 6066 8856
rect 6048 8856 6066 8874
rect 6048 8874 6066 8892
rect 6048 8892 6066 8910
rect 6048 8910 6066 8928
rect 6048 8928 6066 8946
rect 6048 8946 6066 8964
rect 6048 8964 6066 8982
rect 6048 8982 6066 9000
rect 6048 9000 6066 9018
rect 6048 9018 6066 9036
rect 6048 9036 6066 9054
rect 6048 9054 6066 9072
rect 6048 9072 6066 9090
rect 6048 9090 6066 9108
rect 6048 9108 6066 9126
rect 6048 9126 6066 9144
rect 6048 9144 6066 9162
rect 6048 9162 6066 9180
rect 6048 9180 6066 9198
rect 6048 9198 6066 9216
rect 6048 9216 6066 9234
rect 6048 9234 6066 9252
rect 6048 9252 6066 9270
rect 6048 9270 6066 9288
rect 6066 972 6084 990
rect 6066 990 6084 1008
rect 6066 1008 6084 1026
rect 6066 1026 6084 1044
rect 6066 1044 6084 1062
rect 6066 1062 6084 1080
rect 6066 1080 6084 1098
rect 6066 1098 6084 1116
rect 6066 1116 6084 1134
rect 6066 1278 6084 1296
rect 6066 1296 6084 1314
rect 6066 1314 6084 1332
rect 6066 1332 6084 1350
rect 6066 1350 6084 1368
rect 6066 1368 6084 1386
rect 6066 1386 6084 1404
rect 6066 1404 6084 1422
rect 6066 1422 6084 1440
rect 6066 1440 6084 1458
rect 6066 1458 6084 1476
rect 6066 1476 6084 1494
rect 6066 1494 6084 1512
rect 6066 1512 6084 1530
rect 6066 1530 6084 1548
rect 6066 1548 6084 1566
rect 6066 1566 6084 1584
rect 6066 1584 6084 1602
rect 6066 1602 6084 1620
rect 6066 1620 6084 1638
rect 6066 1638 6084 1656
rect 6066 1656 6084 1674
rect 6066 1674 6084 1692
rect 6066 1692 6084 1710
rect 6066 1710 6084 1728
rect 6066 1728 6084 1746
rect 6066 1746 6084 1764
rect 6066 1764 6084 1782
rect 6066 1782 6084 1800
rect 6066 1800 6084 1818
rect 6066 1818 6084 1836
rect 6066 1836 6084 1854
rect 6066 1854 6084 1872
rect 6066 1872 6084 1890
rect 6066 1890 6084 1908
rect 6066 1908 6084 1926
rect 6066 1926 6084 1944
rect 6066 1944 6084 1962
rect 6066 1962 6084 1980
rect 6066 1980 6084 1998
rect 6066 1998 6084 2016
rect 6066 2016 6084 2034
rect 6066 2034 6084 2052
rect 6066 2052 6084 2070
rect 6066 2070 6084 2088
rect 6066 2088 6084 2106
rect 6066 2106 6084 2124
rect 6066 2124 6084 2142
rect 6066 2142 6084 2160
rect 6066 2160 6084 2178
rect 6066 2178 6084 2196
rect 6066 2196 6084 2214
rect 6066 2214 6084 2232
rect 6066 2232 6084 2250
rect 6066 2250 6084 2268
rect 6066 2268 6084 2286
rect 6066 2286 6084 2304
rect 6066 2304 6084 2322
rect 6066 2322 6084 2340
rect 6066 2340 6084 2358
rect 6066 2358 6084 2376
rect 6066 2376 6084 2394
rect 6066 2394 6084 2412
rect 6066 2412 6084 2430
rect 6066 2430 6084 2448
rect 6066 2448 6084 2466
rect 6066 2466 6084 2484
rect 6066 2484 6084 2502
rect 6066 2502 6084 2520
rect 6066 2520 6084 2538
rect 6066 2538 6084 2556
rect 6066 2556 6084 2574
rect 6066 2574 6084 2592
rect 6066 2592 6084 2610
rect 6066 2610 6084 2628
rect 6066 2628 6084 2646
rect 6066 2646 6084 2664
rect 6066 2664 6084 2682
rect 6066 2682 6084 2700
rect 6066 2700 6084 2718
rect 6066 2718 6084 2736
rect 6066 2736 6084 2754
rect 6066 2754 6084 2772
rect 6066 3024 6084 3042
rect 6066 3042 6084 3060
rect 6066 3060 6084 3078
rect 6066 3078 6084 3096
rect 6066 3096 6084 3114
rect 6066 3114 6084 3132
rect 6066 3132 6084 3150
rect 6066 3150 6084 3168
rect 6066 3168 6084 3186
rect 6066 3186 6084 3204
rect 6066 3204 6084 3222
rect 6066 3222 6084 3240
rect 6066 3240 6084 3258
rect 6066 3258 6084 3276
rect 6066 3276 6084 3294
rect 6066 3294 6084 3312
rect 6066 3312 6084 3330
rect 6066 3330 6084 3348
rect 6066 3348 6084 3366
rect 6066 3366 6084 3384
rect 6066 3384 6084 3402
rect 6066 3402 6084 3420
rect 6066 3420 6084 3438
rect 6066 3438 6084 3456
rect 6066 3456 6084 3474
rect 6066 3474 6084 3492
rect 6066 3492 6084 3510
rect 6066 3510 6084 3528
rect 6066 3528 6084 3546
rect 6066 3546 6084 3564
rect 6066 3564 6084 3582
rect 6066 3582 6084 3600
rect 6066 3600 6084 3618
rect 6066 3618 6084 3636
rect 6066 3636 6084 3654
rect 6066 3654 6084 3672
rect 6066 3672 6084 3690
rect 6066 3690 6084 3708
rect 6066 3708 6084 3726
rect 6066 3726 6084 3744
rect 6066 3744 6084 3762
rect 6066 3762 6084 3780
rect 6066 3780 6084 3798
rect 6066 3798 6084 3816
rect 6066 3816 6084 3834
rect 6066 3834 6084 3852
rect 6066 3852 6084 3870
rect 6066 3870 6084 3888
rect 6066 3888 6084 3906
rect 6066 3906 6084 3924
rect 6066 3924 6084 3942
rect 6066 3942 6084 3960
rect 6066 3960 6084 3978
rect 6066 3978 6084 3996
rect 6066 3996 6084 4014
rect 6066 4014 6084 4032
rect 6066 4032 6084 4050
rect 6066 4050 6084 4068
rect 6066 4068 6084 4086
rect 6066 4086 6084 4104
rect 6066 4104 6084 4122
rect 6066 4122 6084 4140
rect 6066 4140 6084 4158
rect 6066 4158 6084 4176
rect 6066 4176 6084 4194
rect 6066 4194 6084 4212
rect 6066 4212 6084 4230
rect 6066 4230 6084 4248
rect 6066 4248 6084 4266
rect 6066 4266 6084 4284
rect 6066 4284 6084 4302
rect 6066 4302 6084 4320
rect 6066 4320 6084 4338
rect 6066 4338 6084 4356
rect 6066 4356 6084 4374
rect 6066 4374 6084 4392
rect 6066 4392 6084 4410
rect 6066 4410 6084 4428
rect 6066 4428 6084 4446
rect 6066 4446 6084 4464
rect 6066 4464 6084 4482
rect 6066 4482 6084 4500
rect 6066 4500 6084 4518
rect 6066 4518 6084 4536
rect 6066 4536 6084 4554
rect 6066 4554 6084 4572
rect 6066 4572 6084 4590
rect 6066 4590 6084 4608
rect 6066 4608 6084 4626
rect 6066 4626 6084 4644
rect 6066 4644 6084 4662
rect 6066 4662 6084 4680
rect 6066 4680 6084 4698
rect 6066 4698 6084 4716
rect 6066 4716 6084 4734
rect 6066 4734 6084 4752
rect 6066 4752 6084 4770
rect 6066 4770 6084 4788
rect 6066 4788 6084 4806
rect 6066 4806 6084 4824
rect 6066 4824 6084 4842
rect 6066 4842 6084 4860
rect 6066 4860 6084 4878
rect 6066 4878 6084 4896
rect 6066 4896 6084 4914
rect 6066 4914 6084 4932
rect 6066 4932 6084 4950
rect 6066 4950 6084 4968
rect 6066 4968 6084 4986
rect 6066 4986 6084 5004
rect 6066 5004 6084 5022
rect 6066 5022 6084 5040
rect 6066 5040 6084 5058
rect 6066 5058 6084 5076
rect 6066 5076 6084 5094
rect 6066 5094 6084 5112
rect 6066 5112 6084 5130
rect 6066 5130 6084 5148
rect 6066 5148 6084 5166
rect 6066 5166 6084 5184
rect 6066 5184 6084 5202
rect 6066 5202 6084 5220
rect 6066 5220 6084 5238
rect 6066 5238 6084 5256
rect 6066 5256 6084 5274
rect 6066 5274 6084 5292
rect 6066 5292 6084 5310
rect 6066 5310 6084 5328
rect 6066 5328 6084 5346
rect 6066 5346 6084 5364
rect 6066 5364 6084 5382
rect 6066 5382 6084 5400
rect 6066 5400 6084 5418
rect 6066 5418 6084 5436
rect 6066 5436 6084 5454
rect 6066 5706 6084 5724
rect 6066 5724 6084 5742
rect 6066 5742 6084 5760
rect 6066 5760 6084 5778
rect 6066 5778 6084 5796
rect 6066 5796 6084 5814
rect 6066 5814 6084 5832
rect 6066 5832 6084 5850
rect 6066 5850 6084 5868
rect 6066 5868 6084 5886
rect 6066 5886 6084 5904
rect 6066 5904 6084 5922
rect 6066 5922 6084 5940
rect 6066 5940 6084 5958
rect 6066 5958 6084 5976
rect 6066 5976 6084 5994
rect 6066 5994 6084 6012
rect 6066 6012 6084 6030
rect 6066 6030 6084 6048
rect 6066 6048 6084 6066
rect 6066 6066 6084 6084
rect 6066 6084 6084 6102
rect 6066 6102 6084 6120
rect 6066 6120 6084 6138
rect 6066 6138 6084 6156
rect 6066 6156 6084 6174
rect 6066 6174 6084 6192
rect 6066 6192 6084 6210
rect 6066 6210 6084 6228
rect 6066 6228 6084 6246
rect 6066 6246 6084 6264
rect 6066 6264 6084 6282
rect 6066 6282 6084 6300
rect 6066 6300 6084 6318
rect 6066 6318 6084 6336
rect 6066 6336 6084 6354
rect 6066 6354 6084 6372
rect 6066 6372 6084 6390
rect 6066 6390 6084 6408
rect 6066 6408 6084 6426
rect 6066 6426 6084 6444
rect 6066 6444 6084 6462
rect 6066 6462 6084 6480
rect 6066 6480 6084 6498
rect 6066 6498 6084 6516
rect 6066 6516 6084 6534
rect 6066 6534 6084 6552
rect 6066 6552 6084 6570
rect 6066 6570 6084 6588
rect 6066 6588 6084 6606
rect 6066 6606 6084 6624
rect 6066 6624 6084 6642
rect 6066 6642 6084 6660
rect 6066 6660 6084 6678
rect 6066 6678 6084 6696
rect 6066 6696 6084 6714
rect 6066 6714 6084 6732
rect 6066 6732 6084 6750
rect 6066 6750 6084 6768
rect 6066 6768 6084 6786
rect 6066 6786 6084 6804
rect 6066 6804 6084 6822
rect 6066 6822 6084 6840
rect 6066 6840 6084 6858
rect 6066 6858 6084 6876
rect 6066 6876 6084 6894
rect 6066 6894 6084 6912
rect 6066 6912 6084 6930
rect 6066 6930 6084 6948
rect 6066 6948 6084 6966
rect 6066 6966 6084 6984
rect 6066 6984 6084 7002
rect 6066 7002 6084 7020
rect 6066 7020 6084 7038
rect 6066 7038 6084 7056
rect 6066 7056 6084 7074
rect 6066 7074 6084 7092
rect 6066 7092 6084 7110
rect 6066 7110 6084 7128
rect 6066 7128 6084 7146
rect 6066 7146 6084 7164
rect 6066 7164 6084 7182
rect 6066 7182 6084 7200
rect 6066 7200 6084 7218
rect 6066 7218 6084 7236
rect 6066 7236 6084 7254
rect 6066 7254 6084 7272
rect 6066 7272 6084 7290
rect 6066 7290 6084 7308
rect 6066 7308 6084 7326
rect 6066 7326 6084 7344
rect 6066 7344 6084 7362
rect 6066 7362 6084 7380
rect 6066 7380 6084 7398
rect 6066 7398 6084 7416
rect 6066 7416 6084 7434
rect 6066 7434 6084 7452
rect 6066 7452 6084 7470
rect 6066 7470 6084 7488
rect 6066 7488 6084 7506
rect 6066 7506 6084 7524
rect 6066 7524 6084 7542
rect 6066 7542 6084 7560
rect 6066 7560 6084 7578
rect 6066 7578 6084 7596
rect 6066 7596 6084 7614
rect 6066 7614 6084 7632
rect 6066 7632 6084 7650
rect 6066 7650 6084 7668
rect 6066 7668 6084 7686
rect 6066 7686 6084 7704
rect 6066 7704 6084 7722
rect 6066 7722 6084 7740
rect 6066 7740 6084 7758
rect 6066 7758 6084 7776
rect 6066 7776 6084 7794
rect 6066 7794 6084 7812
rect 6066 7812 6084 7830
rect 6066 7830 6084 7848
rect 6066 7848 6084 7866
rect 6066 7866 6084 7884
rect 6066 7884 6084 7902
rect 6066 7902 6084 7920
rect 6066 7920 6084 7938
rect 6066 7938 6084 7956
rect 6066 7956 6084 7974
rect 6066 7974 6084 7992
rect 6066 7992 6084 8010
rect 6066 8010 6084 8028
rect 6066 8028 6084 8046
rect 6066 8046 6084 8064
rect 6066 8064 6084 8082
rect 6066 8082 6084 8100
rect 6066 8100 6084 8118
rect 6066 8118 6084 8136
rect 6066 8136 6084 8154
rect 6066 8154 6084 8172
rect 6066 8172 6084 8190
rect 6066 8190 6084 8208
rect 6066 8208 6084 8226
rect 6066 8226 6084 8244
rect 6066 8244 6084 8262
rect 6066 8262 6084 8280
rect 6066 8280 6084 8298
rect 6066 8298 6084 8316
rect 6066 8316 6084 8334
rect 6066 8334 6084 8352
rect 6066 8352 6084 8370
rect 6066 8370 6084 8388
rect 6066 8388 6084 8406
rect 6066 8406 6084 8424
rect 6066 8424 6084 8442
rect 6066 8442 6084 8460
rect 6066 8460 6084 8478
rect 6066 8478 6084 8496
rect 6066 8496 6084 8514
rect 6066 8514 6084 8532
rect 6066 8532 6084 8550
rect 6066 8550 6084 8568
rect 6066 8568 6084 8586
rect 6066 8586 6084 8604
rect 6066 8604 6084 8622
rect 6066 8622 6084 8640
rect 6066 8640 6084 8658
rect 6066 8658 6084 8676
rect 6066 8676 6084 8694
rect 6066 8694 6084 8712
rect 6066 8712 6084 8730
rect 6066 8730 6084 8748
rect 6066 8748 6084 8766
rect 6066 8766 6084 8784
rect 6066 8784 6084 8802
rect 6066 8802 6084 8820
rect 6066 8820 6084 8838
rect 6066 8838 6084 8856
rect 6066 8856 6084 8874
rect 6066 8874 6084 8892
rect 6066 8892 6084 8910
rect 6066 8910 6084 8928
rect 6066 8928 6084 8946
rect 6066 8946 6084 8964
rect 6066 8964 6084 8982
rect 6066 8982 6084 9000
rect 6066 9000 6084 9018
rect 6066 9018 6084 9036
rect 6066 9036 6084 9054
rect 6066 9054 6084 9072
rect 6066 9072 6084 9090
rect 6066 9090 6084 9108
rect 6066 9108 6084 9126
rect 6066 9126 6084 9144
rect 6066 9144 6084 9162
rect 6066 9162 6084 9180
rect 6066 9180 6084 9198
rect 6066 9198 6084 9216
rect 6066 9216 6084 9234
rect 6066 9234 6084 9252
rect 6066 9252 6084 9270
rect 6066 9270 6084 9288
rect 6066 9288 6084 9306
rect 6066 9306 6084 9324
rect 6084 990 6102 1008
rect 6084 1008 6102 1026
rect 6084 1026 6102 1044
rect 6084 1044 6102 1062
rect 6084 1062 6102 1080
rect 6084 1080 6102 1098
rect 6084 1098 6102 1116
rect 6084 1116 6102 1134
rect 6084 1278 6102 1296
rect 6084 1296 6102 1314
rect 6084 1314 6102 1332
rect 6084 1332 6102 1350
rect 6084 1350 6102 1368
rect 6084 1368 6102 1386
rect 6084 1386 6102 1404
rect 6084 1404 6102 1422
rect 6084 1422 6102 1440
rect 6084 1440 6102 1458
rect 6084 1458 6102 1476
rect 6084 1476 6102 1494
rect 6084 1494 6102 1512
rect 6084 1512 6102 1530
rect 6084 1530 6102 1548
rect 6084 1548 6102 1566
rect 6084 1566 6102 1584
rect 6084 1584 6102 1602
rect 6084 1602 6102 1620
rect 6084 1620 6102 1638
rect 6084 1638 6102 1656
rect 6084 1656 6102 1674
rect 6084 1674 6102 1692
rect 6084 1692 6102 1710
rect 6084 1710 6102 1728
rect 6084 1728 6102 1746
rect 6084 1746 6102 1764
rect 6084 1764 6102 1782
rect 6084 1782 6102 1800
rect 6084 1800 6102 1818
rect 6084 1818 6102 1836
rect 6084 1836 6102 1854
rect 6084 1854 6102 1872
rect 6084 1872 6102 1890
rect 6084 1890 6102 1908
rect 6084 1908 6102 1926
rect 6084 1926 6102 1944
rect 6084 1944 6102 1962
rect 6084 1962 6102 1980
rect 6084 1980 6102 1998
rect 6084 1998 6102 2016
rect 6084 2016 6102 2034
rect 6084 2034 6102 2052
rect 6084 2052 6102 2070
rect 6084 2070 6102 2088
rect 6084 2088 6102 2106
rect 6084 2106 6102 2124
rect 6084 2124 6102 2142
rect 6084 2142 6102 2160
rect 6084 2160 6102 2178
rect 6084 2178 6102 2196
rect 6084 2196 6102 2214
rect 6084 2214 6102 2232
rect 6084 2232 6102 2250
rect 6084 2250 6102 2268
rect 6084 2268 6102 2286
rect 6084 2286 6102 2304
rect 6084 2304 6102 2322
rect 6084 2322 6102 2340
rect 6084 2340 6102 2358
rect 6084 2358 6102 2376
rect 6084 2376 6102 2394
rect 6084 2394 6102 2412
rect 6084 2412 6102 2430
rect 6084 2430 6102 2448
rect 6084 2448 6102 2466
rect 6084 2466 6102 2484
rect 6084 2484 6102 2502
rect 6084 2502 6102 2520
rect 6084 2520 6102 2538
rect 6084 2538 6102 2556
rect 6084 2556 6102 2574
rect 6084 2574 6102 2592
rect 6084 2592 6102 2610
rect 6084 2610 6102 2628
rect 6084 2628 6102 2646
rect 6084 2646 6102 2664
rect 6084 2664 6102 2682
rect 6084 2682 6102 2700
rect 6084 2700 6102 2718
rect 6084 2718 6102 2736
rect 6084 2736 6102 2754
rect 6084 2754 6102 2772
rect 6084 2772 6102 2790
rect 6084 3024 6102 3042
rect 6084 3042 6102 3060
rect 6084 3060 6102 3078
rect 6084 3078 6102 3096
rect 6084 3096 6102 3114
rect 6084 3114 6102 3132
rect 6084 3132 6102 3150
rect 6084 3150 6102 3168
rect 6084 3168 6102 3186
rect 6084 3186 6102 3204
rect 6084 3204 6102 3222
rect 6084 3222 6102 3240
rect 6084 3240 6102 3258
rect 6084 3258 6102 3276
rect 6084 3276 6102 3294
rect 6084 3294 6102 3312
rect 6084 3312 6102 3330
rect 6084 3330 6102 3348
rect 6084 3348 6102 3366
rect 6084 3366 6102 3384
rect 6084 3384 6102 3402
rect 6084 3402 6102 3420
rect 6084 3420 6102 3438
rect 6084 3438 6102 3456
rect 6084 3456 6102 3474
rect 6084 3474 6102 3492
rect 6084 3492 6102 3510
rect 6084 3510 6102 3528
rect 6084 3528 6102 3546
rect 6084 3546 6102 3564
rect 6084 3564 6102 3582
rect 6084 3582 6102 3600
rect 6084 3600 6102 3618
rect 6084 3618 6102 3636
rect 6084 3636 6102 3654
rect 6084 3654 6102 3672
rect 6084 3672 6102 3690
rect 6084 3690 6102 3708
rect 6084 3708 6102 3726
rect 6084 3726 6102 3744
rect 6084 3744 6102 3762
rect 6084 3762 6102 3780
rect 6084 3780 6102 3798
rect 6084 3798 6102 3816
rect 6084 3816 6102 3834
rect 6084 3834 6102 3852
rect 6084 3852 6102 3870
rect 6084 3870 6102 3888
rect 6084 3888 6102 3906
rect 6084 3906 6102 3924
rect 6084 3924 6102 3942
rect 6084 3942 6102 3960
rect 6084 3960 6102 3978
rect 6084 3978 6102 3996
rect 6084 3996 6102 4014
rect 6084 4014 6102 4032
rect 6084 4032 6102 4050
rect 6084 4050 6102 4068
rect 6084 4068 6102 4086
rect 6084 4086 6102 4104
rect 6084 4104 6102 4122
rect 6084 4122 6102 4140
rect 6084 4140 6102 4158
rect 6084 4158 6102 4176
rect 6084 4176 6102 4194
rect 6084 4194 6102 4212
rect 6084 4212 6102 4230
rect 6084 4230 6102 4248
rect 6084 4248 6102 4266
rect 6084 4266 6102 4284
rect 6084 4284 6102 4302
rect 6084 4302 6102 4320
rect 6084 4320 6102 4338
rect 6084 4338 6102 4356
rect 6084 4356 6102 4374
rect 6084 4374 6102 4392
rect 6084 4392 6102 4410
rect 6084 4410 6102 4428
rect 6084 4428 6102 4446
rect 6084 4446 6102 4464
rect 6084 4464 6102 4482
rect 6084 4482 6102 4500
rect 6084 4500 6102 4518
rect 6084 4518 6102 4536
rect 6084 4536 6102 4554
rect 6084 4554 6102 4572
rect 6084 4572 6102 4590
rect 6084 4590 6102 4608
rect 6084 4608 6102 4626
rect 6084 4626 6102 4644
rect 6084 4644 6102 4662
rect 6084 4662 6102 4680
rect 6084 4680 6102 4698
rect 6084 4698 6102 4716
rect 6084 4716 6102 4734
rect 6084 4734 6102 4752
rect 6084 4752 6102 4770
rect 6084 4770 6102 4788
rect 6084 4788 6102 4806
rect 6084 4806 6102 4824
rect 6084 4824 6102 4842
rect 6084 4842 6102 4860
rect 6084 4860 6102 4878
rect 6084 4878 6102 4896
rect 6084 4896 6102 4914
rect 6084 4914 6102 4932
rect 6084 4932 6102 4950
rect 6084 4950 6102 4968
rect 6084 4968 6102 4986
rect 6084 4986 6102 5004
rect 6084 5004 6102 5022
rect 6084 5022 6102 5040
rect 6084 5040 6102 5058
rect 6084 5058 6102 5076
rect 6084 5076 6102 5094
rect 6084 5094 6102 5112
rect 6084 5112 6102 5130
rect 6084 5130 6102 5148
rect 6084 5148 6102 5166
rect 6084 5166 6102 5184
rect 6084 5184 6102 5202
rect 6084 5202 6102 5220
rect 6084 5220 6102 5238
rect 6084 5238 6102 5256
rect 6084 5256 6102 5274
rect 6084 5274 6102 5292
rect 6084 5292 6102 5310
rect 6084 5310 6102 5328
rect 6084 5328 6102 5346
rect 6084 5346 6102 5364
rect 6084 5364 6102 5382
rect 6084 5382 6102 5400
rect 6084 5400 6102 5418
rect 6084 5418 6102 5436
rect 6084 5436 6102 5454
rect 6084 5724 6102 5742
rect 6084 5742 6102 5760
rect 6084 5760 6102 5778
rect 6084 5778 6102 5796
rect 6084 5796 6102 5814
rect 6084 5814 6102 5832
rect 6084 5832 6102 5850
rect 6084 5850 6102 5868
rect 6084 5868 6102 5886
rect 6084 5886 6102 5904
rect 6084 5904 6102 5922
rect 6084 5922 6102 5940
rect 6084 5940 6102 5958
rect 6084 5958 6102 5976
rect 6084 5976 6102 5994
rect 6084 5994 6102 6012
rect 6084 6012 6102 6030
rect 6084 6030 6102 6048
rect 6084 6048 6102 6066
rect 6084 6066 6102 6084
rect 6084 6084 6102 6102
rect 6084 6102 6102 6120
rect 6084 6120 6102 6138
rect 6084 6138 6102 6156
rect 6084 6156 6102 6174
rect 6084 6174 6102 6192
rect 6084 6192 6102 6210
rect 6084 6210 6102 6228
rect 6084 6228 6102 6246
rect 6084 6246 6102 6264
rect 6084 6264 6102 6282
rect 6084 6282 6102 6300
rect 6084 6300 6102 6318
rect 6084 6318 6102 6336
rect 6084 6336 6102 6354
rect 6084 6354 6102 6372
rect 6084 6372 6102 6390
rect 6084 6390 6102 6408
rect 6084 6408 6102 6426
rect 6084 6426 6102 6444
rect 6084 6444 6102 6462
rect 6084 6462 6102 6480
rect 6084 6480 6102 6498
rect 6084 6498 6102 6516
rect 6084 6516 6102 6534
rect 6084 6534 6102 6552
rect 6084 6552 6102 6570
rect 6084 6570 6102 6588
rect 6084 6588 6102 6606
rect 6084 6606 6102 6624
rect 6084 6624 6102 6642
rect 6084 6642 6102 6660
rect 6084 6660 6102 6678
rect 6084 6678 6102 6696
rect 6084 6696 6102 6714
rect 6084 6714 6102 6732
rect 6084 6732 6102 6750
rect 6084 6750 6102 6768
rect 6084 6768 6102 6786
rect 6084 6786 6102 6804
rect 6084 6804 6102 6822
rect 6084 6822 6102 6840
rect 6084 6840 6102 6858
rect 6084 6858 6102 6876
rect 6084 6876 6102 6894
rect 6084 6894 6102 6912
rect 6084 6912 6102 6930
rect 6084 6930 6102 6948
rect 6084 6948 6102 6966
rect 6084 6966 6102 6984
rect 6084 6984 6102 7002
rect 6084 7002 6102 7020
rect 6084 7020 6102 7038
rect 6084 7038 6102 7056
rect 6084 7056 6102 7074
rect 6084 7074 6102 7092
rect 6084 7092 6102 7110
rect 6084 7110 6102 7128
rect 6084 7128 6102 7146
rect 6084 7146 6102 7164
rect 6084 7164 6102 7182
rect 6084 7182 6102 7200
rect 6084 7200 6102 7218
rect 6084 7218 6102 7236
rect 6084 7236 6102 7254
rect 6084 7254 6102 7272
rect 6084 7272 6102 7290
rect 6084 7290 6102 7308
rect 6084 7308 6102 7326
rect 6084 7326 6102 7344
rect 6084 7344 6102 7362
rect 6084 7362 6102 7380
rect 6084 7380 6102 7398
rect 6084 7398 6102 7416
rect 6084 7416 6102 7434
rect 6084 7434 6102 7452
rect 6084 7452 6102 7470
rect 6084 7470 6102 7488
rect 6084 7488 6102 7506
rect 6084 7506 6102 7524
rect 6084 7524 6102 7542
rect 6084 7542 6102 7560
rect 6084 7560 6102 7578
rect 6084 7578 6102 7596
rect 6084 7596 6102 7614
rect 6084 7614 6102 7632
rect 6084 7632 6102 7650
rect 6084 7650 6102 7668
rect 6084 7668 6102 7686
rect 6084 7686 6102 7704
rect 6084 7704 6102 7722
rect 6084 7722 6102 7740
rect 6084 7740 6102 7758
rect 6084 7758 6102 7776
rect 6084 7776 6102 7794
rect 6084 7794 6102 7812
rect 6084 7812 6102 7830
rect 6084 7830 6102 7848
rect 6084 7848 6102 7866
rect 6084 7866 6102 7884
rect 6084 7884 6102 7902
rect 6084 7902 6102 7920
rect 6084 7920 6102 7938
rect 6084 7938 6102 7956
rect 6084 7956 6102 7974
rect 6084 7974 6102 7992
rect 6084 7992 6102 8010
rect 6084 8010 6102 8028
rect 6084 8028 6102 8046
rect 6084 8046 6102 8064
rect 6084 8064 6102 8082
rect 6084 8082 6102 8100
rect 6084 8100 6102 8118
rect 6084 8118 6102 8136
rect 6084 8136 6102 8154
rect 6084 8154 6102 8172
rect 6084 8172 6102 8190
rect 6084 8190 6102 8208
rect 6084 8208 6102 8226
rect 6084 8226 6102 8244
rect 6084 8244 6102 8262
rect 6084 8262 6102 8280
rect 6084 8280 6102 8298
rect 6084 8298 6102 8316
rect 6084 8316 6102 8334
rect 6084 8334 6102 8352
rect 6084 8352 6102 8370
rect 6084 8370 6102 8388
rect 6084 8388 6102 8406
rect 6084 8406 6102 8424
rect 6084 8424 6102 8442
rect 6084 8442 6102 8460
rect 6084 8460 6102 8478
rect 6084 8478 6102 8496
rect 6084 8496 6102 8514
rect 6084 8514 6102 8532
rect 6084 8532 6102 8550
rect 6084 8550 6102 8568
rect 6084 8568 6102 8586
rect 6084 8586 6102 8604
rect 6084 8604 6102 8622
rect 6084 8622 6102 8640
rect 6084 8640 6102 8658
rect 6084 8658 6102 8676
rect 6084 8676 6102 8694
rect 6084 8694 6102 8712
rect 6084 8712 6102 8730
rect 6084 8730 6102 8748
rect 6084 8748 6102 8766
rect 6084 8766 6102 8784
rect 6084 8784 6102 8802
rect 6084 8802 6102 8820
rect 6084 8820 6102 8838
rect 6084 8838 6102 8856
rect 6084 8856 6102 8874
rect 6084 8874 6102 8892
rect 6084 8892 6102 8910
rect 6084 8910 6102 8928
rect 6084 8928 6102 8946
rect 6084 8946 6102 8964
rect 6084 8964 6102 8982
rect 6084 8982 6102 9000
rect 6084 9000 6102 9018
rect 6084 9018 6102 9036
rect 6084 9036 6102 9054
rect 6084 9054 6102 9072
rect 6084 9072 6102 9090
rect 6084 9090 6102 9108
rect 6084 9108 6102 9126
rect 6084 9126 6102 9144
rect 6084 9144 6102 9162
rect 6084 9162 6102 9180
rect 6084 9180 6102 9198
rect 6084 9198 6102 9216
rect 6084 9216 6102 9234
rect 6084 9234 6102 9252
rect 6084 9252 6102 9270
rect 6084 9270 6102 9288
rect 6084 9288 6102 9306
rect 6084 9306 6102 9324
rect 6084 9324 6102 9342
rect 6102 1008 6120 1026
rect 6102 1026 6120 1044
rect 6102 1044 6120 1062
rect 6102 1062 6120 1080
rect 6102 1080 6120 1098
rect 6102 1098 6120 1116
rect 6102 1116 6120 1134
rect 6102 1134 6120 1152
rect 6102 1296 6120 1314
rect 6102 1314 6120 1332
rect 6102 1332 6120 1350
rect 6102 1350 6120 1368
rect 6102 1368 6120 1386
rect 6102 1386 6120 1404
rect 6102 1404 6120 1422
rect 6102 1422 6120 1440
rect 6102 1440 6120 1458
rect 6102 1458 6120 1476
rect 6102 1476 6120 1494
rect 6102 1494 6120 1512
rect 6102 1512 6120 1530
rect 6102 1530 6120 1548
rect 6102 1548 6120 1566
rect 6102 1566 6120 1584
rect 6102 1584 6120 1602
rect 6102 1602 6120 1620
rect 6102 1620 6120 1638
rect 6102 1638 6120 1656
rect 6102 1656 6120 1674
rect 6102 1674 6120 1692
rect 6102 1692 6120 1710
rect 6102 1710 6120 1728
rect 6102 1728 6120 1746
rect 6102 1746 6120 1764
rect 6102 1764 6120 1782
rect 6102 1782 6120 1800
rect 6102 1800 6120 1818
rect 6102 1818 6120 1836
rect 6102 1836 6120 1854
rect 6102 1854 6120 1872
rect 6102 1872 6120 1890
rect 6102 1890 6120 1908
rect 6102 1908 6120 1926
rect 6102 1926 6120 1944
rect 6102 1944 6120 1962
rect 6102 1962 6120 1980
rect 6102 1980 6120 1998
rect 6102 1998 6120 2016
rect 6102 2016 6120 2034
rect 6102 2034 6120 2052
rect 6102 2052 6120 2070
rect 6102 2070 6120 2088
rect 6102 2088 6120 2106
rect 6102 2106 6120 2124
rect 6102 2124 6120 2142
rect 6102 2142 6120 2160
rect 6102 2160 6120 2178
rect 6102 2178 6120 2196
rect 6102 2196 6120 2214
rect 6102 2214 6120 2232
rect 6102 2232 6120 2250
rect 6102 2250 6120 2268
rect 6102 2268 6120 2286
rect 6102 2286 6120 2304
rect 6102 2304 6120 2322
rect 6102 2322 6120 2340
rect 6102 2340 6120 2358
rect 6102 2358 6120 2376
rect 6102 2376 6120 2394
rect 6102 2394 6120 2412
rect 6102 2412 6120 2430
rect 6102 2430 6120 2448
rect 6102 2448 6120 2466
rect 6102 2466 6120 2484
rect 6102 2484 6120 2502
rect 6102 2502 6120 2520
rect 6102 2520 6120 2538
rect 6102 2538 6120 2556
rect 6102 2556 6120 2574
rect 6102 2574 6120 2592
rect 6102 2592 6120 2610
rect 6102 2610 6120 2628
rect 6102 2628 6120 2646
rect 6102 2646 6120 2664
rect 6102 2664 6120 2682
rect 6102 2682 6120 2700
rect 6102 2700 6120 2718
rect 6102 2718 6120 2736
rect 6102 2736 6120 2754
rect 6102 2754 6120 2772
rect 6102 2772 6120 2790
rect 6102 3042 6120 3060
rect 6102 3060 6120 3078
rect 6102 3078 6120 3096
rect 6102 3096 6120 3114
rect 6102 3114 6120 3132
rect 6102 3132 6120 3150
rect 6102 3150 6120 3168
rect 6102 3168 6120 3186
rect 6102 3186 6120 3204
rect 6102 3204 6120 3222
rect 6102 3222 6120 3240
rect 6102 3240 6120 3258
rect 6102 3258 6120 3276
rect 6102 3276 6120 3294
rect 6102 3294 6120 3312
rect 6102 3312 6120 3330
rect 6102 3330 6120 3348
rect 6102 3348 6120 3366
rect 6102 3366 6120 3384
rect 6102 3384 6120 3402
rect 6102 3402 6120 3420
rect 6102 3420 6120 3438
rect 6102 3438 6120 3456
rect 6102 3456 6120 3474
rect 6102 3474 6120 3492
rect 6102 3492 6120 3510
rect 6102 3510 6120 3528
rect 6102 3528 6120 3546
rect 6102 3546 6120 3564
rect 6102 3564 6120 3582
rect 6102 3582 6120 3600
rect 6102 3600 6120 3618
rect 6102 3618 6120 3636
rect 6102 3636 6120 3654
rect 6102 3654 6120 3672
rect 6102 3672 6120 3690
rect 6102 3690 6120 3708
rect 6102 3708 6120 3726
rect 6102 3726 6120 3744
rect 6102 3744 6120 3762
rect 6102 3762 6120 3780
rect 6102 3780 6120 3798
rect 6102 3798 6120 3816
rect 6102 3816 6120 3834
rect 6102 3834 6120 3852
rect 6102 3852 6120 3870
rect 6102 3870 6120 3888
rect 6102 3888 6120 3906
rect 6102 3906 6120 3924
rect 6102 3924 6120 3942
rect 6102 3942 6120 3960
rect 6102 3960 6120 3978
rect 6102 3978 6120 3996
rect 6102 3996 6120 4014
rect 6102 4014 6120 4032
rect 6102 4032 6120 4050
rect 6102 4050 6120 4068
rect 6102 4068 6120 4086
rect 6102 4086 6120 4104
rect 6102 4104 6120 4122
rect 6102 4122 6120 4140
rect 6102 4140 6120 4158
rect 6102 4158 6120 4176
rect 6102 4176 6120 4194
rect 6102 4194 6120 4212
rect 6102 4212 6120 4230
rect 6102 4230 6120 4248
rect 6102 4248 6120 4266
rect 6102 4266 6120 4284
rect 6102 4284 6120 4302
rect 6102 4302 6120 4320
rect 6102 4320 6120 4338
rect 6102 4338 6120 4356
rect 6102 4356 6120 4374
rect 6102 4374 6120 4392
rect 6102 4392 6120 4410
rect 6102 4410 6120 4428
rect 6102 4428 6120 4446
rect 6102 4446 6120 4464
rect 6102 4464 6120 4482
rect 6102 4482 6120 4500
rect 6102 4500 6120 4518
rect 6102 4518 6120 4536
rect 6102 4536 6120 4554
rect 6102 4554 6120 4572
rect 6102 4572 6120 4590
rect 6102 4590 6120 4608
rect 6102 4608 6120 4626
rect 6102 4626 6120 4644
rect 6102 4644 6120 4662
rect 6102 4662 6120 4680
rect 6102 4680 6120 4698
rect 6102 4698 6120 4716
rect 6102 4716 6120 4734
rect 6102 4734 6120 4752
rect 6102 4752 6120 4770
rect 6102 4770 6120 4788
rect 6102 4788 6120 4806
rect 6102 4806 6120 4824
rect 6102 4824 6120 4842
rect 6102 4842 6120 4860
rect 6102 4860 6120 4878
rect 6102 4878 6120 4896
rect 6102 4896 6120 4914
rect 6102 4914 6120 4932
rect 6102 4932 6120 4950
rect 6102 4950 6120 4968
rect 6102 4968 6120 4986
rect 6102 4986 6120 5004
rect 6102 5004 6120 5022
rect 6102 5022 6120 5040
rect 6102 5040 6120 5058
rect 6102 5058 6120 5076
rect 6102 5076 6120 5094
rect 6102 5094 6120 5112
rect 6102 5112 6120 5130
rect 6102 5130 6120 5148
rect 6102 5148 6120 5166
rect 6102 5166 6120 5184
rect 6102 5184 6120 5202
rect 6102 5202 6120 5220
rect 6102 5220 6120 5238
rect 6102 5238 6120 5256
rect 6102 5256 6120 5274
rect 6102 5274 6120 5292
rect 6102 5292 6120 5310
rect 6102 5310 6120 5328
rect 6102 5328 6120 5346
rect 6102 5346 6120 5364
rect 6102 5364 6120 5382
rect 6102 5382 6120 5400
rect 6102 5400 6120 5418
rect 6102 5418 6120 5436
rect 6102 5436 6120 5454
rect 6102 5454 6120 5472
rect 6102 5742 6120 5760
rect 6102 5760 6120 5778
rect 6102 5778 6120 5796
rect 6102 5796 6120 5814
rect 6102 5814 6120 5832
rect 6102 5832 6120 5850
rect 6102 5850 6120 5868
rect 6102 5868 6120 5886
rect 6102 5886 6120 5904
rect 6102 5904 6120 5922
rect 6102 5922 6120 5940
rect 6102 5940 6120 5958
rect 6102 5958 6120 5976
rect 6102 5976 6120 5994
rect 6102 5994 6120 6012
rect 6102 6012 6120 6030
rect 6102 6030 6120 6048
rect 6102 6048 6120 6066
rect 6102 6066 6120 6084
rect 6102 6084 6120 6102
rect 6102 6102 6120 6120
rect 6102 6120 6120 6138
rect 6102 6138 6120 6156
rect 6102 6156 6120 6174
rect 6102 6174 6120 6192
rect 6102 6192 6120 6210
rect 6102 6210 6120 6228
rect 6102 6228 6120 6246
rect 6102 6246 6120 6264
rect 6102 6264 6120 6282
rect 6102 6282 6120 6300
rect 6102 6300 6120 6318
rect 6102 6318 6120 6336
rect 6102 6336 6120 6354
rect 6102 6354 6120 6372
rect 6102 6372 6120 6390
rect 6102 6390 6120 6408
rect 6102 6408 6120 6426
rect 6102 6426 6120 6444
rect 6102 6444 6120 6462
rect 6102 6462 6120 6480
rect 6102 6480 6120 6498
rect 6102 6498 6120 6516
rect 6102 6516 6120 6534
rect 6102 6534 6120 6552
rect 6102 6552 6120 6570
rect 6102 6570 6120 6588
rect 6102 6588 6120 6606
rect 6102 6606 6120 6624
rect 6102 6624 6120 6642
rect 6102 6642 6120 6660
rect 6102 6660 6120 6678
rect 6102 6678 6120 6696
rect 6102 6696 6120 6714
rect 6102 6714 6120 6732
rect 6102 6732 6120 6750
rect 6102 6750 6120 6768
rect 6102 6768 6120 6786
rect 6102 6786 6120 6804
rect 6102 6804 6120 6822
rect 6102 6822 6120 6840
rect 6102 6840 6120 6858
rect 6102 6858 6120 6876
rect 6102 6876 6120 6894
rect 6102 6894 6120 6912
rect 6102 6912 6120 6930
rect 6102 6930 6120 6948
rect 6102 6948 6120 6966
rect 6102 6966 6120 6984
rect 6102 6984 6120 7002
rect 6102 7002 6120 7020
rect 6102 7020 6120 7038
rect 6102 7038 6120 7056
rect 6102 7056 6120 7074
rect 6102 7074 6120 7092
rect 6102 7092 6120 7110
rect 6102 7110 6120 7128
rect 6102 7128 6120 7146
rect 6102 7146 6120 7164
rect 6102 7164 6120 7182
rect 6102 7182 6120 7200
rect 6102 7200 6120 7218
rect 6102 7218 6120 7236
rect 6102 7236 6120 7254
rect 6102 7254 6120 7272
rect 6102 7272 6120 7290
rect 6102 7290 6120 7308
rect 6102 7308 6120 7326
rect 6102 7326 6120 7344
rect 6102 7344 6120 7362
rect 6102 7362 6120 7380
rect 6102 7380 6120 7398
rect 6102 7398 6120 7416
rect 6102 7416 6120 7434
rect 6102 7434 6120 7452
rect 6102 7452 6120 7470
rect 6102 7470 6120 7488
rect 6102 7488 6120 7506
rect 6102 7506 6120 7524
rect 6102 7524 6120 7542
rect 6102 7542 6120 7560
rect 6102 7560 6120 7578
rect 6102 7578 6120 7596
rect 6102 7596 6120 7614
rect 6102 7614 6120 7632
rect 6102 7632 6120 7650
rect 6102 7650 6120 7668
rect 6102 7668 6120 7686
rect 6102 7686 6120 7704
rect 6102 7704 6120 7722
rect 6102 7722 6120 7740
rect 6102 7740 6120 7758
rect 6102 7758 6120 7776
rect 6102 7776 6120 7794
rect 6102 7794 6120 7812
rect 6102 7812 6120 7830
rect 6102 7830 6120 7848
rect 6102 7848 6120 7866
rect 6102 7866 6120 7884
rect 6102 7884 6120 7902
rect 6102 7902 6120 7920
rect 6102 7920 6120 7938
rect 6102 7938 6120 7956
rect 6102 7956 6120 7974
rect 6102 7974 6120 7992
rect 6102 7992 6120 8010
rect 6102 8010 6120 8028
rect 6102 8028 6120 8046
rect 6102 8046 6120 8064
rect 6102 8064 6120 8082
rect 6102 8082 6120 8100
rect 6102 8100 6120 8118
rect 6102 8118 6120 8136
rect 6102 8136 6120 8154
rect 6102 8154 6120 8172
rect 6102 8172 6120 8190
rect 6102 8190 6120 8208
rect 6102 8208 6120 8226
rect 6102 8226 6120 8244
rect 6102 8244 6120 8262
rect 6102 8262 6120 8280
rect 6102 8280 6120 8298
rect 6102 8298 6120 8316
rect 6102 8316 6120 8334
rect 6102 8334 6120 8352
rect 6102 8352 6120 8370
rect 6102 8370 6120 8388
rect 6102 8388 6120 8406
rect 6102 8406 6120 8424
rect 6102 8424 6120 8442
rect 6102 8442 6120 8460
rect 6102 8460 6120 8478
rect 6102 8478 6120 8496
rect 6102 8496 6120 8514
rect 6102 8514 6120 8532
rect 6102 8532 6120 8550
rect 6102 8550 6120 8568
rect 6102 8568 6120 8586
rect 6102 8586 6120 8604
rect 6102 8604 6120 8622
rect 6102 8622 6120 8640
rect 6102 8640 6120 8658
rect 6102 8658 6120 8676
rect 6102 8676 6120 8694
rect 6102 8694 6120 8712
rect 6102 8712 6120 8730
rect 6102 8730 6120 8748
rect 6102 8748 6120 8766
rect 6102 8766 6120 8784
rect 6102 8784 6120 8802
rect 6102 8802 6120 8820
rect 6102 8820 6120 8838
rect 6102 8838 6120 8856
rect 6102 8856 6120 8874
rect 6102 8874 6120 8892
rect 6102 8892 6120 8910
rect 6102 8910 6120 8928
rect 6102 8928 6120 8946
rect 6102 8946 6120 8964
rect 6102 8964 6120 8982
rect 6102 8982 6120 9000
rect 6102 9000 6120 9018
rect 6102 9018 6120 9036
rect 6102 9036 6120 9054
rect 6102 9054 6120 9072
rect 6102 9072 6120 9090
rect 6102 9090 6120 9108
rect 6102 9108 6120 9126
rect 6102 9126 6120 9144
rect 6102 9144 6120 9162
rect 6102 9162 6120 9180
rect 6102 9180 6120 9198
rect 6102 9198 6120 9216
rect 6102 9216 6120 9234
rect 6102 9234 6120 9252
rect 6102 9252 6120 9270
rect 6102 9270 6120 9288
rect 6102 9288 6120 9306
rect 6102 9306 6120 9324
rect 6102 9324 6120 9342
rect 6102 9342 6120 9360
rect 6120 1026 6138 1044
rect 6120 1044 6138 1062
rect 6120 1062 6138 1080
rect 6120 1080 6138 1098
rect 6120 1098 6138 1116
rect 6120 1116 6138 1134
rect 6120 1134 6138 1152
rect 6120 1296 6138 1314
rect 6120 1314 6138 1332
rect 6120 1332 6138 1350
rect 6120 1350 6138 1368
rect 6120 1368 6138 1386
rect 6120 1386 6138 1404
rect 6120 1404 6138 1422
rect 6120 1422 6138 1440
rect 6120 1440 6138 1458
rect 6120 1458 6138 1476
rect 6120 1476 6138 1494
rect 6120 1494 6138 1512
rect 6120 1512 6138 1530
rect 6120 1530 6138 1548
rect 6120 1548 6138 1566
rect 6120 1566 6138 1584
rect 6120 1584 6138 1602
rect 6120 1602 6138 1620
rect 6120 1620 6138 1638
rect 6120 1638 6138 1656
rect 6120 1656 6138 1674
rect 6120 1674 6138 1692
rect 6120 1692 6138 1710
rect 6120 1710 6138 1728
rect 6120 1728 6138 1746
rect 6120 1746 6138 1764
rect 6120 1764 6138 1782
rect 6120 1782 6138 1800
rect 6120 1800 6138 1818
rect 6120 1818 6138 1836
rect 6120 1836 6138 1854
rect 6120 1854 6138 1872
rect 6120 1872 6138 1890
rect 6120 1890 6138 1908
rect 6120 1908 6138 1926
rect 6120 1926 6138 1944
rect 6120 1944 6138 1962
rect 6120 1962 6138 1980
rect 6120 1980 6138 1998
rect 6120 1998 6138 2016
rect 6120 2016 6138 2034
rect 6120 2034 6138 2052
rect 6120 2052 6138 2070
rect 6120 2070 6138 2088
rect 6120 2088 6138 2106
rect 6120 2106 6138 2124
rect 6120 2124 6138 2142
rect 6120 2142 6138 2160
rect 6120 2160 6138 2178
rect 6120 2178 6138 2196
rect 6120 2196 6138 2214
rect 6120 2214 6138 2232
rect 6120 2232 6138 2250
rect 6120 2250 6138 2268
rect 6120 2268 6138 2286
rect 6120 2286 6138 2304
rect 6120 2304 6138 2322
rect 6120 2322 6138 2340
rect 6120 2340 6138 2358
rect 6120 2358 6138 2376
rect 6120 2376 6138 2394
rect 6120 2394 6138 2412
rect 6120 2412 6138 2430
rect 6120 2430 6138 2448
rect 6120 2448 6138 2466
rect 6120 2466 6138 2484
rect 6120 2484 6138 2502
rect 6120 2502 6138 2520
rect 6120 2520 6138 2538
rect 6120 2538 6138 2556
rect 6120 2556 6138 2574
rect 6120 2574 6138 2592
rect 6120 2592 6138 2610
rect 6120 2610 6138 2628
rect 6120 2628 6138 2646
rect 6120 2646 6138 2664
rect 6120 2664 6138 2682
rect 6120 2682 6138 2700
rect 6120 2700 6138 2718
rect 6120 2718 6138 2736
rect 6120 2736 6138 2754
rect 6120 2754 6138 2772
rect 6120 2772 6138 2790
rect 6120 3042 6138 3060
rect 6120 3060 6138 3078
rect 6120 3078 6138 3096
rect 6120 3096 6138 3114
rect 6120 3114 6138 3132
rect 6120 3132 6138 3150
rect 6120 3150 6138 3168
rect 6120 3168 6138 3186
rect 6120 3186 6138 3204
rect 6120 3204 6138 3222
rect 6120 3222 6138 3240
rect 6120 3240 6138 3258
rect 6120 3258 6138 3276
rect 6120 3276 6138 3294
rect 6120 3294 6138 3312
rect 6120 3312 6138 3330
rect 6120 3330 6138 3348
rect 6120 3348 6138 3366
rect 6120 3366 6138 3384
rect 6120 3384 6138 3402
rect 6120 3402 6138 3420
rect 6120 3420 6138 3438
rect 6120 3438 6138 3456
rect 6120 3456 6138 3474
rect 6120 3474 6138 3492
rect 6120 3492 6138 3510
rect 6120 3510 6138 3528
rect 6120 3528 6138 3546
rect 6120 3546 6138 3564
rect 6120 3564 6138 3582
rect 6120 3582 6138 3600
rect 6120 3600 6138 3618
rect 6120 3618 6138 3636
rect 6120 3636 6138 3654
rect 6120 3654 6138 3672
rect 6120 3672 6138 3690
rect 6120 3690 6138 3708
rect 6120 3708 6138 3726
rect 6120 3726 6138 3744
rect 6120 3744 6138 3762
rect 6120 3762 6138 3780
rect 6120 3780 6138 3798
rect 6120 3798 6138 3816
rect 6120 3816 6138 3834
rect 6120 3834 6138 3852
rect 6120 3852 6138 3870
rect 6120 3870 6138 3888
rect 6120 3888 6138 3906
rect 6120 3906 6138 3924
rect 6120 3924 6138 3942
rect 6120 3942 6138 3960
rect 6120 3960 6138 3978
rect 6120 3978 6138 3996
rect 6120 3996 6138 4014
rect 6120 4014 6138 4032
rect 6120 4032 6138 4050
rect 6120 4050 6138 4068
rect 6120 4068 6138 4086
rect 6120 4086 6138 4104
rect 6120 4104 6138 4122
rect 6120 4122 6138 4140
rect 6120 4140 6138 4158
rect 6120 4158 6138 4176
rect 6120 4176 6138 4194
rect 6120 4194 6138 4212
rect 6120 4212 6138 4230
rect 6120 4230 6138 4248
rect 6120 4248 6138 4266
rect 6120 4266 6138 4284
rect 6120 4284 6138 4302
rect 6120 4302 6138 4320
rect 6120 4320 6138 4338
rect 6120 4338 6138 4356
rect 6120 4356 6138 4374
rect 6120 4374 6138 4392
rect 6120 4392 6138 4410
rect 6120 4410 6138 4428
rect 6120 4428 6138 4446
rect 6120 4446 6138 4464
rect 6120 4464 6138 4482
rect 6120 4482 6138 4500
rect 6120 4500 6138 4518
rect 6120 4518 6138 4536
rect 6120 4536 6138 4554
rect 6120 4554 6138 4572
rect 6120 4572 6138 4590
rect 6120 4590 6138 4608
rect 6120 4608 6138 4626
rect 6120 4626 6138 4644
rect 6120 4644 6138 4662
rect 6120 4662 6138 4680
rect 6120 4680 6138 4698
rect 6120 4698 6138 4716
rect 6120 4716 6138 4734
rect 6120 4734 6138 4752
rect 6120 4752 6138 4770
rect 6120 4770 6138 4788
rect 6120 4788 6138 4806
rect 6120 4806 6138 4824
rect 6120 4824 6138 4842
rect 6120 4842 6138 4860
rect 6120 4860 6138 4878
rect 6120 4878 6138 4896
rect 6120 4896 6138 4914
rect 6120 4914 6138 4932
rect 6120 4932 6138 4950
rect 6120 4950 6138 4968
rect 6120 4968 6138 4986
rect 6120 4986 6138 5004
rect 6120 5004 6138 5022
rect 6120 5022 6138 5040
rect 6120 5040 6138 5058
rect 6120 5058 6138 5076
rect 6120 5076 6138 5094
rect 6120 5094 6138 5112
rect 6120 5112 6138 5130
rect 6120 5130 6138 5148
rect 6120 5148 6138 5166
rect 6120 5166 6138 5184
rect 6120 5184 6138 5202
rect 6120 5202 6138 5220
rect 6120 5220 6138 5238
rect 6120 5238 6138 5256
rect 6120 5256 6138 5274
rect 6120 5274 6138 5292
rect 6120 5292 6138 5310
rect 6120 5310 6138 5328
rect 6120 5328 6138 5346
rect 6120 5346 6138 5364
rect 6120 5364 6138 5382
rect 6120 5382 6138 5400
rect 6120 5400 6138 5418
rect 6120 5418 6138 5436
rect 6120 5436 6138 5454
rect 6120 5454 6138 5472
rect 6120 5472 6138 5490
rect 6120 5760 6138 5778
rect 6120 5778 6138 5796
rect 6120 5796 6138 5814
rect 6120 5814 6138 5832
rect 6120 5832 6138 5850
rect 6120 5850 6138 5868
rect 6120 5868 6138 5886
rect 6120 5886 6138 5904
rect 6120 5904 6138 5922
rect 6120 5922 6138 5940
rect 6120 5940 6138 5958
rect 6120 5958 6138 5976
rect 6120 5976 6138 5994
rect 6120 5994 6138 6012
rect 6120 6012 6138 6030
rect 6120 6030 6138 6048
rect 6120 6048 6138 6066
rect 6120 6066 6138 6084
rect 6120 6084 6138 6102
rect 6120 6102 6138 6120
rect 6120 6120 6138 6138
rect 6120 6138 6138 6156
rect 6120 6156 6138 6174
rect 6120 6174 6138 6192
rect 6120 6192 6138 6210
rect 6120 6210 6138 6228
rect 6120 6228 6138 6246
rect 6120 6246 6138 6264
rect 6120 6264 6138 6282
rect 6120 6282 6138 6300
rect 6120 6300 6138 6318
rect 6120 6318 6138 6336
rect 6120 6336 6138 6354
rect 6120 6354 6138 6372
rect 6120 6372 6138 6390
rect 6120 6390 6138 6408
rect 6120 6408 6138 6426
rect 6120 6426 6138 6444
rect 6120 6444 6138 6462
rect 6120 6462 6138 6480
rect 6120 6480 6138 6498
rect 6120 6498 6138 6516
rect 6120 6516 6138 6534
rect 6120 6534 6138 6552
rect 6120 6552 6138 6570
rect 6120 6570 6138 6588
rect 6120 6588 6138 6606
rect 6120 6606 6138 6624
rect 6120 6624 6138 6642
rect 6120 6642 6138 6660
rect 6120 6660 6138 6678
rect 6120 6678 6138 6696
rect 6120 6696 6138 6714
rect 6120 6714 6138 6732
rect 6120 6732 6138 6750
rect 6120 6750 6138 6768
rect 6120 6768 6138 6786
rect 6120 6786 6138 6804
rect 6120 6804 6138 6822
rect 6120 6822 6138 6840
rect 6120 6840 6138 6858
rect 6120 6858 6138 6876
rect 6120 6876 6138 6894
rect 6120 6894 6138 6912
rect 6120 6912 6138 6930
rect 6120 6930 6138 6948
rect 6120 6948 6138 6966
rect 6120 6966 6138 6984
rect 6120 6984 6138 7002
rect 6120 7002 6138 7020
rect 6120 7020 6138 7038
rect 6120 7038 6138 7056
rect 6120 7056 6138 7074
rect 6120 7074 6138 7092
rect 6120 7092 6138 7110
rect 6120 7110 6138 7128
rect 6120 7128 6138 7146
rect 6120 7146 6138 7164
rect 6120 7164 6138 7182
rect 6120 7182 6138 7200
rect 6120 7200 6138 7218
rect 6120 7218 6138 7236
rect 6120 7236 6138 7254
rect 6120 7254 6138 7272
rect 6120 7272 6138 7290
rect 6120 7290 6138 7308
rect 6120 7308 6138 7326
rect 6120 7326 6138 7344
rect 6120 7344 6138 7362
rect 6120 7362 6138 7380
rect 6120 7380 6138 7398
rect 6120 7398 6138 7416
rect 6120 7416 6138 7434
rect 6120 7434 6138 7452
rect 6120 7452 6138 7470
rect 6120 7470 6138 7488
rect 6120 7488 6138 7506
rect 6120 7506 6138 7524
rect 6120 7524 6138 7542
rect 6120 7542 6138 7560
rect 6120 7560 6138 7578
rect 6120 7578 6138 7596
rect 6120 7596 6138 7614
rect 6120 7614 6138 7632
rect 6120 7632 6138 7650
rect 6120 7650 6138 7668
rect 6120 7668 6138 7686
rect 6120 7686 6138 7704
rect 6120 7704 6138 7722
rect 6120 7722 6138 7740
rect 6120 7740 6138 7758
rect 6120 7758 6138 7776
rect 6120 7776 6138 7794
rect 6120 7794 6138 7812
rect 6120 7812 6138 7830
rect 6120 7830 6138 7848
rect 6120 7848 6138 7866
rect 6120 7866 6138 7884
rect 6120 7884 6138 7902
rect 6120 7902 6138 7920
rect 6120 7920 6138 7938
rect 6120 7938 6138 7956
rect 6120 7956 6138 7974
rect 6120 7974 6138 7992
rect 6120 7992 6138 8010
rect 6120 8010 6138 8028
rect 6120 8028 6138 8046
rect 6120 8046 6138 8064
rect 6120 8064 6138 8082
rect 6120 8082 6138 8100
rect 6120 8100 6138 8118
rect 6120 8118 6138 8136
rect 6120 8136 6138 8154
rect 6120 8154 6138 8172
rect 6120 8172 6138 8190
rect 6120 8190 6138 8208
rect 6120 8208 6138 8226
rect 6120 8226 6138 8244
rect 6120 8244 6138 8262
rect 6120 8262 6138 8280
rect 6120 8280 6138 8298
rect 6120 8298 6138 8316
rect 6120 8316 6138 8334
rect 6120 8334 6138 8352
rect 6120 8352 6138 8370
rect 6120 8370 6138 8388
rect 6120 8388 6138 8406
rect 6120 8406 6138 8424
rect 6120 8424 6138 8442
rect 6120 8442 6138 8460
rect 6120 8460 6138 8478
rect 6120 8478 6138 8496
rect 6120 8496 6138 8514
rect 6120 8514 6138 8532
rect 6120 8532 6138 8550
rect 6120 8550 6138 8568
rect 6120 8568 6138 8586
rect 6120 8586 6138 8604
rect 6120 8604 6138 8622
rect 6120 8622 6138 8640
rect 6120 8640 6138 8658
rect 6120 8658 6138 8676
rect 6120 8676 6138 8694
rect 6120 8694 6138 8712
rect 6120 8712 6138 8730
rect 6120 8730 6138 8748
rect 6120 8748 6138 8766
rect 6120 8766 6138 8784
rect 6120 8784 6138 8802
rect 6120 8802 6138 8820
rect 6120 8820 6138 8838
rect 6120 8838 6138 8856
rect 6120 8856 6138 8874
rect 6120 8874 6138 8892
rect 6120 8892 6138 8910
rect 6120 8910 6138 8928
rect 6120 8928 6138 8946
rect 6120 8946 6138 8964
rect 6120 8964 6138 8982
rect 6120 8982 6138 9000
rect 6120 9000 6138 9018
rect 6120 9018 6138 9036
rect 6120 9036 6138 9054
rect 6120 9054 6138 9072
rect 6120 9072 6138 9090
rect 6120 9090 6138 9108
rect 6120 9108 6138 9126
rect 6120 9126 6138 9144
rect 6120 9144 6138 9162
rect 6120 9162 6138 9180
rect 6120 9180 6138 9198
rect 6120 9198 6138 9216
rect 6120 9216 6138 9234
rect 6120 9234 6138 9252
rect 6120 9252 6138 9270
rect 6120 9270 6138 9288
rect 6120 9288 6138 9306
rect 6120 9306 6138 9324
rect 6120 9324 6138 9342
rect 6120 9342 6138 9360
rect 6120 9360 6138 9378
rect 6138 1044 6156 1062
rect 6138 1062 6156 1080
rect 6138 1080 6156 1098
rect 6138 1098 6156 1116
rect 6138 1116 6156 1134
rect 6138 1134 6156 1152
rect 6138 1314 6156 1332
rect 6138 1332 6156 1350
rect 6138 1350 6156 1368
rect 6138 1368 6156 1386
rect 6138 1386 6156 1404
rect 6138 1404 6156 1422
rect 6138 1422 6156 1440
rect 6138 1440 6156 1458
rect 6138 1458 6156 1476
rect 6138 1476 6156 1494
rect 6138 1494 6156 1512
rect 6138 1512 6156 1530
rect 6138 1530 6156 1548
rect 6138 1548 6156 1566
rect 6138 1566 6156 1584
rect 6138 1584 6156 1602
rect 6138 1602 6156 1620
rect 6138 1620 6156 1638
rect 6138 1638 6156 1656
rect 6138 1656 6156 1674
rect 6138 1674 6156 1692
rect 6138 1692 6156 1710
rect 6138 1710 6156 1728
rect 6138 1728 6156 1746
rect 6138 1746 6156 1764
rect 6138 1764 6156 1782
rect 6138 1782 6156 1800
rect 6138 1800 6156 1818
rect 6138 1818 6156 1836
rect 6138 1836 6156 1854
rect 6138 1854 6156 1872
rect 6138 1872 6156 1890
rect 6138 1890 6156 1908
rect 6138 1908 6156 1926
rect 6138 1926 6156 1944
rect 6138 1944 6156 1962
rect 6138 1962 6156 1980
rect 6138 1980 6156 1998
rect 6138 1998 6156 2016
rect 6138 2016 6156 2034
rect 6138 2034 6156 2052
rect 6138 2052 6156 2070
rect 6138 2070 6156 2088
rect 6138 2088 6156 2106
rect 6138 2106 6156 2124
rect 6138 2124 6156 2142
rect 6138 2142 6156 2160
rect 6138 2160 6156 2178
rect 6138 2178 6156 2196
rect 6138 2196 6156 2214
rect 6138 2214 6156 2232
rect 6138 2232 6156 2250
rect 6138 2250 6156 2268
rect 6138 2268 6156 2286
rect 6138 2286 6156 2304
rect 6138 2304 6156 2322
rect 6138 2322 6156 2340
rect 6138 2340 6156 2358
rect 6138 2358 6156 2376
rect 6138 2376 6156 2394
rect 6138 2394 6156 2412
rect 6138 2412 6156 2430
rect 6138 2430 6156 2448
rect 6138 2448 6156 2466
rect 6138 2466 6156 2484
rect 6138 2484 6156 2502
rect 6138 2502 6156 2520
rect 6138 2520 6156 2538
rect 6138 2538 6156 2556
rect 6138 2556 6156 2574
rect 6138 2574 6156 2592
rect 6138 2592 6156 2610
rect 6138 2610 6156 2628
rect 6138 2628 6156 2646
rect 6138 2646 6156 2664
rect 6138 2664 6156 2682
rect 6138 2682 6156 2700
rect 6138 2700 6156 2718
rect 6138 2718 6156 2736
rect 6138 2736 6156 2754
rect 6138 2754 6156 2772
rect 6138 2772 6156 2790
rect 6138 2790 6156 2808
rect 6138 3060 6156 3078
rect 6138 3078 6156 3096
rect 6138 3096 6156 3114
rect 6138 3114 6156 3132
rect 6138 3132 6156 3150
rect 6138 3150 6156 3168
rect 6138 3168 6156 3186
rect 6138 3186 6156 3204
rect 6138 3204 6156 3222
rect 6138 3222 6156 3240
rect 6138 3240 6156 3258
rect 6138 3258 6156 3276
rect 6138 3276 6156 3294
rect 6138 3294 6156 3312
rect 6138 3312 6156 3330
rect 6138 3330 6156 3348
rect 6138 3348 6156 3366
rect 6138 3366 6156 3384
rect 6138 3384 6156 3402
rect 6138 3402 6156 3420
rect 6138 3420 6156 3438
rect 6138 3438 6156 3456
rect 6138 3456 6156 3474
rect 6138 3474 6156 3492
rect 6138 3492 6156 3510
rect 6138 3510 6156 3528
rect 6138 3528 6156 3546
rect 6138 3546 6156 3564
rect 6138 3564 6156 3582
rect 6138 3582 6156 3600
rect 6138 3600 6156 3618
rect 6138 3618 6156 3636
rect 6138 3636 6156 3654
rect 6138 3654 6156 3672
rect 6138 3672 6156 3690
rect 6138 3690 6156 3708
rect 6138 3708 6156 3726
rect 6138 3726 6156 3744
rect 6138 3744 6156 3762
rect 6138 3762 6156 3780
rect 6138 3780 6156 3798
rect 6138 3798 6156 3816
rect 6138 3816 6156 3834
rect 6138 3834 6156 3852
rect 6138 3852 6156 3870
rect 6138 3870 6156 3888
rect 6138 3888 6156 3906
rect 6138 3906 6156 3924
rect 6138 3924 6156 3942
rect 6138 3942 6156 3960
rect 6138 3960 6156 3978
rect 6138 3978 6156 3996
rect 6138 3996 6156 4014
rect 6138 4014 6156 4032
rect 6138 4032 6156 4050
rect 6138 4050 6156 4068
rect 6138 4068 6156 4086
rect 6138 4086 6156 4104
rect 6138 4104 6156 4122
rect 6138 4122 6156 4140
rect 6138 4140 6156 4158
rect 6138 4158 6156 4176
rect 6138 4176 6156 4194
rect 6138 4194 6156 4212
rect 6138 4212 6156 4230
rect 6138 4230 6156 4248
rect 6138 4248 6156 4266
rect 6138 4266 6156 4284
rect 6138 4284 6156 4302
rect 6138 4302 6156 4320
rect 6138 4320 6156 4338
rect 6138 4338 6156 4356
rect 6138 4356 6156 4374
rect 6138 4374 6156 4392
rect 6138 4392 6156 4410
rect 6138 4410 6156 4428
rect 6138 4428 6156 4446
rect 6138 4446 6156 4464
rect 6138 4464 6156 4482
rect 6138 4482 6156 4500
rect 6138 4500 6156 4518
rect 6138 4518 6156 4536
rect 6138 4536 6156 4554
rect 6138 4554 6156 4572
rect 6138 4572 6156 4590
rect 6138 4590 6156 4608
rect 6138 4608 6156 4626
rect 6138 4626 6156 4644
rect 6138 4644 6156 4662
rect 6138 4662 6156 4680
rect 6138 4680 6156 4698
rect 6138 4698 6156 4716
rect 6138 4716 6156 4734
rect 6138 4734 6156 4752
rect 6138 4752 6156 4770
rect 6138 4770 6156 4788
rect 6138 4788 6156 4806
rect 6138 4806 6156 4824
rect 6138 4824 6156 4842
rect 6138 4842 6156 4860
rect 6138 4860 6156 4878
rect 6138 4878 6156 4896
rect 6138 4896 6156 4914
rect 6138 4914 6156 4932
rect 6138 4932 6156 4950
rect 6138 4950 6156 4968
rect 6138 4968 6156 4986
rect 6138 4986 6156 5004
rect 6138 5004 6156 5022
rect 6138 5022 6156 5040
rect 6138 5040 6156 5058
rect 6138 5058 6156 5076
rect 6138 5076 6156 5094
rect 6138 5094 6156 5112
rect 6138 5112 6156 5130
rect 6138 5130 6156 5148
rect 6138 5148 6156 5166
rect 6138 5166 6156 5184
rect 6138 5184 6156 5202
rect 6138 5202 6156 5220
rect 6138 5220 6156 5238
rect 6138 5238 6156 5256
rect 6138 5256 6156 5274
rect 6138 5274 6156 5292
rect 6138 5292 6156 5310
rect 6138 5310 6156 5328
rect 6138 5328 6156 5346
rect 6138 5346 6156 5364
rect 6138 5364 6156 5382
rect 6138 5382 6156 5400
rect 6138 5400 6156 5418
rect 6138 5418 6156 5436
rect 6138 5436 6156 5454
rect 6138 5454 6156 5472
rect 6138 5472 6156 5490
rect 6138 5490 6156 5508
rect 6138 5778 6156 5796
rect 6138 5796 6156 5814
rect 6138 5814 6156 5832
rect 6138 5832 6156 5850
rect 6138 5850 6156 5868
rect 6138 5868 6156 5886
rect 6138 5886 6156 5904
rect 6138 5904 6156 5922
rect 6138 5922 6156 5940
rect 6138 5940 6156 5958
rect 6138 5958 6156 5976
rect 6138 5976 6156 5994
rect 6138 5994 6156 6012
rect 6138 6012 6156 6030
rect 6138 6030 6156 6048
rect 6138 6048 6156 6066
rect 6138 6066 6156 6084
rect 6138 6084 6156 6102
rect 6138 6102 6156 6120
rect 6138 6120 6156 6138
rect 6138 6138 6156 6156
rect 6138 6156 6156 6174
rect 6138 6174 6156 6192
rect 6138 6192 6156 6210
rect 6138 6210 6156 6228
rect 6138 6228 6156 6246
rect 6138 6246 6156 6264
rect 6138 6264 6156 6282
rect 6138 6282 6156 6300
rect 6138 6300 6156 6318
rect 6138 6318 6156 6336
rect 6138 6336 6156 6354
rect 6138 6354 6156 6372
rect 6138 6372 6156 6390
rect 6138 6390 6156 6408
rect 6138 6408 6156 6426
rect 6138 6426 6156 6444
rect 6138 6444 6156 6462
rect 6138 6462 6156 6480
rect 6138 6480 6156 6498
rect 6138 6498 6156 6516
rect 6138 6516 6156 6534
rect 6138 6534 6156 6552
rect 6138 6552 6156 6570
rect 6138 6570 6156 6588
rect 6138 6588 6156 6606
rect 6138 6606 6156 6624
rect 6138 6624 6156 6642
rect 6138 6642 6156 6660
rect 6138 6660 6156 6678
rect 6138 6678 6156 6696
rect 6138 6696 6156 6714
rect 6138 6714 6156 6732
rect 6138 6732 6156 6750
rect 6138 6750 6156 6768
rect 6138 6768 6156 6786
rect 6138 6786 6156 6804
rect 6138 6804 6156 6822
rect 6138 6822 6156 6840
rect 6138 6840 6156 6858
rect 6138 6858 6156 6876
rect 6138 6876 6156 6894
rect 6138 6894 6156 6912
rect 6138 6912 6156 6930
rect 6138 6930 6156 6948
rect 6138 6948 6156 6966
rect 6138 6966 6156 6984
rect 6138 6984 6156 7002
rect 6138 7002 6156 7020
rect 6138 7020 6156 7038
rect 6138 7038 6156 7056
rect 6138 7056 6156 7074
rect 6138 7074 6156 7092
rect 6138 7092 6156 7110
rect 6138 7110 6156 7128
rect 6138 7128 6156 7146
rect 6138 7146 6156 7164
rect 6138 7164 6156 7182
rect 6138 7182 6156 7200
rect 6138 7200 6156 7218
rect 6138 7218 6156 7236
rect 6138 7236 6156 7254
rect 6138 7254 6156 7272
rect 6138 7272 6156 7290
rect 6138 7290 6156 7308
rect 6138 7308 6156 7326
rect 6138 7326 6156 7344
rect 6138 7344 6156 7362
rect 6138 7362 6156 7380
rect 6138 7380 6156 7398
rect 6138 7398 6156 7416
rect 6138 7416 6156 7434
rect 6138 7434 6156 7452
rect 6138 7452 6156 7470
rect 6138 7470 6156 7488
rect 6138 7488 6156 7506
rect 6138 7506 6156 7524
rect 6138 7524 6156 7542
rect 6138 7542 6156 7560
rect 6138 7560 6156 7578
rect 6138 7578 6156 7596
rect 6138 7596 6156 7614
rect 6138 7614 6156 7632
rect 6138 7632 6156 7650
rect 6138 7650 6156 7668
rect 6138 7668 6156 7686
rect 6138 7686 6156 7704
rect 6138 7704 6156 7722
rect 6138 7722 6156 7740
rect 6138 7740 6156 7758
rect 6138 7758 6156 7776
rect 6138 7776 6156 7794
rect 6138 7794 6156 7812
rect 6138 7812 6156 7830
rect 6138 7830 6156 7848
rect 6138 7848 6156 7866
rect 6138 7866 6156 7884
rect 6138 7884 6156 7902
rect 6138 7902 6156 7920
rect 6138 7920 6156 7938
rect 6138 7938 6156 7956
rect 6138 7956 6156 7974
rect 6138 7974 6156 7992
rect 6138 7992 6156 8010
rect 6138 8010 6156 8028
rect 6138 8028 6156 8046
rect 6138 8046 6156 8064
rect 6138 8064 6156 8082
rect 6138 8082 6156 8100
rect 6138 8100 6156 8118
rect 6138 8118 6156 8136
rect 6138 8136 6156 8154
rect 6138 8154 6156 8172
rect 6138 8172 6156 8190
rect 6138 8190 6156 8208
rect 6138 8208 6156 8226
rect 6138 8226 6156 8244
rect 6138 8244 6156 8262
rect 6138 8262 6156 8280
rect 6138 8280 6156 8298
rect 6138 8298 6156 8316
rect 6138 8316 6156 8334
rect 6138 8334 6156 8352
rect 6138 8352 6156 8370
rect 6138 8370 6156 8388
rect 6138 8388 6156 8406
rect 6138 8406 6156 8424
rect 6138 8424 6156 8442
rect 6138 8442 6156 8460
rect 6138 8460 6156 8478
rect 6138 8478 6156 8496
rect 6138 8496 6156 8514
rect 6138 8514 6156 8532
rect 6138 8532 6156 8550
rect 6138 8550 6156 8568
rect 6138 8568 6156 8586
rect 6138 8586 6156 8604
rect 6138 8604 6156 8622
rect 6138 8622 6156 8640
rect 6138 8640 6156 8658
rect 6138 8658 6156 8676
rect 6138 8676 6156 8694
rect 6138 8694 6156 8712
rect 6138 8712 6156 8730
rect 6138 8730 6156 8748
rect 6138 8748 6156 8766
rect 6138 8766 6156 8784
rect 6138 8784 6156 8802
rect 6138 8802 6156 8820
rect 6138 8820 6156 8838
rect 6138 8838 6156 8856
rect 6138 8856 6156 8874
rect 6138 8874 6156 8892
rect 6138 8892 6156 8910
rect 6138 8910 6156 8928
rect 6138 8928 6156 8946
rect 6138 8946 6156 8964
rect 6138 8964 6156 8982
rect 6138 8982 6156 9000
rect 6138 9000 6156 9018
rect 6138 9018 6156 9036
rect 6138 9036 6156 9054
rect 6138 9054 6156 9072
rect 6138 9072 6156 9090
rect 6138 9090 6156 9108
rect 6138 9108 6156 9126
rect 6138 9126 6156 9144
rect 6138 9144 6156 9162
rect 6138 9162 6156 9180
rect 6138 9180 6156 9198
rect 6138 9198 6156 9216
rect 6138 9216 6156 9234
rect 6138 9234 6156 9252
rect 6138 9252 6156 9270
rect 6138 9270 6156 9288
rect 6138 9288 6156 9306
rect 6138 9306 6156 9324
rect 6138 9324 6156 9342
rect 6138 9342 6156 9360
rect 6138 9360 6156 9378
rect 6138 9378 6156 9396
rect 6138 9396 6156 9414
rect 6156 1062 6174 1080
rect 6156 1080 6174 1098
rect 6156 1098 6174 1116
rect 6156 1116 6174 1134
rect 6156 1134 6174 1152
rect 6156 1152 6174 1170
rect 6156 1314 6174 1332
rect 6156 1332 6174 1350
rect 6156 1350 6174 1368
rect 6156 1368 6174 1386
rect 6156 1386 6174 1404
rect 6156 1404 6174 1422
rect 6156 1422 6174 1440
rect 6156 1440 6174 1458
rect 6156 1458 6174 1476
rect 6156 1476 6174 1494
rect 6156 1494 6174 1512
rect 6156 1512 6174 1530
rect 6156 1530 6174 1548
rect 6156 1548 6174 1566
rect 6156 1566 6174 1584
rect 6156 1584 6174 1602
rect 6156 1602 6174 1620
rect 6156 1620 6174 1638
rect 6156 1638 6174 1656
rect 6156 1656 6174 1674
rect 6156 1674 6174 1692
rect 6156 1692 6174 1710
rect 6156 1710 6174 1728
rect 6156 1728 6174 1746
rect 6156 1746 6174 1764
rect 6156 1764 6174 1782
rect 6156 1782 6174 1800
rect 6156 1800 6174 1818
rect 6156 1818 6174 1836
rect 6156 1836 6174 1854
rect 6156 1854 6174 1872
rect 6156 1872 6174 1890
rect 6156 1890 6174 1908
rect 6156 1908 6174 1926
rect 6156 1926 6174 1944
rect 6156 1944 6174 1962
rect 6156 1962 6174 1980
rect 6156 1980 6174 1998
rect 6156 1998 6174 2016
rect 6156 2016 6174 2034
rect 6156 2034 6174 2052
rect 6156 2052 6174 2070
rect 6156 2070 6174 2088
rect 6156 2088 6174 2106
rect 6156 2106 6174 2124
rect 6156 2124 6174 2142
rect 6156 2142 6174 2160
rect 6156 2160 6174 2178
rect 6156 2178 6174 2196
rect 6156 2196 6174 2214
rect 6156 2214 6174 2232
rect 6156 2232 6174 2250
rect 6156 2250 6174 2268
rect 6156 2268 6174 2286
rect 6156 2286 6174 2304
rect 6156 2304 6174 2322
rect 6156 2322 6174 2340
rect 6156 2340 6174 2358
rect 6156 2358 6174 2376
rect 6156 2376 6174 2394
rect 6156 2394 6174 2412
rect 6156 2412 6174 2430
rect 6156 2430 6174 2448
rect 6156 2448 6174 2466
rect 6156 2466 6174 2484
rect 6156 2484 6174 2502
rect 6156 2502 6174 2520
rect 6156 2520 6174 2538
rect 6156 2538 6174 2556
rect 6156 2556 6174 2574
rect 6156 2574 6174 2592
rect 6156 2592 6174 2610
rect 6156 2610 6174 2628
rect 6156 2628 6174 2646
rect 6156 2646 6174 2664
rect 6156 2664 6174 2682
rect 6156 2682 6174 2700
rect 6156 2700 6174 2718
rect 6156 2718 6174 2736
rect 6156 2736 6174 2754
rect 6156 2754 6174 2772
rect 6156 2772 6174 2790
rect 6156 2790 6174 2808
rect 6156 3060 6174 3078
rect 6156 3078 6174 3096
rect 6156 3096 6174 3114
rect 6156 3114 6174 3132
rect 6156 3132 6174 3150
rect 6156 3150 6174 3168
rect 6156 3168 6174 3186
rect 6156 3186 6174 3204
rect 6156 3204 6174 3222
rect 6156 3222 6174 3240
rect 6156 3240 6174 3258
rect 6156 3258 6174 3276
rect 6156 3276 6174 3294
rect 6156 3294 6174 3312
rect 6156 3312 6174 3330
rect 6156 3330 6174 3348
rect 6156 3348 6174 3366
rect 6156 3366 6174 3384
rect 6156 3384 6174 3402
rect 6156 3402 6174 3420
rect 6156 3420 6174 3438
rect 6156 3438 6174 3456
rect 6156 3456 6174 3474
rect 6156 3474 6174 3492
rect 6156 3492 6174 3510
rect 6156 3510 6174 3528
rect 6156 3528 6174 3546
rect 6156 3546 6174 3564
rect 6156 3564 6174 3582
rect 6156 3582 6174 3600
rect 6156 3600 6174 3618
rect 6156 3618 6174 3636
rect 6156 3636 6174 3654
rect 6156 3654 6174 3672
rect 6156 3672 6174 3690
rect 6156 3690 6174 3708
rect 6156 3708 6174 3726
rect 6156 3726 6174 3744
rect 6156 3744 6174 3762
rect 6156 3762 6174 3780
rect 6156 3780 6174 3798
rect 6156 3798 6174 3816
rect 6156 3816 6174 3834
rect 6156 3834 6174 3852
rect 6156 3852 6174 3870
rect 6156 3870 6174 3888
rect 6156 3888 6174 3906
rect 6156 3906 6174 3924
rect 6156 3924 6174 3942
rect 6156 3942 6174 3960
rect 6156 3960 6174 3978
rect 6156 3978 6174 3996
rect 6156 3996 6174 4014
rect 6156 4014 6174 4032
rect 6156 4032 6174 4050
rect 6156 4050 6174 4068
rect 6156 4068 6174 4086
rect 6156 4086 6174 4104
rect 6156 4104 6174 4122
rect 6156 4122 6174 4140
rect 6156 4140 6174 4158
rect 6156 4158 6174 4176
rect 6156 4176 6174 4194
rect 6156 4194 6174 4212
rect 6156 4212 6174 4230
rect 6156 4230 6174 4248
rect 6156 4248 6174 4266
rect 6156 4266 6174 4284
rect 6156 4284 6174 4302
rect 6156 4302 6174 4320
rect 6156 4320 6174 4338
rect 6156 4338 6174 4356
rect 6156 4356 6174 4374
rect 6156 4374 6174 4392
rect 6156 4392 6174 4410
rect 6156 4410 6174 4428
rect 6156 4428 6174 4446
rect 6156 4446 6174 4464
rect 6156 4464 6174 4482
rect 6156 4482 6174 4500
rect 6156 4500 6174 4518
rect 6156 4518 6174 4536
rect 6156 4536 6174 4554
rect 6156 4554 6174 4572
rect 6156 4572 6174 4590
rect 6156 4590 6174 4608
rect 6156 4608 6174 4626
rect 6156 4626 6174 4644
rect 6156 4644 6174 4662
rect 6156 4662 6174 4680
rect 6156 4680 6174 4698
rect 6156 4698 6174 4716
rect 6156 4716 6174 4734
rect 6156 4734 6174 4752
rect 6156 4752 6174 4770
rect 6156 4770 6174 4788
rect 6156 4788 6174 4806
rect 6156 4806 6174 4824
rect 6156 4824 6174 4842
rect 6156 4842 6174 4860
rect 6156 4860 6174 4878
rect 6156 4878 6174 4896
rect 6156 4896 6174 4914
rect 6156 4914 6174 4932
rect 6156 4932 6174 4950
rect 6156 4950 6174 4968
rect 6156 4968 6174 4986
rect 6156 4986 6174 5004
rect 6156 5004 6174 5022
rect 6156 5022 6174 5040
rect 6156 5040 6174 5058
rect 6156 5058 6174 5076
rect 6156 5076 6174 5094
rect 6156 5094 6174 5112
rect 6156 5112 6174 5130
rect 6156 5130 6174 5148
rect 6156 5148 6174 5166
rect 6156 5166 6174 5184
rect 6156 5184 6174 5202
rect 6156 5202 6174 5220
rect 6156 5220 6174 5238
rect 6156 5238 6174 5256
rect 6156 5256 6174 5274
rect 6156 5274 6174 5292
rect 6156 5292 6174 5310
rect 6156 5310 6174 5328
rect 6156 5328 6174 5346
rect 6156 5346 6174 5364
rect 6156 5364 6174 5382
rect 6156 5382 6174 5400
rect 6156 5400 6174 5418
rect 6156 5418 6174 5436
rect 6156 5436 6174 5454
rect 6156 5454 6174 5472
rect 6156 5472 6174 5490
rect 6156 5490 6174 5508
rect 6156 5508 6174 5526
rect 6156 5796 6174 5814
rect 6156 5814 6174 5832
rect 6156 5832 6174 5850
rect 6156 5850 6174 5868
rect 6156 5868 6174 5886
rect 6156 5886 6174 5904
rect 6156 5904 6174 5922
rect 6156 5922 6174 5940
rect 6156 5940 6174 5958
rect 6156 5958 6174 5976
rect 6156 5976 6174 5994
rect 6156 5994 6174 6012
rect 6156 6012 6174 6030
rect 6156 6030 6174 6048
rect 6156 6048 6174 6066
rect 6156 6066 6174 6084
rect 6156 6084 6174 6102
rect 6156 6102 6174 6120
rect 6156 6120 6174 6138
rect 6156 6138 6174 6156
rect 6156 6156 6174 6174
rect 6156 6174 6174 6192
rect 6156 6192 6174 6210
rect 6156 6210 6174 6228
rect 6156 6228 6174 6246
rect 6156 6246 6174 6264
rect 6156 6264 6174 6282
rect 6156 6282 6174 6300
rect 6156 6300 6174 6318
rect 6156 6318 6174 6336
rect 6156 6336 6174 6354
rect 6156 6354 6174 6372
rect 6156 6372 6174 6390
rect 6156 6390 6174 6408
rect 6156 6408 6174 6426
rect 6156 6426 6174 6444
rect 6156 6444 6174 6462
rect 6156 6462 6174 6480
rect 6156 6480 6174 6498
rect 6156 6498 6174 6516
rect 6156 6516 6174 6534
rect 6156 6534 6174 6552
rect 6156 6552 6174 6570
rect 6156 6570 6174 6588
rect 6156 6588 6174 6606
rect 6156 6606 6174 6624
rect 6156 6624 6174 6642
rect 6156 6642 6174 6660
rect 6156 6660 6174 6678
rect 6156 6678 6174 6696
rect 6156 6696 6174 6714
rect 6156 6714 6174 6732
rect 6156 6732 6174 6750
rect 6156 6750 6174 6768
rect 6156 6768 6174 6786
rect 6156 6786 6174 6804
rect 6156 6804 6174 6822
rect 6156 6822 6174 6840
rect 6156 6840 6174 6858
rect 6156 6858 6174 6876
rect 6156 6876 6174 6894
rect 6156 6894 6174 6912
rect 6156 6912 6174 6930
rect 6156 6930 6174 6948
rect 6156 6948 6174 6966
rect 6156 6966 6174 6984
rect 6156 6984 6174 7002
rect 6156 7002 6174 7020
rect 6156 7020 6174 7038
rect 6156 7038 6174 7056
rect 6156 7056 6174 7074
rect 6156 7074 6174 7092
rect 6156 7092 6174 7110
rect 6156 7110 6174 7128
rect 6156 7128 6174 7146
rect 6156 7146 6174 7164
rect 6156 7164 6174 7182
rect 6156 7182 6174 7200
rect 6156 7200 6174 7218
rect 6156 7218 6174 7236
rect 6156 7236 6174 7254
rect 6156 7254 6174 7272
rect 6156 7272 6174 7290
rect 6156 7290 6174 7308
rect 6156 7308 6174 7326
rect 6156 7326 6174 7344
rect 6156 7344 6174 7362
rect 6156 7362 6174 7380
rect 6156 7380 6174 7398
rect 6156 7398 6174 7416
rect 6156 7416 6174 7434
rect 6156 7434 6174 7452
rect 6156 7452 6174 7470
rect 6156 7470 6174 7488
rect 6156 7488 6174 7506
rect 6156 7506 6174 7524
rect 6156 7524 6174 7542
rect 6156 7542 6174 7560
rect 6156 7560 6174 7578
rect 6156 7578 6174 7596
rect 6156 7596 6174 7614
rect 6156 7614 6174 7632
rect 6156 7632 6174 7650
rect 6156 7650 6174 7668
rect 6156 7668 6174 7686
rect 6156 7686 6174 7704
rect 6156 7704 6174 7722
rect 6156 7722 6174 7740
rect 6156 7740 6174 7758
rect 6156 7758 6174 7776
rect 6156 7776 6174 7794
rect 6156 7794 6174 7812
rect 6156 7812 6174 7830
rect 6156 7830 6174 7848
rect 6156 7848 6174 7866
rect 6156 7866 6174 7884
rect 6156 7884 6174 7902
rect 6156 7902 6174 7920
rect 6156 7920 6174 7938
rect 6156 7938 6174 7956
rect 6156 7956 6174 7974
rect 6156 7974 6174 7992
rect 6156 7992 6174 8010
rect 6156 8010 6174 8028
rect 6156 8028 6174 8046
rect 6156 8046 6174 8064
rect 6156 8064 6174 8082
rect 6156 8082 6174 8100
rect 6156 8100 6174 8118
rect 6156 8118 6174 8136
rect 6156 8136 6174 8154
rect 6156 8154 6174 8172
rect 6156 8172 6174 8190
rect 6156 8190 6174 8208
rect 6156 8208 6174 8226
rect 6156 8226 6174 8244
rect 6156 8244 6174 8262
rect 6156 8262 6174 8280
rect 6156 8280 6174 8298
rect 6156 8298 6174 8316
rect 6156 8316 6174 8334
rect 6156 8334 6174 8352
rect 6156 8352 6174 8370
rect 6156 8370 6174 8388
rect 6156 8388 6174 8406
rect 6156 8406 6174 8424
rect 6156 8424 6174 8442
rect 6156 8442 6174 8460
rect 6156 8460 6174 8478
rect 6156 8478 6174 8496
rect 6156 8496 6174 8514
rect 6156 8514 6174 8532
rect 6156 8532 6174 8550
rect 6156 8550 6174 8568
rect 6156 8568 6174 8586
rect 6156 8586 6174 8604
rect 6156 8604 6174 8622
rect 6156 8622 6174 8640
rect 6156 8640 6174 8658
rect 6156 8658 6174 8676
rect 6156 8676 6174 8694
rect 6156 8694 6174 8712
rect 6156 8712 6174 8730
rect 6156 8730 6174 8748
rect 6156 8748 6174 8766
rect 6156 8766 6174 8784
rect 6156 8784 6174 8802
rect 6156 8802 6174 8820
rect 6156 8820 6174 8838
rect 6156 8838 6174 8856
rect 6156 8856 6174 8874
rect 6156 8874 6174 8892
rect 6156 8892 6174 8910
rect 6156 8910 6174 8928
rect 6156 8928 6174 8946
rect 6156 8946 6174 8964
rect 6156 8964 6174 8982
rect 6156 8982 6174 9000
rect 6156 9000 6174 9018
rect 6156 9018 6174 9036
rect 6156 9036 6174 9054
rect 6156 9054 6174 9072
rect 6156 9072 6174 9090
rect 6156 9090 6174 9108
rect 6156 9108 6174 9126
rect 6156 9126 6174 9144
rect 6156 9144 6174 9162
rect 6156 9162 6174 9180
rect 6156 9180 6174 9198
rect 6156 9198 6174 9216
rect 6156 9216 6174 9234
rect 6156 9234 6174 9252
rect 6156 9252 6174 9270
rect 6156 9270 6174 9288
rect 6156 9288 6174 9306
rect 6156 9306 6174 9324
rect 6156 9324 6174 9342
rect 6156 9342 6174 9360
rect 6156 9360 6174 9378
rect 6156 9378 6174 9396
rect 6156 9396 6174 9414
rect 6156 9414 6174 9432
rect 6174 1062 6192 1080
rect 6174 1080 6192 1098
rect 6174 1098 6192 1116
rect 6174 1116 6192 1134
rect 6174 1134 6192 1152
rect 6174 1152 6192 1170
rect 6174 1314 6192 1332
rect 6174 1332 6192 1350
rect 6174 1350 6192 1368
rect 6174 1368 6192 1386
rect 6174 1386 6192 1404
rect 6174 1404 6192 1422
rect 6174 1422 6192 1440
rect 6174 1440 6192 1458
rect 6174 1458 6192 1476
rect 6174 1476 6192 1494
rect 6174 1494 6192 1512
rect 6174 1512 6192 1530
rect 6174 1530 6192 1548
rect 6174 1548 6192 1566
rect 6174 1566 6192 1584
rect 6174 1584 6192 1602
rect 6174 1602 6192 1620
rect 6174 1620 6192 1638
rect 6174 1638 6192 1656
rect 6174 1656 6192 1674
rect 6174 1674 6192 1692
rect 6174 1692 6192 1710
rect 6174 1710 6192 1728
rect 6174 1728 6192 1746
rect 6174 1746 6192 1764
rect 6174 1764 6192 1782
rect 6174 1782 6192 1800
rect 6174 1800 6192 1818
rect 6174 1818 6192 1836
rect 6174 1836 6192 1854
rect 6174 1854 6192 1872
rect 6174 1872 6192 1890
rect 6174 1890 6192 1908
rect 6174 1908 6192 1926
rect 6174 1926 6192 1944
rect 6174 1944 6192 1962
rect 6174 1962 6192 1980
rect 6174 1980 6192 1998
rect 6174 1998 6192 2016
rect 6174 2016 6192 2034
rect 6174 2034 6192 2052
rect 6174 2052 6192 2070
rect 6174 2070 6192 2088
rect 6174 2088 6192 2106
rect 6174 2106 6192 2124
rect 6174 2124 6192 2142
rect 6174 2142 6192 2160
rect 6174 2160 6192 2178
rect 6174 2178 6192 2196
rect 6174 2196 6192 2214
rect 6174 2214 6192 2232
rect 6174 2232 6192 2250
rect 6174 2250 6192 2268
rect 6174 2268 6192 2286
rect 6174 2286 6192 2304
rect 6174 2304 6192 2322
rect 6174 2322 6192 2340
rect 6174 2340 6192 2358
rect 6174 2358 6192 2376
rect 6174 2376 6192 2394
rect 6174 2394 6192 2412
rect 6174 2412 6192 2430
rect 6174 2430 6192 2448
rect 6174 2448 6192 2466
rect 6174 2466 6192 2484
rect 6174 2484 6192 2502
rect 6174 2502 6192 2520
rect 6174 2520 6192 2538
rect 6174 2538 6192 2556
rect 6174 2556 6192 2574
rect 6174 2574 6192 2592
rect 6174 2592 6192 2610
rect 6174 2610 6192 2628
rect 6174 2628 6192 2646
rect 6174 2646 6192 2664
rect 6174 2664 6192 2682
rect 6174 2682 6192 2700
rect 6174 2700 6192 2718
rect 6174 2718 6192 2736
rect 6174 2736 6192 2754
rect 6174 2754 6192 2772
rect 6174 2772 6192 2790
rect 6174 2790 6192 2808
rect 6174 2808 6192 2826
rect 6174 3078 6192 3096
rect 6174 3096 6192 3114
rect 6174 3114 6192 3132
rect 6174 3132 6192 3150
rect 6174 3150 6192 3168
rect 6174 3168 6192 3186
rect 6174 3186 6192 3204
rect 6174 3204 6192 3222
rect 6174 3222 6192 3240
rect 6174 3240 6192 3258
rect 6174 3258 6192 3276
rect 6174 3276 6192 3294
rect 6174 3294 6192 3312
rect 6174 3312 6192 3330
rect 6174 3330 6192 3348
rect 6174 3348 6192 3366
rect 6174 3366 6192 3384
rect 6174 3384 6192 3402
rect 6174 3402 6192 3420
rect 6174 3420 6192 3438
rect 6174 3438 6192 3456
rect 6174 3456 6192 3474
rect 6174 3474 6192 3492
rect 6174 3492 6192 3510
rect 6174 3510 6192 3528
rect 6174 3528 6192 3546
rect 6174 3546 6192 3564
rect 6174 3564 6192 3582
rect 6174 3582 6192 3600
rect 6174 3600 6192 3618
rect 6174 3618 6192 3636
rect 6174 3636 6192 3654
rect 6174 3654 6192 3672
rect 6174 3672 6192 3690
rect 6174 3690 6192 3708
rect 6174 3708 6192 3726
rect 6174 3726 6192 3744
rect 6174 3744 6192 3762
rect 6174 3762 6192 3780
rect 6174 3780 6192 3798
rect 6174 3798 6192 3816
rect 6174 3816 6192 3834
rect 6174 3834 6192 3852
rect 6174 3852 6192 3870
rect 6174 3870 6192 3888
rect 6174 3888 6192 3906
rect 6174 3906 6192 3924
rect 6174 3924 6192 3942
rect 6174 3942 6192 3960
rect 6174 3960 6192 3978
rect 6174 3978 6192 3996
rect 6174 3996 6192 4014
rect 6174 4014 6192 4032
rect 6174 4032 6192 4050
rect 6174 4050 6192 4068
rect 6174 4068 6192 4086
rect 6174 4086 6192 4104
rect 6174 4104 6192 4122
rect 6174 4122 6192 4140
rect 6174 4140 6192 4158
rect 6174 4158 6192 4176
rect 6174 4176 6192 4194
rect 6174 4194 6192 4212
rect 6174 4212 6192 4230
rect 6174 4230 6192 4248
rect 6174 4248 6192 4266
rect 6174 4266 6192 4284
rect 6174 4284 6192 4302
rect 6174 4302 6192 4320
rect 6174 4320 6192 4338
rect 6174 4338 6192 4356
rect 6174 4356 6192 4374
rect 6174 4374 6192 4392
rect 6174 4392 6192 4410
rect 6174 4410 6192 4428
rect 6174 4428 6192 4446
rect 6174 4446 6192 4464
rect 6174 4464 6192 4482
rect 6174 4482 6192 4500
rect 6174 4500 6192 4518
rect 6174 4518 6192 4536
rect 6174 4536 6192 4554
rect 6174 4554 6192 4572
rect 6174 4572 6192 4590
rect 6174 4590 6192 4608
rect 6174 4608 6192 4626
rect 6174 4626 6192 4644
rect 6174 4644 6192 4662
rect 6174 4662 6192 4680
rect 6174 4680 6192 4698
rect 6174 4698 6192 4716
rect 6174 4716 6192 4734
rect 6174 4734 6192 4752
rect 6174 4752 6192 4770
rect 6174 4770 6192 4788
rect 6174 4788 6192 4806
rect 6174 4806 6192 4824
rect 6174 4824 6192 4842
rect 6174 4842 6192 4860
rect 6174 4860 6192 4878
rect 6174 4878 6192 4896
rect 6174 4896 6192 4914
rect 6174 4914 6192 4932
rect 6174 4932 6192 4950
rect 6174 4950 6192 4968
rect 6174 4968 6192 4986
rect 6174 4986 6192 5004
rect 6174 5004 6192 5022
rect 6174 5022 6192 5040
rect 6174 5040 6192 5058
rect 6174 5058 6192 5076
rect 6174 5076 6192 5094
rect 6174 5094 6192 5112
rect 6174 5112 6192 5130
rect 6174 5130 6192 5148
rect 6174 5148 6192 5166
rect 6174 5166 6192 5184
rect 6174 5184 6192 5202
rect 6174 5202 6192 5220
rect 6174 5220 6192 5238
rect 6174 5238 6192 5256
rect 6174 5256 6192 5274
rect 6174 5274 6192 5292
rect 6174 5292 6192 5310
rect 6174 5310 6192 5328
rect 6174 5328 6192 5346
rect 6174 5346 6192 5364
rect 6174 5364 6192 5382
rect 6174 5382 6192 5400
rect 6174 5400 6192 5418
rect 6174 5418 6192 5436
rect 6174 5436 6192 5454
rect 6174 5454 6192 5472
rect 6174 5472 6192 5490
rect 6174 5490 6192 5508
rect 6174 5508 6192 5526
rect 6174 5526 6192 5544
rect 6174 5832 6192 5850
rect 6174 5850 6192 5868
rect 6174 5868 6192 5886
rect 6174 5886 6192 5904
rect 6174 5904 6192 5922
rect 6174 5922 6192 5940
rect 6174 5940 6192 5958
rect 6174 5958 6192 5976
rect 6174 5976 6192 5994
rect 6174 5994 6192 6012
rect 6174 6012 6192 6030
rect 6174 6030 6192 6048
rect 6174 6048 6192 6066
rect 6174 6066 6192 6084
rect 6174 6084 6192 6102
rect 6174 6102 6192 6120
rect 6174 6120 6192 6138
rect 6174 6138 6192 6156
rect 6174 6156 6192 6174
rect 6174 6174 6192 6192
rect 6174 6192 6192 6210
rect 6174 6210 6192 6228
rect 6174 6228 6192 6246
rect 6174 6246 6192 6264
rect 6174 6264 6192 6282
rect 6174 6282 6192 6300
rect 6174 6300 6192 6318
rect 6174 6318 6192 6336
rect 6174 6336 6192 6354
rect 6174 6354 6192 6372
rect 6174 6372 6192 6390
rect 6174 6390 6192 6408
rect 6174 6408 6192 6426
rect 6174 6426 6192 6444
rect 6174 6444 6192 6462
rect 6174 6462 6192 6480
rect 6174 6480 6192 6498
rect 6174 6498 6192 6516
rect 6174 6516 6192 6534
rect 6174 6534 6192 6552
rect 6174 6552 6192 6570
rect 6174 6570 6192 6588
rect 6174 6588 6192 6606
rect 6174 6606 6192 6624
rect 6174 6624 6192 6642
rect 6174 6642 6192 6660
rect 6174 6660 6192 6678
rect 6174 6678 6192 6696
rect 6174 6696 6192 6714
rect 6174 6714 6192 6732
rect 6174 6732 6192 6750
rect 6174 6750 6192 6768
rect 6174 6768 6192 6786
rect 6174 6786 6192 6804
rect 6174 6804 6192 6822
rect 6174 6822 6192 6840
rect 6174 6840 6192 6858
rect 6174 6858 6192 6876
rect 6174 6876 6192 6894
rect 6174 6894 6192 6912
rect 6174 6912 6192 6930
rect 6174 6930 6192 6948
rect 6174 6948 6192 6966
rect 6174 6966 6192 6984
rect 6174 6984 6192 7002
rect 6174 7002 6192 7020
rect 6174 7020 6192 7038
rect 6174 7038 6192 7056
rect 6174 7056 6192 7074
rect 6174 7074 6192 7092
rect 6174 7092 6192 7110
rect 6174 7110 6192 7128
rect 6174 7128 6192 7146
rect 6174 7146 6192 7164
rect 6174 7164 6192 7182
rect 6174 7182 6192 7200
rect 6174 7200 6192 7218
rect 6174 7218 6192 7236
rect 6174 7236 6192 7254
rect 6174 7254 6192 7272
rect 6174 7272 6192 7290
rect 6174 7290 6192 7308
rect 6174 7308 6192 7326
rect 6174 7326 6192 7344
rect 6174 7344 6192 7362
rect 6174 7362 6192 7380
rect 6174 7380 6192 7398
rect 6174 7398 6192 7416
rect 6174 7416 6192 7434
rect 6174 7434 6192 7452
rect 6174 7452 6192 7470
rect 6174 7470 6192 7488
rect 6174 7488 6192 7506
rect 6174 7506 6192 7524
rect 6174 7524 6192 7542
rect 6174 7542 6192 7560
rect 6174 7560 6192 7578
rect 6174 7578 6192 7596
rect 6174 7596 6192 7614
rect 6174 7614 6192 7632
rect 6174 7632 6192 7650
rect 6174 7650 6192 7668
rect 6174 7668 6192 7686
rect 6174 7686 6192 7704
rect 6174 7704 6192 7722
rect 6174 7722 6192 7740
rect 6174 7740 6192 7758
rect 6174 7758 6192 7776
rect 6174 7776 6192 7794
rect 6174 7794 6192 7812
rect 6174 7812 6192 7830
rect 6174 7830 6192 7848
rect 6174 7848 6192 7866
rect 6174 7866 6192 7884
rect 6174 7884 6192 7902
rect 6174 7902 6192 7920
rect 6174 7920 6192 7938
rect 6174 7938 6192 7956
rect 6174 7956 6192 7974
rect 6174 7974 6192 7992
rect 6174 7992 6192 8010
rect 6174 8010 6192 8028
rect 6174 8028 6192 8046
rect 6174 8046 6192 8064
rect 6174 8064 6192 8082
rect 6174 8082 6192 8100
rect 6174 8100 6192 8118
rect 6174 8118 6192 8136
rect 6174 8136 6192 8154
rect 6174 8154 6192 8172
rect 6174 8172 6192 8190
rect 6174 8190 6192 8208
rect 6174 8208 6192 8226
rect 6174 8226 6192 8244
rect 6174 8244 6192 8262
rect 6174 8262 6192 8280
rect 6174 8280 6192 8298
rect 6174 8298 6192 8316
rect 6174 8316 6192 8334
rect 6174 8334 6192 8352
rect 6174 8352 6192 8370
rect 6174 8370 6192 8388
rect 6174 8388 6192 8406
rect 6174 8406 6192 8424
rect 6174 8424 6192 8442
rect 6174 8442 6192 8460
rect 6174 8460 6192 8478
rect 6174 8478 6192 8496
rect 6174 8496 6192 8514
rect 6174 8514 6192 8532
rect 6174 8532 6192 8550
rect 6174 8550 6192 8568
rect 6174 8568 6192 8586
rect 6174 8586 6192 8604
rect 6174 8604 6192 8622
rect 6174 8622 6192 8640
rect 6174 8640 6192 8658
rect 6174 8658 6192 8676
rect 6174 8676 6192 8694
rect 6174 8694 6192 8712
rect 6174 8712 6192 8730
rect 6174 8730 6192 8748
rect 6174 8748 6192 8766
rect 6174 8766 6192 8784
rect 6174 8784 6192 8802
rect 6174 8802 6192 8820
rect 6174 8820 6192 8838
rect 6174 8838 6192 8856
rect 6174 8856 6192 8874
rect 6174 8874 6192 8892
rect 6174 8892 6192 8910
rect 6174 8910 6192 8928
rect 6174 8928 6192 8946
rect 6174 8946 6192 8964
rect 6174 8964 6192 8982
rect 6174 8982 6192 9000
rect 6174 9000 6192 9018
rect 6174 9018 6192 9036
rect 6174 9036 6192 9054
rect 6174 9054 6192 9072
rect 6174 9072 6192 9090
rect 6174 9090 6192 9108
rect 6174 9108 6192 9126
rect 6174 9126 6192 9144
rect 6174 9144 6192 9162
rect 6174 9162 6192 9180
rect 6174 9180 6192 9198
rect 6174 9198 6192 9216
rect 6174 9216 6192 9234
rect 6174 9234 6192 9252
rect 6174 9252 6192 9270
rect 6174 9270 6192 9288
rect 6174 9288 6192 9306
rect 6174 9306 6192 9324
rect 6174 9324 6192 9342
rect 6174 9342 6192 9360
rect 6174 9360 6192 9378
rect 6174 9378 6192 9396
rect 6174 9396 6192 9414
rect 6174 9414 6192 9432
rect 6174 9432 6192 9450
rect 6192 1080 6210 1098
rect 6192 1098 6210 1116
rect 6192 1116 6210 1134
rect 6192 1134 6210 1152
rect 6192 1152 6210 1170
rect 6192 1332 6210 1350
rect 6192 1350 6210 1368
rect 6192 1368 6210 1386
rect 6192 1386 6210 1404
rect 6192 1404 6210 1422
rect 6192 1422 6210 1440
rect 6192 1440 6210 1458
rect 6192 1458 6210 1476
rect 6192 1476 6210 1494
rect 6192 1494 6210 1512
rect 6192 1512 6210 1530
rect 6192 1530 6210 1548
rect 6192 1548 6210 1566
rect 6192 1566 6210 1584
rect 6192 1584 6210 1602
rect 6192 1602 6210 1620
rect 6192 1620 6210 1638
rect 6192 1638 6210 1656
rect 6192 1656 6210 1674
rect 6192 1674 6210 1692
rect 6192 1692 6210 1710
rect 6192 1710 6210 1728
rect 6192 1728 6210 1746
rect 6192 1746 6210 1764
rect 6192 1764 6210 1782
rect 6192 1782 6210 1800
rect 6192 1800 6210 1818
rect 6192 1818 6210 1836
rect 6192 1836 6210 1854
rect 6192 1854 6210 1872
rect 6192 1872 6210 1890
rect 6192 1890 6210 1908
rect 6192 1908 6210 1926
rect 6192 1926 6210 1944
rect 6192 1944 6210 1962
rect 6192 1962 6210 1980
rect 6192 1980 6210 1998
rect 6192 1998 6210 2016
rect 6192 2016 6210 2034
rect 6192 2034 6210 2052
rect 6192 2052 6210 2070
rect 6192 2070 6210 2088
rect 6192 2088 6210 2106
rect 6192 2106 6210 2124
rect 6192 2124 6210 2142
rect 6192 2142 6210 2160
rect 6192 2160 6210 2178
rect 6192 2178 6210 2196
rect 6192 2196 6210 2214
rect 6192 2214 6210 2232
rect 6192 2232 6210 2250
rect 6192 2250 6210 2268
rect 6192 2268 6210 2286
rect 6192 2286 6210 2304
rect 6192 2304 6210 2322
rect 6192 2322 6210 2340
rect 6192 2340 6210 2358
rect 6192 2358 6210 2376
rect 6192 2376 6210 2394
rect 6192 2394 6210 2412
rect 6192 2412 6210 2430
rect 6192 2430 6210 2448
rect 6192 2448 6210 2466
rect 6192 2466 6210 2484
rect 6192 2484 6210 2502
rect 6192 2502 6210 2520
rect 6192 2520 6210 2538
rect 6192 2538 6210 2556
rect 6192 2556 6210 2574
rect 6192 2574 6210 2592
rect 6192 2592 6210 2610
rect 6192 2610 6210 2628
rect 6192 2628 6210 2646
rect 6192 2646 6210 2664
rect 6192 2664 6210 2682
rect 6192 2682 6210 2700
rect 6192 2700 6210 2718
rect 6192 2718 6210 2736
rect 6192 2736 6210 2754
rect 6192 2754 6210 2772
rect 6192 2772 6210 2790
rect 6192 2790 6210 2808
rect 6192 2808 6210 2826
rect 6192 3078 6210 3096
rect 6192 3096 6210 3114
rect 6192 3114 6210 3132
rect 6192 3132 6210 3150
rect 6192 3150 6210 3168
rect 6192 3168 6210 3186
rect 6192 3186 6210 3204
rect 6192 3204 6210 3222
rect 6192 3222 6210 3240
rect 6192 3240 6210 3258
rect 6192 3258 6210 3276
rect 6192 3276 6210 3294
rect 6192 3294 6210 3312
rect 6192 3312 6210 3330
rect 6192 3330 6210 3348
rect 6192 3348 6210 3366
rect 6192 3366 6210 3384
rect 6192 3384 6210 3402
rect 6192 3402 6210 3420
rect 6192 3420 6210 3438
rect 6192 3438 6210 3456
rect 6192 3456 6210 3474
rect 6192 3474 6210 3492
rect 6192 3492 6210 3510
rect 6192 3510 6210 3528
rect 6192 3528 6210 3546
rect 6192 3546 6210 3564
rect 6192 3564 6210 3582
rect 6192 3582 6210 3600
rect 6192 3600 6210 3618
rect 6192 3618 6210 3636
rect 6192 3636 6210 3654
rect 6192 3654 6210 3672
rect 6192 3672 6210 3690
rect 6192 3690 6210 3708
rect 6192 3708 6210 3726
rect 6192 3726 6210 3744
rect 6192 3744 6210 3762
rect 6192 3762 6210 3780
rect 6192 3780 6210 3798
rect 6192 3798 6210 3816
rect 6192 3816 6210 3834
rect 6192 3834 6210 3852
rect 6192 3852 6210 3870
rect 6192 3870 6210 3888
rect 6192 3888 6210 3906
rect 6192 3906 6210 3924
rect 6192 3924 6210 3942
rect 6192 3942 6210 3960
rect 6192 3960 6210 3978
rect 6192 3978 6210 3996
rect 6192 3996 6210 4014
rect 6192 4014 6210 4032
rect 6192 4032 6210 4050
rect 6192 4050 6210 4068
rect 6192 4068 6210 4086
rect 6192 4086 6210 4104
rect 6192 4104 6210 4122
rect 6192 4122 6210 4140
rect 6192 4140 6210 4158
rect 6192 4158 6210 4176
rect 6192 4176 6210 4194
rect 6192 4194 6210 4212
rect 6192 4212 6210 4230
rect 6192 4230 6210 4248
rect 6192 4248 6210 4266
rect 6192 4266 6210 4284
rect 6192 4284 6210 4302
rect 6192 4302 6210 4320
rect 6192 4320 6210 4338
rect 6192 4338 6210 4356
rect 6192 4356 6210 4374
rect 6192 4374 6210 4392
rect 6192 4392 6210 4410
rect 6192 4410 6210 4428
rect 6192 4428 6210 4446
rect 6192 4446 6210 4464
rect 6192 4464 6210 4482
rect 6192 4482 6210 4500
rect 6192 4500 6210 4518
rect 6192 4518 6210 4536
rect 6192 4536 6210 4554
rect 6192 4554 6210 4572
rect 6192 4572 6210 4590
rect 6192 4590 6210 4608
rect 6192 4608 6210 4626
rect 6192 4626 6210 4644
rect 6192 4644 6210 4662
rect 6192 4662 6210 4680
rect 6192 4680 6210 4698
rect 6192 4698 6210 4716
rect 6192 4716 6210 4734
rect 6192 4734 6210 4752
rect 6192 4752 6210 4770
rect 6192 4770 6210 4788
rect 6192 4788 6210 4806
rect 6192 4806 6210 4824
rect 6192 4824 6210 4842
rect 6192 4842 6210 4860
rect 6192 4860 6210 4878
rect 6192 4878 6210 4896
rect 6192 4896 6210 4914
rect 6192 4914 6210 4932
rect 6192 4932 6210 4950
rect 6192 4950 6210 4968
rect 6192 4968 6210 4986
rect 6192 4986 6210 5004
rect 6192 5004 6210 5022
rect 6192 5022 6210 5040
rect 6192 5040 6210 5058
rect 6192 5058 6210 5076
rect 6192 5076 6210 5094
rect 6192 5094 6210 5112
rect 6192 5112 6210 5130
rect 6192 5130 6210 5148
rect 6192 5148 6210 5166
rect 6192 5166 6210 5184
rect 6192 5184 6210 5202
rect 6192 5202 6210 5220
rect 6192 5220 6210 5238
rect 6192 5238 6210 5256
rect 6192 5256 6210 5274
rect 6192 5274 6210 5292
rect 6192 5292 6210 5310
rect 6192 5310 6210 5328
rect 6192 5328 6210 5346
rect 6192 5346 6210 5364
rect 6192 5364 6210 5382
rect 6192 5382 6210 5400
rect 6192 5400 6210 5418
rect 6192 5418 6210 5436
rect 6192 5436 6210 5454
rect 6192 5454 6210 5472
rect 6192 5472 6210 5490
rect 6192 5490 6210 5508
rect 6192 5508 6210 5526
rect 6192 5526 6210 5544
rect 6192 5544 6210 5562
rect 6192 5868 6210 5886
rect 6192 5886 6210 5904
rect 6192 5904 6210 5922
rect 6192 5922 6210 5940
rect 6192 5940 6210 5958
rect 6192 5958 6210 5976
rect 6192 5976 6210 5994
rect 6192 5994 6210 6012
rect 6192 6012 6210 6030
rect 6192 6030 6210 6048
rect 6192 6048 6210 6066
rect 6192 6066 6210 6084
rect 6192 6084 6210 6102
rect 6192 6102 6210 6120
rect 6192 6120 6210 6138
rect 6192 6138 6210 6156
rect 6192 6156 6210 6174
rect 6192 6174 6210 6192
rect 6192 6192 6210 6210
rect 6192 6210 6210 6228
rect 6192 6228 6210 6246
rect 6192 6246 6210 6264
rect 6192 6264 6210 6282
rect 6192 6282 6210 6300
rect 6192 6300 6210 6318
rect 6192 6318 6210 6336
rect 6192 6336 6210 6354
rect 6192 6354 6210 6372
rect 6192 6372 6210 6390
rect 6192 6390 6210 6408
rect 6192 6408 6210 6426
rect 6192 6426 6210 6444
rect 6192 6444 6210 6462
rect 6192 6462 6210 6480
rect 6192 6480 6210 6498
rect 6192 6498 6210 6516
rect 6192 6516 6210 6534
rect 6192 6534 6210 6552
rect 6192 6552 6210 6570
rect 6192 6570 6210 6588
rect 6192 6588 6210 6606
rect 6192 6606 6210 6624
rect 6192 6624 6210 6642
rect 6192 6642 6210 6660
rect 6192 6660 6210 6678
rect 6192 6678 6210 6696
rect 6192 6696 6210 6714
rect 6192 6714 6210 6732
rect 6192 6732 6210 6750
rect 6192 6750 6210 6768
rect 6192 6768 6210 6786
rect 6192 6786 6210 6804
rect 6192 6804 6210 6822
rect 6192 6822 6210 6840
rect 6192 6840 6210 6858
rect 6192 6858 6210 6876
rect 6192 6876 6210 6894
rect 6192 6894 6210 6912
rect 6192 6912 6210 6930
rect 6192 6930 6210 6948
rect 6192 6948 6210 6966
rect 6192 6966 6210 6984
rect 6192 6984 6210 7002
rect 6192 7002 6210 7020
rect 6192 7020 6210 7038
rect 6192 7038 6210 7056
rect 6192 7056 6210 7074
rect 6192 7074 6210 7092
rect 6192 7092 6210 7110
rect 6192 7110 6210 7128
rect 6192 7128 6210 7146
rect 6192 7146 6210 7164
rect 6192 7164 6210 7182
rect 6192 7182 6210 7200
rect 6192 7200 6210 7218
rect 6192 7218 6210 7236
rect 6192 7236 6210 7254
rect 6192 7254 6210 7272
rect 6192 7272 6210 7290
rect 6192 7290 6210 7308
rect 6192 7308 6210 7326
rect 6192 7326 6210 7344
rect 6192 7344 6210 7362
rect 6192 7362 6210 7380
rect 6192 7380 6210 7398
rect 6192 7398 6210 7416
rect 6192 7416 6210 7434
rect 6192 7434 6210 7452
rect 6192 7452 6210 7470
rect 6192 7470 6210 7488
rect 6192 7488 6210 7506
rect 6192 7506 6210 7524
rect 6192 7524 6210 7542
rect 6192 7542 6210 7560
rect 6192 7560 6210 7578
rect 6192 7578 6210 7596
rect 6192 7596 6210 7614
rect 6192 7614 6210 7632
rect 6192 7632 6210 7650
rect 6192 7650 6210 7668
rect 6192 7668 6210 7686
rect 6192 7686 6210 7704
rect 6192 7704 6210 7722
rect 6192 7722 6210 7740
rect 6192 7740 6210 7758
rect 6192 7758 6210 7776
rect 6192 7776 6210 7794
rect 6192 7794 6210 7812
rect 6192 7812 6210 7830
rect 6192 7830 6210 7848
rect 6192 7848 6210 7866
rect 6192 7866 6210 7884
rect 6192 7884 6210 7902
rect 6192 7902 6210 7920
rect 6192 7920 6210 7938
rect 6192 7938 6210 7956
rect 6192 7956 6210 7974
rect 6192 7974 6210 7992
rect 6192 7992 6210 8010
rect 6192 8010 6210 8028
rect 6192 8028 6210 8046
rect 6192 8046 6210 8064
rect 6192 8064 6210 8082
rect 6192 8082 6210 8100
rect 6192 8100 6210 8118
rect 6192 8118 6210 8136
rect 6192 8136 6210 8154
rect 6192 8154 6210 8172
rect 6192 8172 6210 8190
rect 6192 8190 6210 8208
rect 6192 8208 6210 8226
rect 6192 8226 6210 8244
rect 6192 8244 6210 8262
rect 6192 8262 6210 8280
rect 6192 8280 6210 8298
rect 6192 8298 6210 8316
rect 6192 8316 6210 8334
rect 6192 8334 6210 8352
rect 6192 8352 6210 8370
rect 6192 8370 6210 8388
rect 6192 8388 6210 8406
rect 6192 8406 6210 8424
rect 6192 8424 6210 8442
rect 6192 8442 6210 8460
rect 6192 8460 6210 8478
rect 6192 8478 6210 8496
rect 6192 8496 6210 8514
rect 6192 8514 6210 8532
rect 6192 8532 6210 8550
rect 6192 8550 6210 8568
rect 6192 8568 6210 8586
rect 6192 8586 6210 8604
rect 6192 8604 6210 8622
rect 6192 8622 6210 8640
rect 6192 8640 6210 8658
rect 6192 8658 6210 8676
rect 6192 8676 6210 8694
rect 6192 8694 6210 8712
rect 6192 8712 6210 8730
rect 6192 8730 6210 8748
rect 6192 8748 6210 8766
rect 6192 8766 6210 8784
rect 6192 8784 6210 8802
rect 6192 8802 6210 8820
rect 6192 8820 6210 8838
rect 6192 8838 6210 8856
rect 6192 8856 6210 8874
rect 6192 8874 6210 8892
rect 6192 8892 6210 8910
rect 6192 8910 6210 8928
rect 6192 8928 6210 8946
rect 6192 8946 6210 8964
rect 6192 8964 6210 8982
rect 6192 8982 6210 9000
rect 6192 9000 6210 9018
rect 6192 9018 6210 9036
rect 6192 9036 6210 9054
rect 6192 9054 6210 9072
rect 6192 9072 6210 9090
rect 6192 9090 6210 9108
rect 6192 9108 6210 9126
rect 6192 9126 6210 9144
rect 6192 9144 6210 9162
rect 6192 9162 6210 9180
rect 6192 9180 6210 9198
rect 6192 9198 6210 9216
rect 6192 9216 6210 9234
rect 6192 9234 6210 9252
rect 6192 9252 6210 9270
rect 6192 9270 6210 9288
rect 6192 9288 6210 9306
rect 6192 9306 6210 9324
rect 6192 9324 6210 9342
rect 6192 9342 6210 9360
rect 6192 9360 6210 9378
rect 6192 9378 6210 9396
rect 6192 9396 6210 9414
rect 6192 9414 6210 9432
rect 6192 9432 6210 9450
rect 6192 9450 6210 9468
rect 6192 9468 6210 9486
rect 6210 1098 6228 1116
rect 6210 1116 6228 1134
rect 6210 1134 6228 1152
rect 6210 1152 6228 1170
rect 6210 1170 6228 1188
rect 6210 1332 6228 1350
rect 6210 1350 6228 1368
rect 6210 1368 6228 1386
rect 6210 1386 6228 1404
rect 6210 1404 6228 1422
rect 6210 1422 6228 1440
rect 6210 1440 6228 1458
rect 6210 1458 6228 1476
rect 6210 1476 6228 1494
rect 6210 1494 6228 1512
rect 6210 1512 6228 1530
rect 6210 1530 6228 1548
rect 6210 1548 6228 1566
rect 6210 1566 6228 1584
rect 6210 1584 6228 1602
rect 6210 1602 6228 1620
rect 6210 1620 6228 1638
rect 6210 1638 6228 1656
rect 6210 1656 6228 1674
rect 6210 1674 6228 1692
rect 6210 1692 6228 1710
rect 6210 1710 6228 1728
rect 6210 1728 6228 1746
rect 6210 1746 6228 1764
rect 6210 1764 6228 1782
rect 6210 1782 6228 1800
rect 6210 1800 6228 1818
rect 6210 1818 6228 1836
rect 6210 1836 6228 1854
rect 6210 1854 6228 1872
rect 6210 1872 6228 1890
rect 6210 1890 6228 1908
rect 6210 1908 6228 1926
rect 6210 1926 6228 1944
rect 6210 1944 6228 1962
rect 6210 1962 6228 1980
rect 6210 1980 6228 1998
rect 6210 1998 6228 2016
rect 6210 2016 6228 2034
rect 6210 2034 6228 2052
rect 6210 2052 6228 2070
rect 6210 2070 6228 2088
rect 6210 2088 6228 2106
rect 6210 2106 6228 2124
rect 6210 2124 6228 2142
rect 6210 2142 6228 2160
rect 6210 2160 6228 2178
rect 6210 2178 6228 2196
rect 6210 2196 6228 2214
rect 6210 2214 6228 2232
rect 6210 2232 6228 2250
rect 6210 2250 6228 2268
rect 6210 2268 6228 2286
rect 6210 2286 6228 2304
rect 6210 2304 6228 2322
rect 6210 2322 6228 2340
rect 6210 2340 6228 2358
rect 6210 2358 6228 2376
rect 6210 2376 6228 2394
rect 6210 2394 6228 2412
rect 6210 2412 6228 2430
rect 6210 2430 6228 2448
rect 6210 2448 6228 2466
rect 6210 2466 6228 2484
rect 6210 2484 6228 2502
rect 6210 2502 6228 2520
rect 6210 2520 6228 2538
rect 6210 2538 6228 2556
rect 6210 2556 6228 2574
rect 6210 2574 6228 2592
rect 6210 2592 6228 2610
rect 6210 2610 6228 2628
rect 6210 2628 6228 2646
rect 6210 2646 6228 2664
rect 6210 2664 6228 2682
rect 6210 2682 6228 2700
rect 6210 2700 6228 2718
rect 6210 2718 6228 2736
rect 6210 2736 6228 2754
rect 6210 2754 6228 2772
rect 6210 2772 6228 2790
rect 6210 2790 6228 2808
rect 6210 2808 6228 2826
rect 6210 3096 6228 3114
rect 6210 3114 6228 3132
rect 6210 3132 6228 3150
rect 6210 3150 6228 3168
rect 6210 3168 6228 3186
rect 6210 3186 6228 3204
rect 6210 3204 6228 3222
rect 6210 3222 6228 3240
rect 6210 3240 6228 3258
rect 6210 3258 6228 3276
rect 6210 3276 6228 3294
rect 6210 3294 6228 3312
rect 6210 3312 6228 3330
rect 6210 3330 6228 3348
rect 6210 3348 6228 3366
rect 6210 3366 6228 3384
rect 6210 3384 6228 3402
rect 6210 3402 6228 3420
rect 6210 3420 6228 3438
rect 6210 3438 6228 3456
rect 6210 3456 6228 3474
rect 6210 3474 6228 3492
rect 6210 3492 6228 3510
rect 6210 3510 6228 3528
rect 6210 3528 6228 3546
rect 6210 3546 6228 3564
rect 6210 3564 6228 3582
rect 6210 3582 6228 3600
rect 6210 3600 6228 3618
rect 6210 3618 6228 3636
rect 6210 3636 6228 3654
rect 6210 3654 6228 3672
rect 6210 3672 6228 3690
rect 6210 3690 6228 3708
rect 6210 3708 6228 3726
rect 6210 3726 6228 3744
rect 6210 3744 6228 3762
rect 6210 3762 6228 3780
rect 6210 3780 6228 3798
rect 6210 3798 6228 3816
rect 6210 3816 6228 3834
rect 6210 3834 6228 3852
rect 6210 3852 6228 3870
rect 6210 3870 6228 3888
rect 6210 3888 6228 3906
rect 6210 3906 6228 3924
rect 6210 3924 6228 3942
rect 6210 3942 6228 3960
rect 6210 3960 6228 3978
rect 6210 3978 6228 3996
rect 6210 3996 6228 4014
rect 6210 4014 6228 4032
rect 6210 4032 6228 4050
rect 6210 4050 6228 4068
rect 6210 4068 6228 4086
rect 6210 4086 6228 4104
rect 6210 4104 6228 4122
rect 6210 4122 6228 4140
rect 6210 4140 6228 4158
rect 6210 4158 6228 4176
rect 6210 4176 6228 4194
rect 6210 4194 6228 4212
rect 6210 4212 6228 4230
rect 6210 4230 6228 4248
rect 6210 4248 6228 4266
rect 6210 4266 6228 4284
rect 6210 4284 6228 4302
rect 6210 4302 6228 4320
rect 6210 4320 6228 4338
rect 6210 4338 6228 4356
rect 6210 4356 6228 4374
rect 6210 4374 6228 4392
rect 6210 4392 6228 4410
rect 6210 4410 6228 4428
rect 6210 4428 6228 4446
rect 6210 4446 6228 4464
rect 6210 4464 6228 4482
rect 6210 4482 6228 4500
rect 6210 4500 6228 4518
rect 6210 4518 6228 4536
rect 6210 4536 6228 4554
rect 6210 4554 6228 4572
rect 6210 4572 6228 4590
rect 6210 4590 6228 4608
rect 6210 4608 6228 4626
rect 6210 4626 6228 4644
rect 6210 4644 6228 4662
rect 6210 4662 6228 4680
rect 6210 4680 6228 4698
rect 6210 4698 6228 4716
rect 6210 4716 6228 4734
rect 6210 4734 6228 4752
rect 6210 4752 6228 4770
rect 6210 4770 6228 4788
rect 6210 4788 6228 4806
rect 6210 4806 6228 4824
rect 6210 4824 6228 4842
rect 6210 4842 6228 4860
rect 6210 4860 6228 4878
rect 6210 4878 6228 4896
rect 6210 4896 6228 4914
rect 6210 4914 6228 4932
rect 6210 4932 6228 4950
rect 6210 4950 6228 4968
rect 6210 4968 6228 4986
rect 6210 4986 6228 5004
rect 6210 5004 6228 5022
rect 6210 5022 6228 5040
rect 6210 5040 6228 5058
rect 6210 5058 6228 5076
rect 6210 5076 6228 5094
rect 6210 5094 6228 5112
rect 6210 5112 6228 5130
rect 6210 5130 6228 5148
rect 6210 5148 6228 5166
rect 6210 5166 6228 5184
rect 6210 5184 6228 5202
rect 6210 5202 6228 5220
rect 6210 5220 6228 5238
rect 6210 5238 6228 5256
rect 6210 5256 6228 5274
rect 6210 5274 6228 5292
rect 6210 5292 6228 5310
rect 6210 5310 6228 5328
rect 6210 5328 6228 5346
rect 6210 5346 6228 5364
rect 6210 5364 6228 5382
rect 6210 5382 6228 5400
rect 6210 5400 6228 5418
rect 6210 5418 6228 5436
rect 6210 5436 6228 5454
rect 6210 5454 6228 5472
rect 6210 5472 6228 5490
rect 6210 5490 6228 5508
rect 6210 5508 6228 5526
rect 6210 5526 6228 5544
rect 6210 5544 6228 5562
rect 6210 5562 6228 5580
rect 6210 5904 6228 5922
rect 6210 5922 6228 5940
rect 6210 5940 6228 5958
rect 6210 5958 6228 5976
rect 6210 5976 6228 5994
rect 6210 5994 6228 6012
rect 6210 6012 6228 6030
rect 6210 6030 6228 6048
rect 6210 6048 6228 6066
rect 6210 6066 6228 6084
rect 6210 6084 6228 6102
rect 6210 6102 6228 6120
rect 6210 6120 6228 6138
rect 6210 6138 6228 6156
rect 6210 6156 6228 6174
rect 6210 6174 6228 6192
rect 6210 6192 6228 6210
rect 6210 6210 6228 6228
rect 6210 6228 6228 6246
rect 6210 6246 6228 6264
rect 6210 6264 6228 6282
rect 6210 6282 6228 6300
rect 6210 6300 6228 6318
rect 6210 6318 6228 6336
rect 6210 6336 6228 6354
rect 6210 6354 6228 6372
rect 6210 6372 6228 6390
rect 6210 6390 6228 6408
rect 6210 6408 6228 6426
rect 6210 6426 6228 6444
rect 6210 6444 6228 6462
rect 6210 6462 6228 6480
rect 6210 6480 6228 6498
rect 6210 6498 6228 6516
rect 6210 6516 6228 6534
rect 6210 6534 6228 6552
rect 6210 6552 6228 6570
rect 6210 6570 6228 6588
rect 6210 6588 6228 6606
rect 6210 6606 6228 6624
rect 6210 6624 6228 6642
rect 6210 6642 6228 6660
rect 6210 6660 6228 6678
rect 6210 6678 6228 6696
rect 6210 6696 6228 6714
rect 6210 6714 6228 6732
rect 6210 6732 6228 6750
rect 6210 6750 6228 6768
rect 6210 6768 6228 6786
rect 6210 6786 6228 6804
rect 6210 6804 6228 6822
rect 6210 6822 6228 6840
rect 6210 6840 6228 6858
rect 6210 6858 6228 6876
rect 6210 6876 6228 6894
rect 6210 6894 6228 6912
rect 6210 6912 6228 6930
rect 6210 6930 6228 6948
rect 6210 6948 6228 6966
rect 6210 6966 6228 6984
rect 6210 6984 6228 7002
rect 6210 7002 6228 7020
rect 6210 7020 6228 7038
rect 6210 7038 6228 7056
rect 6210 7056 6228 7074
rect 6210 7074 6228 7092
rect 6210 7092 6228 7110
rect 6210 7110 6228 7128
rect 6210 7128 6228 7146
rect 6210 7146 6228 7164
rect 6210 7164 6228 7182
rect 6210 7182 6228 7200
rect 6210 7200 6228 7218
rect 6210 7218 6228 7236
rect 6210 7236 6228 7254
rect 6210 7254 6228 7272
rect 6210 7272 6228 7290
rect 6210 7290 6228 7308
rect 6210 7308 6228 7326
rect 6210 7326 6228 7344
rect 6210 7344 6228 7362
rect 6210 7362 6228 7380
rect 6210 7380 6228 7398
rect 6210 7398 6228 7416
rect 6210 7416 6228 7434
rect 6210 7434 6228 7452
rect 6210 7452 6228 7470
rect 6210 7470 6228 7488
rect 6210 7488 6228 7506
rect 6210 7506 6228 7524
rect 6210 7524 6228 7542
rect 6210 7542 6228 7560
rect 6210 7560 6228 7578
rect 6210 7578 6228 7596
rect 6210 7596 6228 7614
rect 6210 7614 6228 7632
rect 6210 7632 6228 7650
rect 6210 7650 6228 7668
rect 6210 7668 6228 7686
rect 6210 7686 6228 7704
rect 6210 7704 6228 7722
rect 6210 7722 6228 7740
rect 6210 7740 6228 7758
rect 6210 7758 6228 7776
rect 6210 7776 6228 7794
rect 6210 7794 6228 7812
rect 6210 7812 6228 7830
rect 6210 7830 6228 7848
rect 6210 7848 6228 7866
rect 6210 7866 6228 7884
rect 6210 7884 6228 7902
rect 6210 7902 6228 7920
rect 6210 7920 6228 7938
rect 6210 7938 6228 7956
rect 6210 7956 6228 7974
rect 6210 7974 6228 7992
rect 6210 7992 6228 8010
rect 6210 8010 6228 8028
rect 6210 8028 6228 8046
rect 6210 8046 6228 8064
rect 6210 8064 6228 8082
rect 6210 8082 6228 8100
rect 6210 8100 6228 8118
rect 6210 8118 6228 8136
rect 6210 8136 6228 8154
rect 6210 8154 6228 8172
rect 6210 8172 6228 8190
rect 6210 8190 6228 8208
rect 6210 8208 6228 8226
rect 6210 8226 6228 8244
rect 6210 8244 6228 8262
rect 6210 8262 6228 8280
rect 6210 8280 6228 8298
rect 6210 8298 6228 8316
rect 6210 8316 6228 8334
rect 6210 8334 6228 8352
rect 6210 8352 6228 8370
rect 6210 8370 6228 8388
rect 6210 8388 6228 8406
rect 6210 8406 6228 8424
rect 6210 8424 6228 8442
rect 6210 8442 6228 8460
rect 6210 8460 6228 8478
rect 6210 8478 6228 8496
rect 6210 8496 6228 8514
rect 6210 8514 6228 8532
rect 6210 8532 6228 8550
rect 6210 8550 6228 8568
rect 6210 8568 6228 8586
rect 6210 8586 6228 8604
rect 6210 8604 6228 8622
rect 6210 8622 6228 8640
rect 6210 8640 6228 8658
rect 6210 8658 6228 8676
rect 6210 8676 6228 8694
rect 6210 8694 6228 8712
rect 6210 8712 6228 8730
rect 6210 8730 6228 8748
rect 6210 8748 6228 8766
rect 6210 8766 6228 8784
rect 6210 8784 6228 8802
rect 6210 8802 6228 8820
rect 6210 8820 6228 8838
rect 6210 8838 6228 8856
rect 6210 8856 6228 8874
rect 6210 8874 6228 8892
rect 6210 8892 6228 8910
rect 6210 8910 6228 8928
rect 6210 8928 6228 8946
rect 6210 8946 6228 8964
rect 6210 8964 6228 8982
rect 6210 8982 6228 9000
rect 6210 9000 6228 9018
rect 6210 9018 6228 9036
rect 6210 9036 6228 9054
rect 6210 9054 6228 9072
rect 6210 9072 6228 9090
rect 6210 9090 6228 9108
rect 6210 9108 6228 9126
rect 6210 9126 6228 9144
rect 6210 9144 6228 9162
rect 6210 9162 6228 9180
rect 6210 9180 6228 9198
rect 6210 9198 6228 9216
rect 6210 9216 6228 9234
rect 6210 9234 6228 9252
rect 6210 9252 6228 9270
rect 6210 9270 6228 9288
rect 6210 9288 6228 9306
rect 6210 9306 6228 9324
rect 6210 9324 6228 9342
rect 6210 9342 6228 9360
rect 6210 9360 6228 9378
rect 6210 9378 6228 9396
rect 6210 9396 6228 9414
rect 6210 9414 6228 9432
rect 6210 9432 6228 9450
rect 6210 9450 6228 9468
rect 6210 9468 6228 9486
rect 6210 9486 6228 9504
rect 6228 1116 6246 1134
rect 6228 1134 6246 1152
rect 6228 1152 6246 1170
rect 6228 1170 6246 1188
rect 6228 1350 6246 1368
rect 6228 1368 6246 1386
rect 6228 1386 6246 1404
rect 6228 1404 6246 1422
rect 6228 1422 6246 1440
rect 6228 1440 6246 1458
rect 6228 1458 6246 1476
rect 6228 1476 6246 1494
rect 6228 1494 6246 1512
rect 6228 1512 6246 1530
rect 6228 1530 6246 1548
rect 6228 1548 6246 1566
rect 6228 1566 6246 1584
rect 6228 1584 6246 1602
rect 6228 1602 6246 1620
rect 6228 1620 6246 1638
rect 6228 1638 6246 1656
rect 6228 1656 6246 1674
rect 6228 1674 6246 1692
rect 6228 1692 6246 1710
rect 6228 1710 6246 1728
rect 6228 1728 6246 1746
rect 6228 1746 6246 1764
rect 6228 1764 6246 1782
rect 6228 1782 6246 1800
rect 6228 1800 6246 1818
rect 6228 1818 6246 1836
rect 6228 1836 6246 1854
rect 6228 1854 6246 1872
rect 6228 1872 6246 1890
rect 6228 1890 6246 1908
rect 6228 1908 6246 1926
rect 6228 1926 6246 1944
rect 6228 1944 6246 1962
rect 6228 1962 6246 1980
rect 6228 1980 6246 1998
rect 6228 1998 6246 2016
rect 6228 2016 6246 2034
rect 6228 2034 6246 2052
rect 6228 2052 6246 2070
rect 6228 2070 6246 2088
rect 6228 2088 6246 2106
rect 6228 2106 6246 2124
rect 6228 2124 6246 2142
rect 6228 2142 6246 2160
rect 6228 2160 6246 2178
rect 6228 2178 6246 2196
rect 6228 2196 6246 2214
rect 6228 2214 6246 2232
rect 6228 2232 6246 2250
rect 6228 2250 6246 2268
rect 6228 2268 6246 2286
rect 6228 2286 6246 2304
rect 6228 2304 6246 2322
rect 6228 2322 6246 2340
rect 6228 2340 6246 2358
rect 6228 2358 6246 2376
rect 6228 2376 6246 2394
rect 6228 2394 6246 2412
rect 6228 2412 6246 2430
rect 6228 2430 6246 2448
rect 6228 2448 6246 2466
rect 6228 2466 6246 2484
rect 6228 2484 6246 2502
rect 6228 2502 6246 2520
rect 6228 2520 6246 2538
rect 6228 2538 6246 2556
rect 6228 2556 6246 2574
rect 6228 2574 6246 2592
rect 6228 2592 6246 2610
rect 6228 2610 6246 2628
rect 6228 2628 6246 2646
rect 6228 2646 6246 2664
rect 6228 2664 6246 2682
rect 6228 2682 6246 2700
rect 6228 2700 6246 2718
rect 6228 2718 6246 2736
rect 6228 2736 6246 2754
rect 6228 2754 6246 2772
rect 6228 2772 6246 2790
rect 6228 2790 6246 2808
rect 6228 2808 6246 2826
rect 6228 2826 6246 2844
rect 6228 3096 6246 3114
rect 6228 3114 6246 3132
rect 6228 3132 6246 3150
rect 6228 3150 6246 3168
rect 6228 3168 6246 3186
rect 6228 3186 6246 3204
rect 6228 3204 6246 3222
rect 6228 3222 6246 3240
rect 6228 3240 6246 3258
rect 6228 3258 6246 3276
rect 6228 3276 6246 3294
rect 6228 3294 6246 3312
rect 6228 3312 6246 3330
rect 6228 3330 6246 3348
rect 6228 3348 6246 3366
rect 6228 3366 6246 3384
rect 6228 3384 6246 3402
rect 6228 3402 6246 3420
rect 6228 3420 6246 3438
rect 6228 3438 6246 3456
rect 6228 3456 6246 3474
rect 6228 3474 6246 3492
rect 6228 3492 6246 3510
rect 6228 3510 6246 3528
rect 6228 3528 6246 3546
rect 6228 3546 6246 3564
rect 6228 3564 6246 3582
rect 6228 3582 6246 3600
rect 6228 3600 6246 3618
rect 6228 3618 6246 3636
rect 6228 3636 6246 3654
rect 6228 3654 6246 3672
rect 6228 3672 6246 3690
rect 6228 3690 6246 3708
rect 6228 3708 6246 3726
rect 6228 3726 6246 3744
rect 6228 3744 6246 3762
rect 6228 3762 6246 3780
rect 6228 3780 6246 3798
rect 6228 3798 6246 3816
rect 6228 3816 6246 3834
rect 6228 3834 6246 3852
rect 6228 3852 6246 3870
rect 6228 3870 6246 3888
rect 6228 3888 6246 3906
rect 6228 3906 6246 3924
rect 6228 3924 6246 3942
rect 6228 3942 6246 3960
rect 6228 3960 6246 3978
rect 6228 3978 6246 3996
rect 6228 3996 6246 4014
rect 6228 4014 6246 4032
rect 6228 4032 6246 4050
rect 6228 4050 6246 4068
rect 6228 4068 6246 4086
rect 6228 4086 6246 4104
rect 6228 4104 6246 4122
rect 6228 4122 6246 4140
rect 6228 4140 6246 4158
rect 6228 4158 6246 4176
rect 6228 4176 6246 4194
rect 6228 4194 6246 4212
rect 6228 4212 6246 4230
rect 6228 4230 6246 4248
rect 6228 4248 6246 4266
rect 6228 4266 6246 4284
rect 6228 4284 6246 4302
rect 6228 4302 6246 4320
rect 6228 4320 6246 4338
rect 6228 4338 6246 4356
rect 6228 4356 6246 4374
rect 6228 4374 6246 4392
rect 6228 4392 6246 4410
rect 6228 4410 6246 4428
rect 6228 4428 6246 4446
rect 6228 4446 6246 4464
rect 6228 4464 6246 4482
rect 6228 4482 6246 4500
rect 6228 4500 6246 4518
rect 6228 4518 6246 4536
rect 6228 4536 6246 4554
rect 6228 4554 6246 4572
rect 6228 4572 6246 4590
rect 6228 4590 6246 4608
rect 6228 4608 6246 4626
rect 6228 4626 6246 4644
rect 6228 4644 6246 4662
rect 6228 4662 6246 4680
rect 6228 4680 6246 4698
rect 6228 4698 6246 4716
rect 6228 4716 6246 4734
rect 6228 4734 6246 4752
rect 6228 4752 6246 4770
rect 6228 4770 6246 4788
rect 6228 4788 6246 4806
rect 6228 4806 6246 4824
rect 6228 4824 6246 4842
rect 6228 4842 6246 4860
rect 6228 4860 6246 4878
rect 6228 4878 6246 4896
rect 6228 4896 6246 4914
rect 6228 4914 6246 4932
rect 6228 4932 6246 4950
rect 6228 4950 6246 4968
rect 6228 4968 6246 4986
rect 6228 4986 6246 5004
rect 6228 5004 6246 5022
rect 6228 5022 6246 5040
rect 6228 5040 6246 5058
rect 6228 5058 6246 5076
rect 6228 5076 6246 5094
rect 6228 5094 6246 5112
rect 6228 5112 6246 5130
rect 6228 5130 6246 5148
rect 6228 5148 6246 5166
rect 6228 5166 6246 5184
rect 6228 5184 6246 5202
rect 6228 5202 6246 5220
rect 6228 5220 6246 5238
rect 6228 5238 6246 5256
rect 6228 5256 6246 5274
rect 6228 5274 6246 5292
rect 6228 5292 6246 5310
rect 6228 5310 6246 5328
rect 6228 5328 6246 5346
rect 6228 5346 6246 5364
rect 6228 5364 6246 5382
rect 6228 5382 6246 5400
rect 6228 5400 6246 5418
rect 6228 5418 6246 5436
rect 6228 5436 6246 5454
rect 6228 5454 6246 5472
rect 6228 5472 6246 5490
rect 6228 5490 6246 5508
rect 6228 5508 6246 5526
rect 6228 5526 6246 5544
rect 6228 5544 6246 5562
rect 6228 5562 6246 5580
rect 6228 5580 6246 5598
rect 6228 5958 6246 5976
rect 6228 5976 6246 5994
rect 6228 5994 6246 6012
rect 6228 6012 6246 6030
rect 6228 6030 6246 6048
rect 6228 6048 6246 6066
rect 6228 6066 6246 6084
rect 6228 6084 6246 6102
rect 6228 6102 6246 6120
rect 6228 6120 6246 6138
rect 6228 6138 6246 6156
rect 6228 6156 6246 6174
rect 6228 6174 6246 6192
rect 6228 6192 6246 6210
rect 6228 6210 6246 6228
rect 6228 6228 6246 6246
rect 6228 6246 6246 6264
rect 6228 6264 6246 6282
rect 6228 6282 6246 6300
rect 6228 6300 6246 6318
rect 6228 6318 6246 6336
rect 6228 6336 6246 6354
rect 6228 6354 6246 6372
rect 6228 6372 6246 6390
rect 6228 6390 6246 6408
rect 6228 6408 6246 6426
rect 6228 6426 6246 6444
rect 6228 6444 6246 6462
rect 6228 6462 6246 6480
rect 6228 6480 6246 6498
rect 6228 6498 6246 6516
rect 6228 6516 6246 6534
rect 6228 6534 6246 6552
rect 6228 6552 6246 6570
rect 6228 6570 6246 6588
rect 6228 6588 6246 6606
rect 6228 6606 6246 6624
rect 6228 6624 6246 6642
rect 6228 6642 6246 6660
rect 6228 6660 6246 6678
rect 6228 6678 6246 6696
rect 6228 6696 6246 6714
rect 6228 6714 6246 6732
rect 6228 6732 6246 6750
rect 6228 6750 6246 6768
rect 6228 6768 6246 6786
rect 6228 6786 6246 6804
rect 6228 6804 6246 6822
rect 6228 6822 6246 6840
rect 6228 6840 6246 6858
rect 6228 6858 6246 6876
rect 6228 6876 6246 6894
rect 6228 6894 6246 6912
rect 6228 6912 6246 6930
rect 6228 6930 6246 6948
rect 6228 6948 6246 6966
rect 6228 6966 6246 6984
rect 6228 6984 6246 7002
rect 6228 7002 6246 7020
rect 6228 7020 6246 7038
rect 6228 7038 6246 7056
rect 6228 7056 6246 7074
rect 6228 7074 6246 7092
rect 6228 7092 6246 7110
rect 6228 7110 6246 7128
rect 6228 7128 6246 7146
rect 6228 7146 6246 7164
rect 6228 7164 6246 7182
rect 6228 7182 6246 7200
rect 6228 7200 6246 7218
rect 6228 7218 6246 7236
rect 6228 7236 6246 7254
rect 6228 7254 6246 7272
rect 6228 7272 6246 7290
rect 6228 7290 6246 7308
rect 6228 7308 6246 7326
rect 6228 7326 6246 7344
rect 6228 7344 6246 7362
rect 6228 7362 6246 7380
rect 6228 7380 6246 7398
rect 6228 7398 6246 7416
rect 6228 7416 6246 7434
rect 6228 7434 6246 7452
rect 6228 7452 6246 7470
rect 6228 7470 6246 7488
rect 6228 7488 6246 7506
rect 6228 7506 6246 7524
rect 6228 7524 6246 7542
rect 6228 7542 6246 7560
rect 6228 7560 6246 7578
rect 6228 7578 6246 7596
rect 6228 7596 6246 7614
rect 6228 7614 6246 7632
rect 6228 7632 6246 7650
rect 6228 7650 6246 7668
rect 6228 7668 6246 7686
rect 6228 7686 6246 7704
rect 6228 7704 6246 7722
rect 6228 7722 6246 7740
rect 6228 7740 6246 7758
rect 6228 7758 6246 7776
rect 6228 7776 6246 7794
rect 6228 7794 6246 7812
rect 6228 7812 6246 7830
rect 6228 7830 6246 7848
rect 6228 7848 6246 7866
rect 6228 7866 6246 7884
rect 6228 7884 6246 7902
rect 6228 7902 6246 7920
rect 6228 7920 6246 7938
rect 6228 7938 6246 7956
rect 6228 7956 6246 7974
rect 6228 7974 6246 7992
rect 6228 7992 6246 8010
rect 6228 8010 6246 8028
rect 6228 8028 6246 8046
rect 6228 8046 6246 8064
rect 6228 8064 6246 8082
rect 6228 8082 6246 8100
rect 6228 8100 6246 8118
rect 6228 8118 6246 8136
rect 6228 8136 6246 8154
rect 6228 8154 6246 8172
rect 6228 8172 6246 8190
rect 6228 8190 6246 8208
rect 6228 8208 6246 8226
rect 6228 8226 6246 8244
rect 6228 8244 6246 8262
rect 6228 8262 6246 8280
rect 6228 8280 6246 8298
rect 6228 8298 6246 8316
rect 6228 8316 6246 8334
rect 6228 8334 6246 8352
rect 6228 8352 6246 8370
rect 6228 8370 6246 8388
rect 6228 8388 6246 8406
rect 6228 8406 6246 8424
rect 6228 8424 6246 8442
rect 6228 8442 6246 8460
rect 6228 8460 6246 8478
rect 6228 8478 6246 8496
rect 6228 8496 6246 8514
rect 6228 8514 6246 8532
rect 6228 8532 6246 8550
rect 6228 8550 6246 8568
rect 6228 8568 6246 8586
rect 6228 8586 6246 8604
rect 6228 8604 6246 8622
rect 6228 8622 6246 8640
rect 6228 8640 6246 8658
rect 6228 8658 6246 8676
rect 6228 8676 6246 8694
rect 6228 8694 6246 8712
rect 6228 8712 6246 8730
rect 6228 8730 6246 8748
rect 6228 8748 6246 8766
rect 6228 8766 6246 8784
rect 6228 8784 6246 8802
rect 6228 8802 6246 8820
rect 6228 8820 6246 8838
rect 6228 8838 6246 8856
rect 6228 8856 6246 8874
rect 6228 8874 6246 8892
rect 6228 8892 6246 8910
rect 6228 8910 6246 8928
rect 6228 8928 6246 8946
rect 6228 8946 6246 8964
rect 6228 8964 6246 8982
rect 6228 8982 6246 9000
rect 6228 9000 6246 9018
rect 6228 9018 6246 9036
rect 6228 9036 6246 9054
rect 6228 9054 6246 9072
rect 6228 9072 6246 9090
rect 6228 9090 6246 9108
rect 6228 9108 6246 9126
rect 6228 9126 6246 9144
rect 6228 9144 6246 9162
rect 6228 9162 6246 9180
rect 6228 9180 6246 9198
rect 6228 9198 6246 9216
rect 6228 9216 6246 9234
rect 6228 9234 6246 9252
rect 6228 9252 6246 9270
rect 6228 9270 6246 9288
rect 6228 9288 6246 9306
rect 6228 9306 6246 9324
rect 6228 9324 6246 9342
rect 6228 9342 6246 9360
rect 6228 9360 6246 9378
rect 6228 9378 6246 9396
rect 6228 9396 6246 9414
rect 6228 9414 6246 9432
rect 6228 9432 6246 9450
rect 6228 9450 6246 9468
rect 6228 9468 6246 9486
rect 6228 9486 6246 9504
rect 6228 9504 6246 9522
rect 6246 1134 6264 1152
rect 6246 1152 6264 1170
rect 6246 1170 6264 1188
rect 6246 1188 6264 1206
rect 6246 1350 6264 1368
rect 6246 1368 6264 1386
rect 6246 1386 6264 1404
rect 6246 1404 6264 1422
rect 6246 1422 6264 1440
rect 6246 1440 6264 1458
rect 6246 1458 6264 1476
rect 6246 1476 6264 1494
rect 6246 1494 6264 1512
rect 6246 1512 6264 1530
rect 6246 1530 6264 1548
rect 6246 1548 6264 1566
rect 6246 1566 6264 1584
rect 6246 1584 6264 1602
rect 6246 1602 6264 1620
rect 6246 1620 6264 1638
rect 6246 1638 6264 1656
rect 6246 1656 6264 1674
rect 6246 1674 6264 1692
rect 6246 1692 6264 1710
rect 6246 1710 6264 1728
rect 6246 1728 6264 1746
rect 6246 1746 6264 1764
rect 6246 1764 6264 1782
rect 6246 1782 6264 1800
rect 6246 1800 6264 1818
rect 6246 1818 6264 1836
rect 6246 1836 6264 1854
rect 6246 1854 6264 1872
rect 6246 1872 6264 1890
rect 6246 1890 6264 1908
rect 6246 1908 6264 1926
rect 6246 1926 6264 1944
rect 6246 1944 6264 1962
rect 6246 1962 6264 1980
rect 6246 1980 6264 1998
rect 6246 1998 6264 2016
rect 6246 2016 6264 2034
rect 6246 2034 6264 2052
rect 6246 2052 6264 2070
rect 6246 2070 6264 2088
rect 6246 2088 6264 2106
rect 6246 2106 6264 2124
rect 6246 2124 6264 2142
rect 6246 2142 6264 2160
rect 6246 2160 6264 2178
rect 6246 2178 6264 2196
rect 6246 2196 6264 2214
rect 6246 2214 6264 2232
rect 6246 2232 6264 2250
rect 6246 2250 6264 2268
rect 6246 2268 6264 2286
rect 6246 2286 6264 2304
rect 6246 2304 6264 2322
rect 6246 2322 6264 2340
rect 6246 2340 6264 2358
rect 6246 2358 6264 2376
rect 6246 2376 6264 2394
rect 6246 2394 6264 2412
rect 6246 2412 6264 2430
rect 6246 2430 6264 2448
rect 6246 2448 6264 2466
rect 6246 2466 6264 2484
rect 6246 2484 6264 2502
rect 6246 2502 6264 2520
rect 6246 2520 6264 2538
rect 6246 2538 6264 2556
rect 6246 2556 6264 2574
rect 6246 2574 6264 2592
rect 6246 2592 6264 2610
rect 6246 2610 6264 2628
rect 6246 2628 6264 2646
rect 6246 2646 6264 2664
rect 6246 2664 6264 2682
rect 6246 2682 6264 2700
rect 6246 2700 6264 2718
rect 6246 2718 6264 2736
rect 6246 2736 6264 2754
rect 6246 2754 6264 2772
rect 6246 2772 6264 2790
rect 6246 2790 6264 2808
rect 6246 2808 6264 2826
rect 6246 2826 6264 2844
rect 6246 3114 6264 3132
rect 6246 3132 6264 3150
rect 6246 3150 6264 3168
rect 6246 3168 6264 3186
rect 6246 3186 6264 3204
rect 6246 3204 6264 3222
rect 6246 3222 6264 3240
rect 6246 3240 6264 3258
rect 6246 3258 6264 3276
rect 6246 3276 6264 3294
rect 6246 3294 6264 3312
rect 6246 3312 6264 3330
rect 6246 3330 6264 3348
rect 6246 3348 6264 3366
rect 6246 3366 6264 3384
rect 6246 3384 6264 3402
rect 6246 3402 6264 3420
rect 6246 3420 6264 3438
rect 6246 3438 6264 3456
rect 6246 3456 6264 3474
rect 6246 3474 6264 3492
rect 6246 3492 6264 3510
rect 6246 3510 6264 3528
rect 6246 3528 6264 3546
rect 6246 3546 6264 3564
rect 6246 3564 6264 3582
rect 6246 3582 6264 3600
rect 6246 3600 6264 3618
rect 6246 3618 6264 3636
rect 6246 3636 6264 3654
rect 6246 3654 6264 3672
rect 6246 3672 6264 3690
rect 6246 3690 6264 3708
rect 6246 3708 6264 3726
rect 6246 3726 6264 3744
rect 6246 3744 6264 3762
rect 6246 3762 6264 3780
rect 6246 3780 6264 3798
rect 6246 3798 6264 3816
rect 6246 3816 6264 3834
rect 6246 3834 6264 3852
rect 6246 3852 6264 3870
rect 6246 3870 6264 3888
rect 6246 3888 6264 3906
rect 6246 3906 6264 3924
rect 6246 3924 6264 3942
rect 6246 3942 6264 3960
rect 6246 3960 6264 3978
rect 6246 3978 6264 3996
rect 6246 3996 6264 4014
rect 6246 4014 6264 4032
rect 6246 4032 6264 4050
rect 6246 4050 6264 4068
rect 6246 4068 6264 4086
rect 6246 4086 6264 4104
rect 6246 4104 6264 4122
rect 6246 4122 6264 4140
rect 6246 4140 6264 4158
rect 6246 4158 6264 4176
rect 6246 4176 6264 4194
rect 6246 4194 6264 4212
rect 6246 4212 6264 4230
rect 6246 4230 6264 4248
rect 6246 4248 6264 4266
rect 6246 4266 6264 4284
rect 6246 4284 6264 4302
rect 6246 4302 6264 4320
rect 6246 4320 6264 4338
rect 6246 4338 6264 4356
rect 6246 4356 6264 4374
rect 6246 4374 6264 4392
rect 6246 4392 6264 4410
rect 6246 4410 6264 4428
rect 6246 4428 6264 4446
rect 6246 4446 6264 4464
rect 6246 4464 6264 4482
rect 6246 4482 6264 4500
rect 6246 4500 6264 4518
rect 6246 4518 6264 4536
rect 6246 4536 6264 4554
rect 6246 4554 6264 4572
rect 6246 4572 6264 4590
rect 6246 4590 6264 4608
rect 6246 4608 6264 4626
rect 6246 4626 6264 4644
rect 6246 4644 6264 4662
rect 6246 4662 6264 4680
rect 6246 4680 6264 4698
rect 6246 4698 6264 4716
rect 6246 4716 6264 4734
rect 6246 4734 6264 4752
rect 6246 4752 6264 4770
rect 6246 4770 6264 4788
rect 6246 4788 6264 4806
rect 6246 4806 6264 4824
rect 6246 4824 6264 4842
rect 6246 4842 6264 4860
rect 6246 4860 6264 4878
rect 6246 4878 6264 4896
rect 6246 4896 6264 4914
rect 6246 4914 6264 4932
rect 6246 4932 6264 4950
rect 6246 4950 6264 4968
rect 6246 4968 6264 4986
rect 6246 4986 6264 5004
rect 6246 5004 6264 5022
rect 6246 5022 6264 5040
rect 6246 5040 6264 5058
rect 6246 5058 6264 5076
rect 6246 5076 6264 5094
rect 6246 5094 6264 5112
rect 6246 5112 6264 5130
rect 6246 5130 6264 5148
rect 6246 5148 6264 5166
rect 6246 5166 6264 5184
rect 6246 5184 6264 5202
rect 6246 5202 6264 5220
rect 6246 5220 6264 5238
rect 6246 5238 6264 5256
rect 6246 5256 6264 5274
rect 6246 5274 6264 5292
rect 6246 5292 6264 5310
rect 6246 5310 6264 5328
rect 6246 5328 6264 5346
rect 6246 5346 6264 5364
rect 6246 5364 6264 5382
rect 6246 5382 6264 5400
rect 6246 5400 6264 5418
rect 6246 5418 6264 5436
rect 6246 5436 6264 5454
rect 6246 5454 6264 5472
rect 6246 5472 6264 5490
rect 6246 5490 6264 5508
rect 6246 5508 6264 5526
rect 6246 5526 6264 5544
rect 6246 5544 6264 5562
rect 6246 5562 6264 5580
rect 6246 5580 6264 5598
rect 6246 5598 6264 5616
rect 6246 5994 6264 6012
rect 6246 6012 6264 6030
rect 6246 6030 6264 6048
rect 6246 6048 6264 6066
rect 6246 6066 6264 6084
rect 6246 6084 6264 6102
rect 6246 6102 6264 6120
rect 6246 6120 6264 6138
rect 6246 6138 6264 6156
rect 6246 6156 6264 6174
rect 6246 6174 6264 6192
rect 6246 6192 6264 6210
rect 6246 6210 6264 6228
rect 6246 6228 6264 6246
rect 6246 6246 6264 6264
rect 6246 6264 6264 6282
rect 6246 6282 6264 6300
rect 6246 6300 6264 6318
rect 6246 6318 6264 6336
rect 6246 6336 6264 6354
rect 6246 6354 6264 6372
rect 6246 6372 6264 6390
rect 6246 6390 6264 6408
rect 6246 6408 6264 6426
rect 6246 6426 6264 6444
rect 6246 6444 6264 6462
rect 6246 6462 6264 6480
rect 6246 6480 6264 6498
rect 6246 6498 6264 6516
rect 6246 6516 6264 6534
rect 6246 6534 6264 6552
rect 6246 6552 6264 6570
rect 6246 6570 6264 6588
rect 6246 6588 6264 6606
rect 6246 6606 6264 6624
rect 6246 6624 6264 6642
rect 6246 6642 6264 6660
rect 6246 6660 6264 6678
rect 6246 6678 6264 6696
rect 6246 6696 6264 6714
rect 6246 6714 6264 6732
rect 6246 6732 6264 6750
rect 6246 6750 6264 6768
rect 6246 6768 6264 6786
rect 6246 6786 6264 6804
rect 6246 6804 6264 6822
rect 6246 6822 6264 6840
rect 6246 6840 6264 6858
rect 6246 6858 6264 6876
rect 6246 6876 6264 6894
rect 6246 6894 6264 6912
rect 6246 6912 6264 6930
rect 6246 6930 6264 6948
rect 6246 6948 6264 6966
rect 6246 6966 6264 6984
rect 6246 6984 6264 7002
rect 6246 7002 6264 7020
rect 6246 7020 6264 7038
rect 6246 7038 6264 7056
rect 6246 7056 6264 7074
rect 6246 7074 6264 7092
rect 6246 7092 6264 7110
rect 6246 7110 6264 7128
rect 6246 7128 6264 7146
rect 6246 7146 6264 7164
rect 6246 7164 6264 7182
rect 6246 7182 6264 7200
rect 6246 7200 6264 7218
rect 6246 7218 6264 7236
rect 6246 7236 6264 7254
rect 6246 7254 6264 7272
rect 6246 7272 6264 7290
rect 6246 7290 6264 7308
rect 6246 7308 6264 7326
rect 6246 7326 6264 7344
rect 6246 7344 6264 7362
rect 6246 7362 6264 7380
rect 6246 7380 6264 7398
rect 6246 7398 6264 7416
rect 6246 7416 6264 7434
rect 6246 7434 6264 7452
rect 6246 7452 6264 7470
rect 6246 7470 6264 7488
rect 6246 7488 6264 7506
rect 6246 7506 6264 7524
rect 6246 7524 6264 7542
rect 6246 7542 6264 7560
rect 6246 7560 6264 7578
rect 6246 7578 6264 7596
rect 6246 7596 6264 7614
rect 6246 7614 6264 7632
rect 6246 7632 6264 7650
rect 6246 7650 6264 7668
rect 6246 7668 6264 7686
rect 6246 7686 6264 7704
rect 6246 7704 6264 7722
rect 6246 7722 6264 7740
rect 6246 7740 6264 7758
rect 6246 7758 6264 7776
rect 6246 7776 6264 7794
rect 6246 7794 6264 7812
rect 6246 7812 6264 7830
rect 6246 7830 6264 7848
rect 6246 7848 6264 7866
rect 6246 7866 6264 7884
rect 6246 7884 6264 7902
rect 6246 7902 6264 7920
rect 6246 7920 6264 7938
rect 6246 7938 6264 7956
rect 6246 7956 6264 7974
rect 6246 7974 6264 7992
rect 6246 7992 6264 8010
rect 6246 8010 6264 8028
rect 6246 8028 6264 8046
rect 6246 8046 6264 8064
rect 6246 8064 6264 8082
rect 6246 8082 6264 8100
rect 6246 8100 6264 8118
rect 6246 8118 6264 8136
rect 6246 8136 6264 8154
rect 6246 8154 6264 8172
rect 6246 8172 6264 8190
rect 6246 8190 6264 8208
rect 6246 8208 6264 8226
rect 6246 8226 6264 8244
rect 6246 8244 6264 8262
rect 6246 8262 6264 8280
rect 6246 8280 6264 8298
rect 6246 8298 6264 8316
rect 6246 8316 6264 8334
rect 6246 8334 6264 8352
rect 6246 8352 6264 8370
rect 6246 8370 6264 8388
rect 6246 8388 6264 8406
rect 6246 8406 6264 8424
rect 6246 8424 6264 8442
rect 6246 8442 6264 8460
rect 6246 8460 6264 8478
rect 6246 8478 6264 8496
rect 6246 8496 6264 8514
rect 6246 8514 6264 8532
rect 6246 8532 6264 8550
rect 6246 8550 6264 8568
rect 6246 8568 6264 8586
rect 6246 8586 6264 8604
rect 6246 8604 6264 8622
rect 6246 8622 6264 8640
rect 6246 8640 6264 8658
rect 6246 8658 6264 8676
rect 6246 8676 6264 8694
rect 6246 8694 6264 8712
rect 6246 8712 6264 8730
rect 6246 8730 6264 8748
rect 6246 8748 6264 8766
rect 6246 8766 6264 8784
rect 6246 8784 6264 8802
rect 6246 8802 6264 8820
rect 6246 8820 6264 8838
rect 6246 8838 6264 8856
rect 6246 8856 6264 8874
rect 6246 8874 6264 8892
rect 6246 8892 6264 8910
rect 6246 8910 6264 8928
rect 6246 8928 6264 8946
rect 6246 8946 6264 8964
rect 6246 8964 6264 8982
rect 6246 8982 6264 9000
rect 6246 9000 6264 9018
rect 6246 9018 6264 9036
rect 6246 9036 6264 9054
rect 6246 9054 6264 9072
rect 6246 9072 6264 9090
rect 6246 9090 6264 9108
rect 6246 9108 6264 9126
rect 6246 9126 6264 9144
rect 6246 9144 6264 9162
rect 6246 9162 6264 9180
rect 6246 9180 6264 9198
rect 6246 9198 6264 9216
rect 6246 9216 6264 9234
rect 6246 9234 6264 9252
rect 6246 9252 6264 9270
rect 6246 9270 6264 9288
rect 6246 9288 6264 9306
rect 6246 9306 6264 9324
rect 6246 9324 6264 9342
rect 6246 9342 6264 9360
rect 6246 9360 6264 9378
rect 6246 9378 6264 9396
rect 6246 9396 6264 9414
rect 6246 9414 6264 9432
rect 6246 9432 6264 9450
rect 6246 9450 6264 9468
rect 6246 9468 6264 9486
rect 6246 9486 6264 9504
rect 6246 9504 6264 9522
rect 6246 9522 6264 9540
rect 6264 1152 6282 1170
rect 6264 1170 6282 1188
rect 6264 1188 6282 1206
rect 6264 1350 6282 1368
rect 6264 1368 6282 1386
rect 6264 1386 6282 1404
rect 6264 1404 6282 1422
rect 6264 1422 6282 1440
rect 6264 1440 6282 1458
rect 6264 1458 6282 1476
rect 6264 1476 6282 1494
rect 6264 1494 6282 1512
rect 6264 1512 6282 1530
rect 6264 1530 6282 1548
rect 6264 1548 6282 1566
rect 6264 1566 6282 1584
rect 6264 1584 6282 1602
rect 6264 1602 6282 1620
rect 6264 1620 6282 1638
rect 6264 1638 6282 1656
rect 6264 1656 6282 1674
rect 6264 1674 6282 1692
rect 6264 1692 6282 1710
rect 6264 1710 6282 1728
rect 6264 1728 6282 1746
rect 6264 1746 6282 1764
rect 6264 1764 6282 1782
rect 6264 1782 6282 1800
rect 6264 1800 6282 1818
rect 6264 1818 6282 1836
rect 6264 1836 6282 1854
rect 6264 1854 6282 1872
rect 6264 1872 6282 1890
rect 6264 1890 6282 1908
rect 6264 1908 6282 1926
rect 6264 1926 6282 1944
rect 6264 1944 6282 1962
rect 6264 1962 6282 1980
rect 6264 1980 6282 1998
rect 6264 1998 6282 2016
rect 6264 2016 6282 2034
rect 6264 2034 6282 2052
rect 6264 2052 6282 2070
rect 6264 2070 6282 2088
rect 6264 2088 6282 2106
rect 6264 2106 6282 2124
rect 6264 2124 6282 2142
rect 6264 2142 6282 2160
rect 6264 2160 6282 2178
rect 6264 2178 6282 2196
rect 6264 2196 6282 2214
rect 6264 2214 6282 2232
rect 6264 2232 6282 2250
rect 6264 2250 6282 2268
rect 6264 2268 6282 2286
rect 6264 2286 6282 2304
rect 6264 2304 6282 2322
rect 6264 2322 6282 2340
rect 6264 2340 6282 2358
rect 6264 2358 6282 2376
rect 6264 2376 6282 2394
rect 6264 2394 6282 2412
rect 6264 2412 6282 2430
rect 6264 2430 6282 2448
rect 6264 2448 6282 2466
rect 6264 2466 6282 2484
rect 6264 2484 6282 2502
rect 6264 2502 6282 2520
rect 6264 2520 6282 2538
rect 6264 2538 6282 2556
rect 6264 2556 6282 2574
rect 6264 2574 6282 2592
rect 6264 2592 6282 2610
rect 6264 2610 6282 2628
rect 6264 2628 6282 2646
rect 6264 2646 6282 2664
rect 6264 2664 6282 2682
rect 6264 2682 6282 2700
rect 6264 2700 6282 2718
rect 6264 2718 6282 2736
rect 6264 2736 6282 2754
rect 6264 2754 6282 2772
rect 6264 2772 6282 2790
rect 6264 2790 6282 2808
rect 6264 2808 6282 2826
rect 6264 2826 6282 2844
rect 6264 3132 6282 3150
rect 6264 3150 6282 3168
rect 6264 3168 6282 3186
rect 6264 3186 6282 3204
rect 6264 3204 6282 3222
rect 6264 3222 6282 3240
rect 6264 3240 6282 3258
rect 6264 3258 6282 3276
rect 6264 3276 6282 3294
rect 6264 3294 6282 3312
rect 6264 3312 6282 3330
rect 6264 3330 6282 3348
rect 6264 3348 6282 3366
rect 6264 3366 6282 3384
rect 6264 3384 6282 3402
rect 6264 3402 6282 3420
rect 6264 3420 6282 3438
rect 6264 3438 6282 3456
rect 6264 3456 6282 3474
rect 6264 3474 6282 3492
rect 6264 3492 6282 3510
rect 6264 3510 6282 3528
rect 6264 3528 6282 3546
rect 6264 3546 6282 3564
rect 6264 3564 6282 3582
rect 6264 3582 6282 3600
rect 6264 3600 6282 3618
rect 6264 3618 6282 3636
rect 6264 3636 6282 3654
rect 6264 3654 6282 3672
rect 6264 3672 6282 3690
rect 6264 3690 6282 3708
rect 6264 3708 6282 3726
rect 6264 3726 6282 3744
rect 6264 3744 6282 3762
rect 6264 3762 6282 3780
rect 6264 3780 6282 3798
rect 6264 3798 6282 3816
rect 6264 3816 6282 3834
rect 6264 3834 6282 3852
rect 6264 3852 6282 3870
rect 6264 3870 6282 3888
rect 6264 3888 6282 3906
rect 6264 3906 6282 3924
rect 6264 3924 6282 3942
rect 6264 3942 6282 3960
rect 6264 3960 6282 3978
rect 6264 3978 6282 3996
rect 6264 3996 6282 4014
rect 6264 4014 6282 4032
rect 6264 4032 6282 4050
rect 6264 4050 6282 4068
rect 6264 4068 6282 4086
rect 6264 4086 6282 4104
rect 6264 4104 6282 4122
rect 6264 4122 6282 4140
rect 6264 4140 6282 4158
rect 6264 4158 6282 4176
rect 6264 4176 6282 4194
rect 6264 4194 6282 4212
rect 6264 4212 6282 4230
rect 6264 4230 6282 4248
rect 6264 4248 6282 4266
rect 6264 4266 6282 4284
rect 6264 4284 6282 4302
rect 6264 4302 6282 4320
rect 6264 4320 6282 4338
rect 6264 4338 6282 4356
rect 6264 4356 6282 4374
rect 6264 4374 6282 4392
rect 6264 4392 6282 4410
rect 6264 4410 6282 4428
rect 6264 4428 6282 4446
rect 6264 4446 6282 4464
rect 6264 4464 6282 4482
rect 6264 4482 6282 4500
rect 6264 4500 6282 4518
rect 6264 4518 6282 4536
rect 6264 4536 6282 4554
rect 6264 4554 6282 4572
rect 6264 4572 6282 4590
rect 6264 4590 6282 4608
rect 6264 4608 6282 4626
rect 6264 4626 6282 4644
rect 6264 4644 6282 4662
rect 6264 4662 6282 4680
rect 6264 4680 6282 4698
rect 6264 4698 6282 4716
rect 6264 4716 6282 4734
rect 6264 4734 6282 4752
rect 6264 4752 6282 4770
rect 6264 4770 6282 4788
rect 6264 4788 6282 4806
rect 6264 4806 6282 4824
rect 6264 4824 6282 4842
rect 6264 4842 6282 4860
rect 6264 4860 6282 4878
rect 6264 4878 6282 4896
rect 6264 4896 6282 4914
rect 6264 4914 6282 4932
rect 6264 4932 6282 4950
rect 6264 4950 6282 4968
rect 6264 4968 6282 4986
rect 6264 4986 6282 5004
rect 6264 5004 6282 5022
rect 6264 5022 6282 5040
rect 6264 5040 6282 5058
rect 6264 5058 6282 5076
rect 6264 5076 6282 5094
rect 6264 5094 6282 5112
rect 6264 5112 6282 5130
rect 6264 5130 6282 5148
rect 6264 5148 6282 5166
rect 6264 5166 6282 5184
rect 6264 5184 6282 5202
rect 6264 5202 6282 5220
rect 6264 5220 6282 5238
rect 6264 5238 6282 5256
rect 6264 5256 6282 5274
rect 6264 5274 6282 5292
rect 6264 5292 6282 5310
rect 6264 5310 6282 5328
rect 6264 5328 6282 5346
rect 6264 5346 6282 5364
rect 6264 5364 6282 5382
rect 6264 5382 6282 5400
rect 6264 5400 6282 5418
rect 6264 5418 6282 5436
rect 6264 5436 6282 5454
rect 6264 5454 6282 5472
rect 6264 5472 6282 5490
rect 6264 5490 6282 5508
rect 6264 5508 6282 5526
rect 6264 5526 6282 5544
rect 6264 5544 6282 5562
rect 6264 5562 6282 5580
rect 6264 5580 6282 5598
rect 6264 5598 6282 5616
rect 6264 5616 6282 5634
rect 6264 6030 6282 6048
rect 6264 6048 6282 6066
rect 6264 6066 6282 6084
rect 6264 6084 6282 6102
rect 6264 6102 6282 6120
rect 6264 6120 6282 6138
rect 6264 6138 6282 6156
rect 6264 6156 6282 6174
rect 6264 6174 6282 6192
rect 6264 6192 6282 6210
rect 6264 6210 6282 6228
rect 6264 6228 6282 6246
rect 6264 6246 6282 6264
rect 6264 6264 6282 6282
rect 6264 6282 6282 6300
rect 6264 6300 6282 6318
rect 6264 6318 6282 6336
rect 6264 6336 6282 6354
rect 6264 6354 6282 6372
rect 6264 6372 6282 6390
rect 6264 6390 6282 6408
rect 6264 6408 6282 6426
rect 6264 6426 6282 6444
rect 6264 6444 6282 6462
rect 6264 6462 6282 6480
rect 6264 6480 6282 6498
rect 6264 6498 6282 6516
rect 6264 6516 6282 6534
rect 6264 6534 6282 6552
rect 6264 6552 6282 6570
rect 6264 6570 6282 6588
rect 6264 6588 6282 6606
rect 6264 6606 6282 6624
rect 6264 6624 6282 6642
rect 6264 6642 6282 6660
rect 6264 6660 6282 6678
rect 6264 6678 6282 6696
rect 6264 6696 6282 6714
rect 6264 6714 6282 6732
rect 6264 6732 6282 6750
rect 6264 6750 6282 6768
rect 6264 6768 6282 6786
rect 6264 6786 6282 6804
rect 6264 6804 6282 6822
rect 6264 6822 6282 6840
rect 6264 6840 6282 6858
rect 6264 6858 6282 6876
rect 6264 6876 6282 6894
rect 6264 6894 6282 6912
rect 6264 6912 6282 6930
rect 6264 6930 6282 6948
rect 6264 6948 6282 6966
rect 6264 6966 6282 6984
rect 6264 6984 6282 7002
rect 6264 7002 6282 7020
rect 6264 7020 6282 7038
rect 6264 7038 6282 7056
rect 6264 7056 6282 7074
rect 6264 7074 6282 7092
rect 6264 7092 6282 7110
rect 6264 7110 6282 7128
rect 6264 7128 6282 7146
rect 6264 7146 6282 7164
rect 6264 7164 6282 7182
rect 6264 7182 6282 7200
rect 6264 7200 6282 7218
rect 6264 7218 6282 7236
rect 6264 7236 6282 7254
rect 6264 7254 6282 7272
rect 6264 7272 6282 7290
rect 6264 7290 6282 7308
rect 6264 7308 6282 7326
rect 6264 7326 6282 7344
rect 6264 7344 6282 7362
rect 6264 7362 6282 7380
rect 6264 7380 6282 7398
rect 6264 7398 6282 7416
rect 6264 7416 6282 7434
rect 6264 7434 6282 7452
rect 6264 7452 6282 7470
rect 6264 7470 6282 7488
rect 6264 7488 6282 7506
rect 6264 7506 6282 7524
rect 6264 7524 6282 7542
rect 6264 7542 6282 7560
rect 6264 7560 6282 7578
rect 6264 7578 6282 7596
rect 6264 7596 6282 7614
rect 6264 7614 6282 7632
rect 6264 7632 6282 7650
rect 6264 7650 6282 7668
rect 6264 7668 6282 7686
rect 6264 7686 6282 7704
rect 6264 7704 6282 7722
rect 6264 7722 6282 7740
rect 6264 7740 6282 7758
rect 6264 7758 6282 7776
rect 6264 7776 6282 7794
rect 6264 7794 6282 7812
rect 6264 7812 6282 7830
rect 6264 7830 6282 7848
rect 6264 7848 6282 7866
rect 6264 7866 6282 7884
rect 6264 7884 6282 7902
rect 6264 7902 6282 7920
rect 6264 7920 6282 7938
rect 6264 7938 6282 7956
rect 6264 7956 6282 7974
rect 6264 7974 6282 7992
rect 6264 7992 6282 8010
rect 6264 8010 6282 8028
rect 6264 8028 6282 8046
rect 6264 8046 6282 8064
rect 6264 8064 6282 8082
rect 6264 8082 6282 8100
rect 6264 8100 6282 8118
rect 6264 8118 6282 8136
rect 6264 8136 6282 8154
rect 6264 8154 6282 8172
rect 6264 8172 6282 8190
rect 6264 8190 6282 8208
rect 6264 8208 6282 8226
rect 6264 8226 6282 8244
rect 6264 8244 6282 8262
rect 6264 8262 6282 8280
rect 6264 8280 6282 8298
rect 6264 8298 6282 8316
rect 6264 8316 6282 8334
rect 6264 8334 6282 8352
rect 6264 8352 6282 8370
rect 6264 8370 6282 8388
rect 6264 8388 6282 8406
rect 6264 8406 6282 8424
rect 6264 8424 6282 8442
rect 6264 8442 6282 8460
rect 6264 8460 6282 8478
rect 6264 8478 6282 8496
rect 6264 8496 6282 8514
rect 6264 8514 6282 8532
rect 6264 8532 6282 8550
rect 6264 8550 6282 8568
rect 6264 8568 6282 8586
rect 6264 8586 6282 8604
rect 6264 8604 6282 8622
rect 6264 8622 6282 8640
rect 6264 8640 6282 8658
rect 6264 8658 6282 8676
rect 6264 8676 6282 8694
rect 6264 8694 6282 8712
rect 6264 8712 6282 8730
rect 6264 8730 6282 8748
rect 6264 8748 6282 8766
rect 6264 8766 6282 8784
rect 6264 8784 6282 8802
rect 6264 8802 6282 8820
rect 6264 8820 6282 8838
rect 6264 8838 6282 8856
rect 6264 8856 6282 8874
rect 6264 8874 6282 8892
rect 6264 8892 6282 8910
rect 6264 8910 6282 8928
rect 6264 8928 6282 8946
rect 6264 8946 6282 8964
rect 6264 8964 6282 8982
rect 6264 8982 6282 9000
rect 6264 9000 6282 9018
rect 6264 9018 6282 9036
rect 6264 9036 6282 9054
rect 6264 9054 6282 9072
rect 6264 9072 6282 9090
rect 6264 9090 6282 9108
rect 6264 9108 6282 9126
rect 6264 9126 6282 9144
rect 6264 9144 6282 9162
rect 6264 9162 6282 9180
rect 6264 9180 6282 9198
rect 6264 9198 6282 9216
rect 6264 9216 6282 9234
rect 6264 9234 6282 9252
rect 6264 9252 6282 9270
rect 6264 9270 6282 9288
rect 6264 9288 6282 9306
rect 6264 9306 6282 9324
rect 6264 9324 6282 9342
rect 6264 9342 6282 9360
rect 6264 9360 6282 9378
rect 6264 9378 6282 9396
rect 6264 9396 6282 9414
rect 6264 9414 6282 9432
rect 6264 9432 6282 9450
rect 6264 9450 6282 9468
rect 6264 9468 6282 9486
rect 6264 9486 6282 9504
rect 6264 9504 6282 9522
rect 6264 9522 6282 9540
rect 6264 9540 6282 9558
rect 6264 9558 6282 9576
rect 6282 1170 6300 1188
rect 6282 1188 6300 1206
rect 6282 1368 6300 1386
rect 6282 1386 6300 1404
rect 6282 1404 6300 1422
rect 6282 1422 6300 1440
rect 6282 1440 6300 1458
rect 6282 1458 6300 1476
rect 6282 1476 6300 1494
rect 6282 1494 6300 1512
rect 6282 1512 6300 1530
rect 6282 1530 6300 1548
rect 6282 1548 6300 1566
rect 6282 1566 6300 1584
rect 6282 1584 6300 1602
rect 6282 1602 6300 1620
rect 6282 1620 6300 1638
rect 6282 1638 6300 1656
rect 6282 1656 6300 1674
rect 6282 1674 6300 1692
rect 6282 1692 6300 1710
rect 6282 1710 6300 1728
rect 6282 1728 6300 1746
rect 6282 1746 6300 1764
rect 6282 1764 6300 1782
rect 6282 1782 6300 1800
rect 6282 1800 6300 1818
rect 6282 1818 6300 1836
rect 6282 1836 6300 1854
rect 6282 1854 6300 1872
rect 6282 1872 6300 1890
rect 6282 1890 6300 1908
rect 6282 1908 6300 1926
rect 6282 1926 6300 1944
rect 6282 1944 6300 1962
rect 6282 1962 6300 1980
rect 6282 1980 6300 1998
rect 6282 1998 6300 2016
rect 6282 2016 6300 2034
rect 6282 2034 6300 2052
rect 6282 2052 6300 2070
rect 6282 2070 6300 2088
rect 6282 2088 6300 2106
rect 6282 2106 6300 2124
rect 6282 2124 6300 2142
rect 6282 2142 6300 2160
rect 6282 2160 6300 2178
rect 6282 2178 6300 2196
rect 6282 2196 6300 2214
rect 6282 2214 6300 2232
rect 6282 2232 6300 2250
rect 6282 2250 6300 2268
rect 6282 2268 6300 2286
rect 6282 2286 6300 2304
rect 6282 2304 6300 2322
rect 6282 2322 6300 2340
rect 6282 2340 6300 2358
rect 6282 2358 6300 2376
rect 6282 2376 6300 2394
rect 6282 2394 6300 2412
rect 6282 2412 6300 2430
rect 6282 2430 6300 2448
rect 6282 2448 6300 2466
rect 6282 2466 6300 2484
rect 6282 2484 6300 2502
rect 6282 2502 6300 2520
rect 6282 2520 6300 2538
rect 6282 2538 6300 2556
rect 6282 2556 6300 2574
rect 6282 2574 6300 2592
rect 6282 2592 6300 2610
rect 6282 2610 6300 2628
rect 6282 2628 6300 2646
rect 6282 2646 6300 2664
rect 6282 2664 6300 2682
rect 6282 2682 6300 2700
rect 6282 2700 6300 2718
rect 6282 2718 6300 2736
rect 6282 2736 6300 2754
rect 6282 2754 6300 2772
rect 6282 2772 6300 2790
rect 6282 2790 6300 2808
rect 6282 2808 6300 2826
rect 6282 2826 6300 2844
rect 6282 2844 6300 2862
rect 6282 3150 6300 3168
rect 6282 3168 6300 3186
rect 6282 3186 6300 3204
rect 6282 3204 6300 3222
rect 6282 3222 6300 3240
rect 6282 3240 6300 3258
rect 6282 3258 6300 3276
rect 6282 3276 6300 3294
rect 6282 3294 6300 3312
rect 6282 3312 6300 3330
rect 6282 3330 6300 3348
rect 6282 3348 6300 3366
rect 6282 3366 6300 3384
rect 6282 3384 6300 3402
rect 6282 3402 6300 3420
rect 6282 3420 6300 3438
rect 6282 3438 6300 3456
rect 6282 3456 6300 3474
rect 6282 3474 6300 3492
rect 6282 3492 6300 3510
rect 6282 3510 6300 3528
rect 6282 3528 6300 3546
rect 6282 3546 6300 3564
rect 6282 3564 6300 3582
rect 6282 3582 6300 3600
rect 6282 3600 6300 3618
rect 6282 3618 6300 3636
rect 6282 3636 6300 3654
rect 6282 3654 6300 3672
rect 6282 3672 6300 3690
rect 6282 3690 6300 3708
rect 6282 3708 6300 3726
rect 6282 3726 6300 3744
rect 6282 3744 6300 3762
rect 6282 3762 6300 3780
rect 6282 3780 6300 3798
rect 6282 3798 6300 3816
rect 6282 3816 6300 3834
rect 6282 3834 6300 3852
rect 6282 3852 6300 3870
rect 6282 3870 6300 3888
rect 6282 3888 6300 3906
rect 6282 3906 6300 3924
rect 6282 3924 6300 3942
rect 6282 3942 6300 3960
rect 6282 3960 6300 3978
rect 6282 3978 6300 3996
rect 6282 3996 6300 4014
rect 6282 4014 6300 4032
rect 6282 4032 6300 4050
rect 6282 4050 6300 4068
rect 6282 4068 6300 4086
rect 6282 4086 6300 4104
rect 6282 4104 6300 4122
rect 6282 4122 6300 4140
rect 6282 4140 6300 4158
rect 6282 4158 6300 4176
rect 6282 4176 6300 4194
rect 6282 4194 6300 4212
rect 6282 4212 6300 4230
rect 6282 4230 6300 4248
rect 6282 4248 6300 4266
rect 6282 4266 6300 4284
rect 6282 4284 6300 4302
rect 6282 4302 6300 4320
rect 6282 4320 6300 4338
rect 6282 4338 6300 4356
rect 6282 4356 6300 4374
rect 6282 4374 6300 4392
rect 6282 4392 6300 4410
rect 6282 4410 6300 4428
rect 6282 4428 6300 4446
rect 6282 4446 6300 4464
rect 6282 4464 6300 4482
rect 6282 4482 6300 4500
rect 6282 4500 6300 4518
rect 6282 4518 6300 4536
rect 6282 4536 6300 4554
rect 6282 4554 6300 4572
rect 6282 4572 6300 4590
rect 6282 4590 6300 4608
rect 6282 4608 6300 4626
rect 6282 4626 6300 4644
rect 6282 4644 6300 4662
rect 6282 4662 6300 4680
rect 6282 4680 6300 4698
rect 6282 4698 6300 4716
rect 6282 4716 6300 4734
rect 6282 4734 6300 4752
rect 6282 4752 6300 4770
rect 6282 4770 6300 4788
rect 6282 4788 6300 4806
rect 6282 4806 6300 4824
rect 6282 4824 6300 4842
rect 6282 4842 6300 4860
rect 6282 4860 6300 4878
rect 6282 4878 6300 4896
rect 6282 4896 6300 4914
rect 6282 4914 6300 4932
rect 6282 4932 6300 4950
rect 6282 4950 6300 4968
rect 6282 4968 6300 4986
rect 6282 4986 6300 5004
rect 6282 5004 6300 5022
rect 6282 5022 6300 5040
rect 6282 5040 6300 5058
rect 6282 5058 6300 5076
rect 6282 5076 6300 5094
rect 6282 5094 6300 5112
rect 6282 5112 6300 5130
rect 6282 5130 6300 5148
rect 6282 5148 6300 5166
rect 6282 5166 6300 5184
rect 6282 5184 6300 5202
rect 6282 5202 6300 5220
rect 6282 5220 6300 5238
rect 6282 5238 6300 5256
rect 6282 5256 6300 5274
rect 6282 5274 6300 5292
rect 6282 5292 6300 5310
rect 6282 5310 6300 5328
rect 6282 5328 6300 5346
rect 6282 5346 6300 5364
rect 6282 5364 6300 5382
rect 6282 5382 6300 5400
rect 6282 5400 6300 5418
rect 6282 5418 6300 5436
rect 6282 5436 6300 5454
rect 6282 5454 6300 5472
rect 6282 5472 6300 5490
rect 6282 5490 6300 5508
rect 6282 5508 6300 5526
rect 6282 5526 6300 5544
rect 6282 5544 6300 5562
rect 6282 5562 6300 5580
rect 6282 5580 6300 5598
rect 6282 5598 6300 5616
rect 6282 5616 6300 5634
rect 6282 5634 6300 5652
rect 6282 6084 6300 6102
rect 6282 6102 6300 6120
rect 6282 6120 6300 6138
rect 6282 6138 6300 6156
rect 6282 6156 6300 6174
rect 6282 6174 6300 6192
rect 6282 6192 6300 6210
rect 6282 6210 6300 6228
rect 6282 6228 6300 6246
rect 6282 6246 6300 6264
rect 6282 6264 6300 6282
rect 6282 6282 6300 6300
rect 6282 6300 6300 6318
rect 6282 6318 6300 6336
rect 6282 6336 6300 6354
rect 6282 6354 6300 6372
rect 6282 6372 6300 6390
rect 6282 6390 6300 6408
rect 6282 6408 6300 6426
rect 6282 6426 6300 6444
rect 6282 6444 6300 6462
rect 6282 6462 6300 6480
rect 6282 6480 6300 6498
rect 6282 6498 6300 6516
rect 6282 6516 6300 6534
rect 6282 6534 6300 6552
rect 6282 6552 6300 6570
rect 6282 6570 6300 6588
rect 6282 6588 6300 6606
rect 6282 6606 6300 6624
rect 6282 6624 6300 6642
rect 6282 6642 6300 6660
rect 6282 6660 6300 6678
rect 6282 6678 6300 6696
rect 6282 6696 6300 6714
rect 6282 6714 6300 6732
rect 6282 6732 6300 6750
rect 6282 6750 6300 6768
rect 6282 6768 6300 6786
rect 6282 6786 6300 6804
rect 6282 6804 6300 6822
rect 6282 6822 6300 6840
rect 6282 6840 6300 6858
rect 6282 6858 6300 6876
rect 6282 6876 6300 6894
rect 6282 6894 6300 6912
rect 6282 6912 6300 6930
rect 6282 6930 6300 6948
rect 6282 6948 6300 6966
rect 6282 6966 6300 6984
rect 6282 6984 6300 7002
rect 6282 7002 6300 7020
rect 6282 7020 6300 7038
rect 6282 7038 6300 7056
rect 6282 7056 6300 7074
rect 6282 7074 6300 7092
rect 6282 7092 6300 7110
rect 6282 7110 6300 7128
rect 6282 7128 6300 7146
rect 6282 7146 6300 7164
rect 6282 7164 6300 7182
rect 6282 7182 6300 7200
rect 6282 7200 6300 7218
rect 6282 7218 6300 7236
rect 6282 7236 6300 7254
rect 6282 7254 6300 7272
rect 6282 7272 6300 7290
rect 6282 7290 6300 7308
rect 6282 7308 6300 7326
rect 6282 7326 6300 7344
rect 6282 7344 6300 7362
rect 6282 7362 6300 7380
rect 6282 7380 6300 7398
rect 6282 7398 6300 7416
rect 6282 7416 6300 7434
rect 6282 7434 6300 7452
rect 6282 7452 6300 7470
rect 6282 7470 6300 7488
rect 6282 7488 6300 7506
rect 6282 7506 6300 7524
rect 6282 7524 6300 7542
rect 6282 7542 6300 7560
rect 6282 7560 6300 7578
rect 6282 7578 6300 7596
rect 6282 7596 6300 7614
rect 6282 7614 6300 7632
rect 6282 7632 6300 7650
rect 6282 7650 6300 7668
rect 6282 7668 6300 7686
rect 6282 7686 6300 7704
rect 6282 7704 6300 7722
rect 6282 7722 6300 7740
rect 6282 7740 6300 7758
rect 6282 7758 6300 7776
rect 6282 7776 6300 7794
rect 6282 7794 6300 7812
rect 6282 7812 6300 7830
rect 6282 7830 6300 7848
rect 6282 7848 6300 7866
rect 6282 7866 6300 7884
rect 6282 7884 6300 7902
rect 6282 7902 6300 7920
rect 6282 7920 6300 7938
rect 6282 7938 6300 7956
rect 6282 7956 6300 7974
rect 6282 7974 6300 7992
rect 6282 7992 6300 8010
rect 6282 8010 6300 8028
rect 6282 8028 6300 8046
rect 6282 8046 6300 8064
rect 6282 8064 6300 8082
rect 6282 8082 6300 8100
rect 6282 8100 6300 8118
rect 6282 8118 6300 8136
rect 6282 8136 6300 8154
rect 6282 8154 6300 8172
rect 6282 8172 6300 8190
rect 6282 8190 6300 8208
rect 6282 8208 6300 8226
rect 6282 8226 6300 8244
rect 6282 8244 6300 8262
rect 6282 8262 6300 8280
rect 6282 8280 6300 8298
rect 6282 8298 6300 8316
rect 6282 8316 6300 8334
rect 6282 8334 6300 8352
rect 6282 8352 6300 8370
rect 6282 8370 6300 8388
rect 6282 8388 6300 8406
rect 6282 8406 6300 8424
rect 6282 8424 6300 8442
rect 6282 8442 6300 8460
rect 6282 8460 6300 8478
rect 6282 8478 6300 8496
rect 6282 8496 6300 8514
rect 6282 8514 6300 8532
rect 6282 8532 6300 8550
rect 6282 8550 6300 8568
rect 6282 8568 6300 8586
rect 6282 8586 6300 8604
rect 6282 8604 6300 8622
rect 6282 8622 6300 8640
rect 6282 8640 6300 8658
rect 6282 8658 6300 8676
rect 6282 8676 6300 8694
rect 6282 8694 6300 8712
rect 6282 8712 6300 8730
rect 6282 8730 6300 8748
rect 6282 8748 6300 8766
rect 6282 8766 6300 8784
rect 6282 8784 6300 8802
rect 6282 8802 6300 8820
rect 6282 8820 6300 8838
rect 6282 8838 6300 8856
rect 6282 8856 6300 8874
rect 6282 8874 6300 8892
rect 6282 8892 6300 8910
rect 6282 8910 6300 8928
rect 6282 8928 6300 8946
rect 6282 8946 6300 8964
rect 6282 8964 6300 8982
rect 6282 8982 6300 9000
rect 6282 9000 6300 9018
rect 6282 9018 6300 9036
rect 6282 9036 6300 9054
rect 6282 9054 6300 9072
rect 6282 9072 6300 9090
rect 6282 9090 6300 9108
rect 6282 9108 6300 9126
rect 6282 9126 6300 9144
rect 6282 9144 6300 9162
rect 6282 9162 6300 9180
rect 6282 9180 6300 9198
rect 6282 9198 6300 9216
rect 6282 9216 6300 9234
rect 6282 9234 6300 9252
rect 6282 9252 6300 9270
rect 6282 9270 6300 9288
rect 6282 9288 6300 9306
rect 6282 9306 6300 9324
rect 6282 9324 6300 9342
rect 6282 9342 6300 9360
rect 6282 9360 6300 9378
rect 6282 9378 6300 9396
rect 6282 9396 6300 9414
rect 6282 9414 6300 9432
rect 6282 9432 6300 9450
rect 6282 9450 6300 9468
rect 6282 9468 6300 9486
rect 6282 9486 6300 9504
rect 6282 9504 6300 9522
rect 6282 9522 6300 9540
rect 6282 9540 6300 9558
rect 6282 9558 6300 9576
rect 6282 9576 6300 9594
rect 6300 1188 6318 1206
rect 6300 1206 6318 1224
rect 6300 1368 6318 1386
rect 6300 1386 6318 1404
rect 6300 1404 6318 1422
rect 6300 1422 6318 1440
rect 6300 1440 6318 1458
rect 6300 1458 6318 1476
rect 6300 1476 6318 1494
rect 6300 1494 6318 1512
rect 6300 1512 6318 1530
rect 6300 1530 6318 1548
rect 6300 1548 6318 1566
rect 6300 1566 6318 1584
rect 6300 1584 6318 1602
rect 6300 1602 6318 1620
rect 6300 1620 6318 1638
rect 6300 1638 6318 1656
rect 6300 1656 6318 1674
rect 6300 1674 6318 1692
rect 6300 1692 6318 1710
rect 6300 1710 6318 1728
rect 6300 1728 6318 1746
rect 6300 1746 6318 1764
rect 6300 1764 6318 1782
rect 6300 1782 6318 1800
rect 6300 1800 6318 1818
rect 6300 1818 6318 1836
rect 6300 1836 6318 1854
rect 6300 1854 6318 1872
rect 6300 1872 6318 1890
rect 6300 1890 6318 1908
rect 6300 1908 6318 1926
rect 6300 1926 6318 1944
rect 6300 1944 6318 1962
rect 6300 1962 6318 1980
rect 6300 1980 6318 1998
rect 6300 1998 6318 2016
rect 6300 2016 6318 2034
rect 6300 2034 6318 2052
rect 6300 2052 6318 2070
rect 6300 2070 6318 2088
rect 6300 2088 6318 2106
rect 6300 2106 6318 2124
rect 6300 2124 6318 2142
rect 6300 2142 6318 2160
rect 6300 2160 6318 2178
rect 6300 2178 6318 2196
rect 6300 2196 6318 2214
rect 6300 2214 6318 2232
rect 6300 2232 6318 2250
rect 6300 2250 6318 2268
rect 6300 2268 6318 2286
rect 6300 2286 6318 2304
rect 6300 2304 6318 2322
rect 6300 2322 6318 2340
rect 6300 2340 6318 2358
rect 6300 2358 6318 2376
rect 6300 2376 6318 2394
rect 6300 2394 6318 2412
rect 6300 2412 6318 2430
rect 6300 2430 6318 2448
rect 6300 2448 6318 2466
rect 6300 2466 6318 2484
rect 6300 2484 6318 2502
rect 6300 2502 6318 2520
rect 6300 2520 6318 2538
rect 6300 2538 6318 2556
rect 6300 2556 6318 2574
rect 6300 2574 6318 2592
rect 6300 2592 6318 2610
rect 6300 2610 6318 2628
rect 6300 2628 6318 2646
rect 6300 2646 6318 2664
rect 6300 2664 6318 2682
rect 6300 2682 6318 2700
rect 6300 2700 6318 2718
rect 6300 2718 6318 2736
rect 6300 2736 6318 2754
rect 6300 2754 6318 2772
rect 6300 2772 6318 2790
rect 6300 2790 6318 2808
rect 6300 2808 6318 2826
rect 6300 2826 6318 2844
rect 6300 2844 6318 2862
rect 6300 3168 6318 3186
rect 6300 3186 6318 3204
rect 6300 3204 6318 3222
rect 6300 3222 6318 3240
rect 6300 3240 6318 3258
rect 6300 3258 6318 3276
rect 6300 3276 6318 3294
rect 6300 3294 6318 3312
rect 6300 3312 6318 3330
rect 6300 3330 6318 3348
rect 6300 3348 6318 3366
rect 6300 3366 6318 3384
rect 6300 3384 6318 3402
rect 6300 3402 6318 3420
rect 6300 3420 6318 3438
rect 6300 3438 6318 3456
rect 6300 3456 6318 3474
rect 6300 3474 6318 3492
rect 6300 3492 6318 3510
rect 6300 3510 6318 3528
rect 6300 3528 6318 3546
rect 6300 3546 6318 3564
rect 6300 3564 6318 3582
rect 6300 3582 6318 3600
rect 6300 3600 6318 3618
rect 6300 3618 6318 3636
rect 6300 3636 6318 3654
rect 6300 3654 6318 3672
rect 6300 3672 6318 3690
rect 6300 3690 6318 3708
rect 6300 3708 6318 3726
rect 6300 3726 6318 3744
rect 6300 3744 6318 3762
rect 6300 3762 6318 3780
rect 6300 3780 6318 3798
rect 6300 3798 6318 3816
rect 6300 3816 6318 3834
rect 6300 3834 6318 3852
rect 6300 3852 6318 3870
rect 6300 3870 6318 3888
rect 6300 3888 6318 3906
rect 6300 3906 6318 3924
rect 6300 3924 6318 3942
rect 6300 3942 6318 3960
rect 6300 3960 6318 3978
rect 6300 3978 6318 3996
rect 6300 3996 6318 4014
rect 6300 4014 6318 4032
rect 6300 4032 6318 4050
rect 6300 4050 6318 4068
rect 6300 4068 6318 4086
rect 6300 4086 6318 4104
rect 6300 4104 6318 4122
rect 6300 4122 6318 4140
rect 6300 4140 6318 4158
rect 6300 4158 6318 4176
rect 6300 4176 6318 4194
rect 6300 4194 6318 4212
rect 6300 4212 6318 4230
rect 6300 4230 6318 4248
rect 6300 4248 6318 4266
rect 6300 4266 6318 4284
rect 6300 4284 6318 4302
rect 6300 4302 6318 4320
rect 6300 4320 6318 4338
rect 6300 4338 6318 4356
rect 6300 4356 6318 4374
rect 6300 4374 6318 4392
rect 6300 4392 6318 4410
rect 6300 4410 6318 4428
rect 6300 4428 6318 4446
rect 6300 4446 6318 4464
rect 6300 4464 6318 4482
rect 6300 4482 6318 4500
rect 6300 4500 6318 4518
rect 6300 4518 6318 4536
rect 6300 4536 6318 4554
rect 6300 4554 6318 4572
rect 6300 4572 6318 4590
rect 6300 4590 6318 4608
rect 6300 4608 6318 4626
rect 6300 4626 6318 4644
rect 6300 4644 6318 4662
rect 6300 4662 6318 4680
rect 6300 4680 6318 4698
rect 6300 4698 6318 4716
rect 6300 4716 6318 4734
rect 6300 4734 6318 4752
rect 6300 4752 6318 4770
rect 6300 4770 6318 4788
rect 6300 4788 6318 4806
rect 6300 4806 6318 4824
rect 6300 4824 6318 4842
rect 6300 4842 6318 4860
rect 6300 4860 6318 4878
rect 6300 4878 6318 4896
rect 6300 4896 6318 4914
rect 6300 4914 6318 4932
rect 6300 4932 6318 4950
rect 6300 4950 6318 4968
rect 6300 4968 6318 4986
rect 6300 4986 6318 5004
rect 6300 5004 6318 5022
rect 6300 5022 6318 5040
rect 6300 5040 6318 5058
rect 6300 5058 6318 5076
rect 6300 5076 6318 5094
rect 6300 5094 6318 5112
rect 6300 5112 6318 5130
rect 6300 5130 6318 5148
rect 6300 5148 6318 5166
rect 6300 5166 6318 5184
rect 6300 5184 6318 5202
rect 6300 5202 6318 5220
rect 6300 5220 6318 5238
rect 6300 5238 6318 5256
rect 6300 5256 6318 5274
rect 6300 5274 6318 5292
rect 6300 5292 6318 5310
rect 6300 5310 6318 5328
rect 6300 5328 6318 5346
rect 6300 5346 6318 5364
rect 6300 5364 6318 5382
rect 6300 5382 6318 5400
rect 6300 5400 6318 5418
rect 6300 5418 6318 5436
rect 6300 5436 6318 5454
rect 6300 5454 6318 5472
rect 6300 5472 6318 5490
rect 6300 5490 6318 5508
rect 6300 5508 6318 5526
rect 6300 5526 6318 5544
rect 6300 5544 6318 5562
rect 6300 5562 6318 5580
rect 6300 5580 6318 5598
rect 6300 5598 6318 5616
rect 6300 5616 6318 5634
rect 6300 5634 6318 5652
rect 6300 6120 6318 6138
rect 6300 6138 6318 6156
rect 6300 6156 6318 6174
rect 6300 6174 6318 6192
rect 6300 6192 6318 6210
rect 6300 6210 6318 6228
rect 6300 6228 6318 6246
rect 6300 6246 6318 6264
rect 6300 6264 6318 6282
rect 6300 6282 6318 6300
rect 6300 6300 6318 6318
rect 6300 6318 6318 6336
rect 6300 6336 6318 6354
rect 6300 6354 6318 6372
rect 6300 6372 6318 6390
rect 6300 6390 6318 6408
rect 6300 6408 6318 6426
rect 6300 6426 6318 6444
rect 6300 6444 6318 6462
rect 6300 6462 6318 6480
rect 6300 6480 6318 6498
rect 6300 6498 6318 6516
rect 6300 6516 6318 6534
rect 6300 6534 6318 6552
rect 6300 6552 6318 6570
rect 6300 6570 6318 6588
rect 6300 6588 6318 6606
rect 6300 6606 6318 6624
rect 6300 6624 6318 6642
rect 6300 6642 6318 6660
rect 6300 6660 6318 6678
rect 6300 6678 6318 6696
rect 6300 6696 6318 6714
rect 6300 6714 6318 6732
rect 6300 6732 6318 6750
rect 6300 6750 6318 6768
rect 6300 6768 6318 6786
rect 6300 6786 6318 6804
rect 6300 6804 6318 6822
rect 6300 6822 6318 6840
rect 6300 6840 6318 6858
rect 6300 6858 6318 6876
rect 6300 6876 6318 6894
rect 6300 6894 6318 6912
rect 6300 6912 6318 6930
rect 6300 6930 6318 6948
rect 6300 6948 6318 6966
rect 6300 6966 6318 6984
rect 6300 6984 6318 7002
rect 6300 7002 6318 7020
rect 6300 7020 6318 7038
rect 6300 7038 6318 7056
rect 6300 7056 6318 7074
rect 6300 7074 6318 7092
rect 6300 7092 6318 7110
rect 6300 7110 6318 7128
rect 6300 7128 6318 7146
rect 6300 7146 6318 7164
rect 6300 7164 6318 7182
rect 6300 7182 6318 7200
rect 6300 7200 6318 7218
rect 6300 7218 6318 7236
rect 6300 7236 6318 7254
rect 6300 7254 6318 7272
rect 6300 7272 6318 7290
rect 6300 7290 6318 7308
rect 6300 7308 6318 7326
rect 6300 7326 6318 7344
rect 6300 7344 6318 7362
rect 6300 7362 6318 7380
rect 6300 7380 6318 7398
rect 6300 7398 6318 7416
rect 6300 7416 6318 7434
rect 6300 7434 6318 7452
rect 6300 7452 6318 7470
rect 6300 7470 6318 7488
rect 6300 7488 6318 7506
rect 6300 7506 6318 7524
rect 6300 7524 6318 7542
rect 6300 7542 6318 7560
rect 6300 7560 6318 7578
rect 6300 7578 6318 7596
rect 6300 7596 6318 7614
rect 6300 7614 6318 7632
rect 6300 7632 6318 7650
rect 6300 7650 6318 7668
rect 6300 7668 6318 7686
rect 6300 7686 6318 7704
rect 6300 7704 6318 7722
rect 6300 7722 6318 7740
rect 6300 7740 6318 7758
rect 6300 7758 6318 7776
rect 6300 7776 6318 7794
rect 6300 7794 6318 7812
rect 6300 7812 6318 7830
rect 6300 7830 6318 7848
rect 6300 7848 6318 7866
rect 6300 7866 6318 7884
rect 6300 7884 6318 7902
rect 6300 7902 6318 7920
rect 6300 7920 6318 7938
rect 6300 7938 6318 7956
rect 6300 7956 6318 7974
rect 6300 7974 6318 7992
rect 6300 7992 6318 8010
rect 6300 8010 6318 8028
rect 6300 8028 6318 8046
rect 6300 8046 6318 8064
rect 6300 8064 6318 8082
rect 6300 8082 6318 8100
rect 6300 8100 6318 8118
rect 6300 8118 6318 8136
rect 6300 8136 6318 8154
rect 6300 8154 6318 8172
rect 6300 8172 6318 8190
rect 6300 8190 6318 8208
rect 6300 8208 6318 8226
rect 6300 8226 6318 8244
rect 6300 8244 6318 8262
rect 6300 8262 6318 8280
rect 6300 8280 6318 8298
rect 6300 8298 6318 8316
rect 6300 8316 6318 8334
rect 6300 8334 6318 8352
rect 6300 8352 6318 8370
rect 6300 8370 6318 8388
rect 6300 8388 6318 8406
rect 6300 8406 6318 8424
rect 6300 8424 6318 8442
rect 6300 8442 6318 8460
rect 6300 8460 6318 8478
rect 6300 8478 6318 8496
rect 6300 8496 6318 8514
rect 6300 8514 6318 8532
rect 6300 8532 6318 8550
rect 6300 8550 6318 8568
rect 6300 8568 6318 8586
rect 6300 8586 6318 8604
rect 6300 8604 6318 8622
rect 6300 8622 6318 8640
rect 6300 8640 6318 8658
rect 6300 8658 6318 8676
rect 6300 8676 6318 8694
rect 6300 8694 6318 8712
rect 6300 8712 6318 8730
rect 6300 8730 6318 8748
rect 6300 8748 6318 8766
rect 6300 8766 6318 8784
rect 6300 8784 6318 8802
rect 6300 8802 6318 8820
rect 6300 8820 6318 8838
rect 6300 8838 6318 8856
rect 6300 8856 6318 8874
rect 6300 8874 6318 8892
rect 6300 8892 6318 8910
rect 6300 8910 6318 8928
rect 6300 8928 6318 8946
rect 6300 8946 6318 8964
rect 6300 8964 6318 8982
rect 6300 8982 6318 9000
rect 6300 9000 6318 9018
rect 6300 9018 6318 9036
rect 6300 9036 6318 9054
rect 6300 9054 6318 9072
rect 6300 9072 6318 9090
rect 6300 9090 6318 9108
rect 6300 9108 6318 9126
rect 6300 9126 6318 9144
rect 6300 9144 6318 9162
rect 6300 9162 6318 9180
rect 6300 9180 6318 9198
rect 6300 9198 6318 9216
rect 6300 9216 6318 9234
rect 6300 9234 6318 9252
rect 6300 9252 6318 9270
rect 6300 9270 6318 9288
rect 6300 9288 6318 9306
rect 6300 9306 6318 9324
rect 6300 9324 6318 9342
rect 6300 9342 6318 9360
rect 6300 9360 6318 9378
rect 6300 9378 6318 9396
rect 6300 9396 6318 9414
rect 6300 9414 6318 9432
rect 6300 9432 6318 9450
rect 6300 9450 6318 9468
rect 6300 9468 6318 9486
rect 6300 9486 6318 9504
rect 6300 9504 6318 9522
rect 6300 9522 6318 9540
rect 6300 9540 6318 9558
rect 6300 9558 6318 9576
rect 6300 9576 6318 9594
rect 6300 9594 6318 9612
rect 6318 1206 6336 1224
rect 6318 1386 6336 1404
rect 6318 1404 6336 1422
rect 6318 1422 6336 1440
rect 6318 1440 6336 1458
rect 6318 1458 6336 1476
rect 6318 1476 6336 1494
rect 6318 1494 6336 1512
rect 6318 1512 6336 1530
rect 6318 1530 6336 1548
rect 6318 1548 6336 1566
rect 6318 1566 6336 1584
rect 6318 1584 6336 1602
rect 6318 1602 6336 1620
rect 6318 1620 6336 1638
rect 6318 1638 6336 1656
rect 6318 1656 6336 1674
rect 6318 1674 6336 1692
rect 6318 1692 6336 1710
rect 6318 1710 6336 1728
rect 6318 1728 6336 1746
rect 6318 1746 6336 1764
rect 6318 1764 6336 1782
rect 6318 1782 6336 1800
rect 6318 1800 6336 1818
rect 6318 1818 6336 1836
rect 6318 1836 6336 1854
rect 6318 1854 6336 1872
rect 6318 1872 6336 1890
rect 6318 1890 6336 1908
rect 6318 1908 6336 1926
rect 6318 1926 6336 1944
rect 6318 1944 6336 1962
rect 6318 1962 6336 1980
rect 6318 1980 6336 1998
rect 6318 1998 6336 2016
rect 6318 2016 6336 2034
rect 6318 2034 6336 2052
rect 6318 2052 6336 2070
rect 6318 2070 6336 2088
rect 6318 2088 6336 2106
rect 6318 2106 6336 2124
rect 6318 2124 6336 2142
rect 6318 2142 6336 2160
rect 6318 2160 6336 2178
rect 6318 2178 6336 2196
rect 6318 2196 6336 2214
rect 6318 2214 6336 2232
rect 6318 2232 6336 2250
rect 6318 2250 6336 2268
rect 6318 2268 6336 2286
rect 6318 2286 6336 2304
rect 6318 2304 6336 2322
rect 6318 2322 6336 2340
rect 6318 2340 6336 2358
rect 6318 2358 6336 2376
rect 6318 2376 6336 2394
rect 6318 2394 6336 2412
rect 6318 2412 6336 2430
rect 6318 2430 6336 2448
rect 6318 2448 6336 2466
rect 6318 2466 6336 2484
rect 6318 2484 6336 2502
rect 6318 2502 6336 2520
rect 6318 2520 6336 2538
rect 6318 2538 6336 2556
rect 6318 2556 6336 2574
rect 6318 2574 6336 2592
rect 6318 2592 6336 2610
rect 6318 2610 6336 2628
rect 6318 2628 6336 2646
rect 6318 2646 6336 2664
rect 6318 2664 6336 2682
rect 6318 2682 6336 2700
rect 6318 2700 6336 2718
rect 6318 2718 6336 2736
rect 6318 2736 6336 2754
rect 6318 2754 6336 2772
rect 6318 2772 6336 2790
rect 6318 2790 6336 2808
rect 6318 2808 6336 2826
rect 6318 2826 6336 2844
rect 6318 2844 6336 2862
rect 6318 2862 6336 2880
rect 6318 3186 6336 3204
rect 6318 3204 6336 3222
rect 6318 3222 6336 3240
rect 6318 3240 6336 3258
rect 6318 3258 6336 3276
rect 6318 3276 6336 3294
rect 6318 3294 6336 3312
rect 6318 3312 6336 3330
rect 6318 3330 6336 3348
rect 6318 3348 6336 3366
rect 6318 3366 6336 3384
rect 6318 3384 6336 3402
rect 6318 3402 6336 3420
rect 6318 3420 6336 3438
rect 6318 3438 6336 3456
rect 6318 3456 6336 3474
rect 6318 3474 6336 3492
rect 6318 3492 6336 3510
rect 6318 3510 6336 3528
rect 6318 3528 6336 3546
rect 6318 3546 6336 3564
rect 6318 3564 6336 3582
rect 6318 3582 6336 3600
rect 6318 3600 6336 3618
rect 6318 3618 6336 3636
rect 6318 3636 6336 3654
rect 6318 3654 6336 3672
rect 6318 3672 6336 3690
rect 6318 3690 6336 3708
rect 6318 3708 6336 3726
rect 6318 3726 6336 3744
rect 6318 3744 6336 3762
rect 6318 3762 6336 3780
rect 6318 3780 6336 3798
rect 6318 3798 6336 3816
rect 6318 3816 6336 3834
rect 6318 3834 6336 3852
rect 6318 3852 6336 3870
rect 6318 3870 6336 3888
rect 6318 3888 6336 3906
rect 6318 3906 6336 3924
rect 6318 3924 6336 3942
rect 6318 3942 6336 3960
rect 6318 3960 6336 3978
rect 6318 3978 6336 3996
rect 6318 3996 6336 4014
rect 6318 4014 6336 4032
rect 6318 4032 6336 4050
rect 6318 4050 6336 4068
rect 6318 4068 6336 4086
rect 6318 4086 6336 4104
rect 6318 4104 6336 4122
rect 6318 4122 6336 4140
rect 6318 4140 6336 4158
rect 6318 4158 6336 4176
rect 6318 4176 6336 4194
rect 6318 4194 6336 4212
rect 6318 4212 6336 4230
rect 6318 4230 6336 4248
rect 6318 4248 6336 4266
rect 6318 4266 6336 4284
rect 6318 4284 6336 4302
rect 6318 4302 6336 4320
rect 6318 4320 6336 4338
rect 6318 4338 6336 4356
rect 6318 4356 6336 4374
rect 6318 4374 6336 4392
rect 6318 4392 6336 4410
rect 6318 4410 6336 4428
rect 6318 4428 6336 4446
rect 6318 4446 6336 4464
rect 6318 4464 6336 4482
rect 6318 4482 6336 4500
rect 6318 4500 6336 4518
rect 6318 4518 6336 4536
rect 6318 4536 6336 4554
rect 6318 4554 6336 4572
rect 6318 4572 6336 4590
rect 6318 4590 6336 4608
rect 6318 4608 6336 4626
rect 6318 4626 6336 4644
rect 6318 4644 6336 4662
rect 6318 4662 6336 4680
rect 6318 4680 6336 4698
rect 6318 4698 6336 4716
rect 6318 4716 6336 4734
rect 6318 4734 6336 4752
rect 6318 4752 6336 4770
rect 6318 4770 6336 4788
rect 6318 4788 6336 4806
rect 6318 4806 6336 4824
rect 6318 4824 6336 4842
rect 6318 4842 6336 4860
rect 6318 4860 6336 4878
rect 6318 4878 6336 4896
rect 6318 4896 6336 4914
rect 6318 4914 6336 4932
rect 6318 4932 6336 4950
rect 6318 4950 6336 4968
rect 6318 4968 6336 4986
rect 6318 4986 6336 5004
rect 6318 5004 6336 5022
rect 6318 5022 6336 5040
rect 6318 5040 6336 5058
rect 6318 5058 6336 5076
rect 6318 5076 6336 5094
rect 6318 5094 6336 5112
rect 6318 5112 6336 5130
rect 6318 5130 6336 5148
rect 6318 5148 6336 5166
rect 6318 5166 6336 5184
rect 6318 5184 6336 5202
rect 6318 5202 6336 5220
rect 6318 5220 6336 5238
rect 6318 5238 6336 5256
rect 6318 5256 6336 5274
rect 6318 5274 6336 5292
rect 6318 5292 6336 5310
rect 6318 5310 6336 5328
rect 6318 5328 6336 5346
rect 6318 5346 6336 5364
rect 6318 5364 6336 5382
rect 6318 5382 6336 5400
rect 6318 5400 6336 5418
rect 6318 5418 6336 5436
rect 6318 5436 6336 5454
rect 6318 5454 6336 5472
rect 6318 5472 6336 5490
rect 6318 5490 6336 5508
rect 6318 5508 6336 5526
rect 6318 5526 6336 5544
rect 6318 5544 6336 5562
rect 6318 5562 6336 5580
rect 6318 5580 6336 5598
rect 6318 5598 6336 5616
rect 6318 5616 6336 5634
rect 6318 5634 6336 5652
rect 6318 5652 6336 5670
rect 6318 6156 6336 6174
rect 6318 6174 6336 6192
rect 6318 6192 6336 6210
rect 6318 6210 6336 6228
rect 6318 6228 6336 6246
rect 6318 6246 6336 6264
rect 6318 6264 6336 6282
rect 6318 6282 6336 6300
rect 6318 6300 6336 6318
rect 6318 6318 6336 6336
rect 6318 6336 6336 6354
rect 6318 6354 6336 6372
rect 6318 6372 6336 6390
rect 6318 6390 6336 6408
rect 6318 6408 6336 6426
rect 6318 6426 6336 6444
rect 6318 6444 6336 6462
rect 6318 6462 6336 6480
rect 6318 6480 6336 6498
rect 6318 6498 6336 6516
rect 6318 6516 6336 6534
rect 6318 6534 6336 6552
rect 6318 6552 6336 6570
rect 6318 6570 6336 6588
rect 6318 6588 6336 6606
rect 6318 6606 6336 6624
rect 6318 6624 6336 6642
rect 6318 6642 6336 6660
rect 6318 6660 6336 6678
rect 6318 6678 6336 6696
rect 6318 6696 6336 6714
rect 6318 6714 6336 6732
rect 6318 6732 6336 6750
rect 6318 6750 6336 6768
rect 6318 6768 6336 6786
rect 6318 6786 6336 6804
rect 6318 6804 6336 6822
rect 6318 6822 6336 6840
rect 6318 6840 6336 6858
rect 6318 6858 6336 6876
rect 6318 6876 6336 6894
rect 6318 6894 6336 6912
rect 6318 6912 6336 6930
rect 6318 6930 6336 6948
rect 6318 6948 6336 6966
rect 6318 6966 6336 6984
rect 6318 6984 6336 7002
rect 6318 7002 6336 7020
rect 6318 7020 6336 7038
rect 6318 7038 6336 7056
rect 6318 7056 6336 7074
rect 6318 7074 6336 7092
rect 6318 7092 6336 7110
rect 6318 7110 6336 7128
rect 6318 7128 6336 7146
rect 6318 7146 6336 7164
rect 6318 7164 6336 7182
rect 6318 7182 6336 7200
rect 6318 7200 6336 7218
rect 6318 7218 6336 7236
rect 6318 7236 6336 7254
rect 6318 7254 6336 7272
rect 6318 7272 6336 7290
rect 6318 7290 6336 7308
rect 6318 7308 6336 7326
rect 6318 7326 6336 7344
rect 6318 7344 6336 7362
rect 6318 7362 6336 7380
rect 6318 7380 6336 7398
rect 6318 7398 6336 7416
rect 6318 7416 6336 7434
rect 6318 7434 6336 7452
rect 6318 7452 6336 7470
rect 6318 7470 6336 7488
rect 6318 7488 6336 7506
rect 6318 7506 6336 7524
rect 6318 7524 6336 7542
rect 6318 7542 6336 7560
rect 6318 7560 6336 7578
rect 6318 7578 6336 7596
rect 6318 7596 6336 7614
rect 6318 7614 6336 7632
rect 6318 7632 6336 7650
rect 6318 7650 6336 7668
rect 6318 7668 6336 7686
rect 6318 7686 6336 7704
rect 6318 7704 6336 7722
rect 6318 7722 6336 7740
rect 6318 7740 6336 7758
rect 6318 7758 6336 7776
rect 6318 7776 6336 7794
rect 6318 7794 6336 7812
rect 6318 7812 6336 7830
rect 6318 7830 6336 7848
rect 6318 7848 6336 7866
rect 6318 7866 6336 7884
rect 6318 7884 6336 7902
rect 6318 7902 6336 7920
rect 6318 7920 6336 7938
rect 6318 7938 6336 7956
rect 6318 7956 6336 7974
rect 6318 7974 6336 7992
rect 6318 7992 6336 8010
rect 6318 8010 6336 8028
rect 6318 8028 6336 8046
rect 6318 8046 6336 8064
rect 6318 8064 6336 8082
rect 6318 8082 6336 8100
rect 6318 8100 6336 8118
rect 6318 8118 6336 8136
rect 6318 8136 6336 8154
rect 6318 8154 6336 8172
rect 6318 8172 6336 8190
rect 6318 8190 6336 8208
rect 6318 8208 6336 8226
rect 6318 8226 6336 8244
rect 6318 8244 6336 8262
rect 6318 8262 6336 8280
rect 6318 8280 6336 8298
rect 6318 8298 6336 8316
rect 6318 8316 6336 8334
rect 6318 8334 6336 8352
rect 6318 8352 6336 8370
rect 6318 8370 6336 8388
rect 6318 8388 6336 8406
rect 6318 8406 6336 8424
rect 6318 8424 6336 8442
rect 6318 8442 6336 8460
rect 6318 8460 6336 8478
rect 6318 8478 6336 8496
rect 6318 8496 6336 8514
rect 6318 8514 6336 8532
rect 6318 8532 6336 8550
rect 6318 8550 6336 8568
rect 6318 8568 6336 8586
rect 6318 8586 6336 8604
rect 6318 8604 6336 8622
rect 6318 8622 6336 8640
rect 6318 8640 6336 8658
rect 6318 8658 6336 8676
rect 6318 8676 6336 8694
rect 6318 8694 6336 8712
rect 6318 8712 6336 8730
rect 6318 8730 6336 8748
rect 6318 8748 6336 8766
rect 6318 8766 6336 8784
rect 6318 8784 6336 8802
rect 6318 8802 6336 8820
rect 6318 8820 6336 8838
rect 6318 8838 6336 8856
rect 6318 8856 6336 8874
rect 6318 8874 6336 8892
rect 6318 8892 6336 8910
rect 6318 8910 6336 8928
rect 6318 8928 6336 8946
rect 6318 8946 6336 8964
rect 6318 8964 6336 8982
rect 6318 8982 6336 9000
rect 6318 9000 6336 9018
rect 6318 9018 6336 9036
rect 6318 9036 6336 9054
rect 6318 9054 6336 9072
rect 6318 9072 6336 9090
rect 6318 9090 6336 9108
rect 6318 9108 6336 9126
rect 6318 9126 6336 9144
rect 6318 9144 6336 9162
rect 6318 9162 6336 9180
rect 6318 9180 6336 9198
rect 6318 9198 6336 9216
rect 6318 9216 6336 9234
rect 6318 9234 6336 9252
rect 6318 9252 6336 9270
rect 6318 9270 6336 9288
rect 6318 9288 6336 9306
rect 6318 9306 6336 9324
rect 6318 9324 6336 9342
rect 6318 9342 6336 9360
rect 6318 9360 6336 9378
rect 6318 9378 6336 9396
rect 6318 9396 6336 9414
rect 6318 9414 6336 9432
rect 6318 9432 6336 9450
rect 6318 9450 6336 9468
rect 6318 9468 6336 9486
rect 6318 9486 6336 9504
rect 6318 9504 6336 9522
rect 6318 9522 6336 9540
rect 6318 9540 6336 9558
rect 6318 9558 6336 9576
rect 6318 9576 6336 9594
rect 6318 9594 6336 9612
rect 6318 9612 6336 9630
rect 6336 1386 6354 1404
rect 6336 1404 6354 1422
rect 6336 1422 6354 1440
rect 6336 1440 6354 1458
rect 6336 1458 6354 1476
rect 6336 1476 6354 1494
rect 6336 1494 6354 1512
rect 6336 1512 6354 1530
rect 6336 1530 6354 1548
rect 6336 1548 6354 1566
rect 6336 1566 6354 1584
rect 6336 1584 6354 1602
rect 6336 1602 6354 1620
rect 6336 1620 6354 1638
rect 6336 1638 6354 1656
rect 6336 1656 6354 1674
rect 6336 1674 6354 1692
rect 6336 1692 6354 1710
rect 6336 1710 6354 1728
rect 6336 1728 6354 1746
rect 6336 1746 6354 1764
rect 6336 1764 6354 1782
rect 6336 1782 6354 1800
rect 6336 1800 6354 1818
rect 6336 1818 6354 1836
rect 6336 1836 6354 1854
rect 6336 1854 6354 1872
rect 6336 1872 6354 1890
rect 6336 1890 6354 1908
rect 6336 1908 6354 1926
rect 6336 1926 6354 1944
rect 6336 1944 6354 1962
rect 6336 1962 6354 1980
rect 6336 1980 6354 1998
rect 6336 1998 6354 2016
rect 6336 2016 6354 2034
rect 6336 2034 6354 2052
rect 6336 2052 6354 2070
rect 6336 2070 6354 2088
rect 6336 2088 6354 2106
rect 6336 2106 6354 2124
rect 6336 2124 6354 2142
rect 6336 2142 6354 2160
rect 6336 2160 6354 2178
rect 6336 2178 6354 2196
rect 6336 2196 6354 2214
rect 6336 2214 6354 2232
rect 6336 2232 6354 2250
rect 6336 2250 6354 2268
rect 6336 2268 6354 2286
rect 6336 2286 6354 2304
rect 6336 2304 6354 2322
rect 6336 2322 6354 2340
rect 6336 2340 6354 2358
rect 6336 2358 6354 2376
rect 6336 2376 6354 2394
rect 6336 2394 6354 2412
rect 6336 2412 6354 2430
rect 6336 2430 6354 2448
rect 6336 2448 6354 2466
rect 6336 2466 6354 2484
rect 6336 2484 6354 2502
rect 6336 2502 6354 2520
rect 6336 2520 6354 2538
rect 6336 2538 6354 2556
rect 6336 2556 6354 2574
rect 6336 2574 6354 2592
rect 6336 2592 6354 2610
rect 6336 2610 6354 2628
rect 6336 2628 6354 2646
rect 6336 2646 6354 2664
rect 6336 2664 6354 2682
rect 6336 2682 6354 2700
rect 6336 2700 6354 2718
rect 6336 2718 6354 2736
rect 6336 2736 6354 2754
rect 6336 2754 6354 2772
rect 6336 2772 6354 2790
rect 6336 2790 6354 2808
rect 6336 2808 6354 2826
rect 6336 2826 6354 2844
rect 6336 2844 6354 2862
rect 6336 2862 6354 2880
rect 6336 3222 6354 3240
rect 6336 3240 6354 3258
rect 6336 3258 6354 3276
rect 6336 3276 6354 3294
rect 6336 3294 6354 3312
rect 6336 3312 6354 3330
rect 6336 3330 6354 3348
rect 6336 3348 6354 3366
rect 6336 3366 6354 3384
rect 6336 3384 6354 3402
rect 6336 3402 6354 3420
rect 6336 3420 6354 3438
rect 6336 3438 6354 3456
rect 6336 3456 6354 3474
rect 6336 3474 6354 3492
rect 6336 3492 6354 3510
rect 6336 3510 6354 3528
rect 6336 3528 6354 3546
rect 6336 3546 6354 3564
rect 6336 3564 6354 3582
rect 6336 3582 6354 3600
rect 6336 3600 6354 3618
rect 6336 3618 6354 3636
rect 6336 3636 6354 3654
rect 6336 3654 6354 3672
rect 6336 3672 6354 3690
rect 6336 3690 6354 3708
rect 6336 3708 6354 3726
rect 6336 3726 6354 3744
rect 6336 3744 6354 3762
rect 6336 3762 6354 3780
rect 6336 3780 6354 3798
rect 6336 3798 6354 3816
rect 6336 3816 6354 3834
rect 6336 3834 6354 3852
rect 6336 3852 6354 3870
rect 6336 3870 6354 3888
rect 6336 3888 6354 3906
rect 6336 3906 6354 3924
rect 6336 3924 6354 3942
rect 6336 3942 6354 3960
rect 6336 3960 6354 3978
rect 6336 3978 6354 3996
rect 6336 3996 6354 4014
rect 6336 4014 6354 4032
rect 6336 4032 6354 4050
rect 6336 4050 6354 4068
rect 6336 4068 6354 4086
rect 6336 4086 6354 4104
rect 6336 4104 6354 4122
rect 6336 4122 6354 4140
rect 6336 4140 6354 4158
rect 6336 4158 6354 4176
rect 6336 4176 6354 4194
rect 6336 4194 6354 4212
rect 6336 4212 6354 4230
rect 6336 4230 6354 4248
rect 6336 4248 6354 4266
rect 6336 4266 6354 4284
rect 6336 4284 6354 4302
rect 6336 4302 6354 4320
rect 6336 4320 6354 4338
rect 6336 4338 6354 4356
rect 6336 4356 6354 4374
rect 6336 4374 6354 4392
rect 6336 4392 6354 4410
rect 6336 4410 6354 4428
rect 6336 4428 6354 4446
rect 6336 4446 6354 4464
rect 6336 4464 6354 4482
rect 6336 4482 6354 4500
rect 6336 4500 6354 4518
rect 6336 4518 6354 4536
rect 6336 4536 6354 4554
rect 6336 4554 6354 4572
rect 6336 4572 6354 4590
rect 6336 4590 6354 4608
rect 6336 4608 6354 4626
rect 6336 4626 6354 4644
rect 6336 4644 6354 4662
rect 6336 4662 6354 4680
rect 6336 4680 6354 4698
rect 6336 4698 6354 4716
rect 6336 4716 6354 4734
rect 6336 4734 6354 4752
rect 6336 4752 6354 4770
rect 6336 4770 6354 4788
rect 6336 4788 6354 4806
rect 6336 4806 6354 4824
rect 6336 4824 6354 4842
rect 6336 4842 6354 4860
rect 6336 4860 6354 4878
rect 6336 4878 6354 4896
rect 6336 4896 6354 4914
rect 6336 4914 6354 4932
rect 6336 4932 6354 4950
rect 6336 4950 6354 4968
rect 6336 4968 6354 4986
rect 6336 4986 6354 5004
rect 6336 5004 6354 5022
rect 6336 5022 6354 5040
rect 6336 5040 6354 5058
rect 6336 5058 6354 5076
rect 6336 5076 6354 5094
rect 6336 5094 6354 5112
rect 6336 5112 6354 5130
rect 6336 5130 6354 5148
rect 6336 5148 6354 5166
rect 6336 5166 6354 5184
rect 6336 5184 6354 5202
rect 6336 5202 6354 5220
rect 6336 5220 6354 5238
rect 6336 5238 6354 5256
rect 6336 5256 6354 5274
rect 6336 5274 6354 5292
rect 6336 5292 6354 5310
rect 6336 5310 6354 5328
rect 6336 5328 6354 5346
rect 6336 5346 6354 5364
rect 6336 5364 6354 5382
rect 6336 5382 6354 5400
rect 6336 5400 6354 5418
rect 6336 5418 6354 5436
rect 6336 5436 6354 5454
rect 6336 5454 6354 5472
rect 6336 5472 6354 5490
rect 6336 5490 6354 5508
rect 6336 5508 6354 5526
rect 6336 5526 6354 5544
rect 6336 5544 6354 5562
rect 6336 5562 6354 5580
rect 6336 5580 6354 5598
rect 6336 5598 6354 5616
rect 6336 5616 6354 5634
rect 6336 5634 6354 5652
rect 6336 5652 6354 5670
rect 6336 5670 6354 5688
rect 6336 6210 6354 6228
rect 6336 6228 6354 6246
rect 6336 6246 6354 6264
rect 6336 6264 6354 6282
rect 6336 6282 6354 6300
rect 6336 6300 6354 6318
rect 6336 6318 6354 6336
rect 6336 6336 6354 6354
rect 6336 6354 6354 6372
rect 6336 6372 6354 6390
rect 6336 6390 6354 6408
rect 6336 6408 6354 6426
rect 6336 6426 6354 6444
rect 6336 6444 6354 6462
rect 6336 6462 6354 6480
rect 6336 6480 6354 6498
rect 6336 6498 6354 6516
rect 6336 6516 6354 6534
rect 6336 6534 6354 6552
rect 6336 6552 6354 6570
rect 6336 6570 6354 6588
rect 6336 6588 6354 6606
rect 6336 6606 6354 6624
rect 6336 6624 6354 6642
rect 6336 6642 6354 6660
rect 6336 6660 6354 6678
rect 6336 6678 6354 6696
rect 6336 6696 6354 6714
rect 6336 6714 6354 6732
rect 6336 6732 6354 6750
rect 6336 6750 6354 6768
rect 6336 6768 6354 6786
rect 6336 6786 6354 6804
rect 6336 6804 6354 6822
rect 6336 6822 6354 6840
rect 6336 6840 6354 6858
rect 6336 6858 6354 6876
rect 6336 6876 6354 6894
rect 6336 6894 6354 6912
rect 6336 6912 6354 6930
rect 6336 6930 6354 6948
rect 6336 6948 6354 6966
rect 6336 6966 6354 6984
rect 6336 6984 6354 7002
rect 6336 7002 6354 7020
rect 6336 7020 6354 7038
rect 6336 7038 6354 7056
rect 6336 7056 6354 7074
rect 6336 7074 6354 7092
rect 6336 7092 6354 7110
rect 6336 7110 6354 7128
rect 6336 7128 6354 7146
rect 6336 7146 6354 7164
rect 6336 7164 6354 7182
rect 6336 7182 6354 7200
rect 6336 7200 6354 7218
rect 6336 7218 6354 7236
rect 6336 7236 6354 7254
rect 6336 7254 6354 7272
rect 6336 7272 6354 7290
rect 6336 7290 6354 7308
rect 6336 7308 6354 7326
rect 6336 7326 6354 7344
rect 6336 7344 6354 7362
rect 6336 7362 6354 7380
rect 6336 7380 6354 7398
rect 6336 7398 6354 7416
rect 6336 7416 6354 7434
rect 6336 7434 6354 7452
rect 6336 7452 6354 7470
rect 6336 7470 6354 7488
rect 6336 7488 6354 7506
rect 6336 7506 6354 7524
rect 6336 7524 6354 7542
rect 6336 7542 6354 7560
rect 6336 7560 6354 7578
rect 6336 7578 6354 7596
rect 6336 7596 6354 7614
rect 6336 7614 6354 7632
rect 6336 7632 6354 7650
rect 6336 7650 6354 7668
rect 6336 7668 6354 7686
rect 6336 7686 6354 7704
rect 6336 7704 6354 7722
rect 6336 7722 6354 7740
rect 6336 7740 6354 7758
rect 6336 7758 6354 7776
rect 6336 7776 6354 7794
rect 6336 7794 6354 7812
rect 6336 7812 6354 7830
rect 6336 7830 6354 7848
rect 6336 7848 6354 7866
rect 6336 7866 6354 7884
rect 6336 7884 6354 7902
rect 6336 7902 6354 7920
rect 6336 7920 6354 7938
rect 6336 7938 6354 7956
rect 6336 7956 6354 7974
rect 6336 7974 6354 7992
rect 6336 7992 6354 8010
rect 6336 8010 6354 8028
rect 6336 8028 6354 8046
rect 6336 8046 6354 8064
rect 6336 8064 6354 8082
rect 6336 8082 6354 8100
rect 6336 8100 6354 8118
rect 6336 8118 6354 8136
rect 6336 8136 6354 8154
rect 6336 8154 6354 8172
rect 6336 8172 6354 8190
rect 6336 8190 6354 8208
rect 6336 8208 6354 8226
rect 6336 8226 6354 8244
rect 6336 8244 6354 8262
rect 6336 8262 6354 8280
rect 6336 8280 6354 8298
rect 6336 8298 6354 8316
rect 6336 8316 6354 8334
rect 6336 8334 6354 8352
rect 6336 8352 6354 8370
rect 6336 8370 6354 8388
rect 6336 8388 6354 8406
rect 6336 8406 6354 8424
rect 6336 8424 6354 8442
rect 6336 8442 6354 8460
rect 6336 8460 6354 8478
rect 6336 8478 6354 8496
rect 6336 8496 6354 8514
rect 6336 8514 6354 8532
rect 6336 8532 6354 8550
rect 6336 8550 6354 8568
rect 6336 8568 6354 8586
rect 6336 8586 6354 8604
rect 6336 8604 6354 8622
rect 6336 8622 6354 8640
rect 6336 8640 6354 8658
rect 6336 8658 6354 8676
rect 6336 8676 6354 8694
rect 6336 8694 6354 8712
rect 6336 8712 6354 8730
rect 6336 8730 6354 8748
rect 6336 8748 6354 8766
rect 6336 8766 6354 8784
rect 6336 8784 6354 8802
rect 6336 8802 6354 8820
rect 6336 8820 6354 8838
rect 6336 8838 6354 8856
rect 6336 8856 6354 8874
rect 6336 8874 6354 8892
rect 6336 8892 6354 8910
rect 6336 8910 6354 8928
rect 6336 8928 6354 8946
rect 6336 8946 6354 8964
rect 6336 8964 6354 8982
rect 6336 8982 6354 9000
rect 6336 9000 6354 9018
rect 6336 9018 6354 9036
rect 6336 9036 6354 9054
rect 6336 9054 6354 9072
rect 6336 9072 6354 9090
rect 6336 9090 6354 9108
rect 6336 9108 6354 9126
rect 6336 9126 6354 9144
rect 6336 9144 6354 9162
rect 6336 9162 6354 9180
rect 6336 9180 6354 9198
rect 6336 9198 6354 9216
rect 6336 9216 6354 9234
rect 6336 9234 6354 9252
rect 6336 9252 6354 9270
rect 6336 9270 6354 9288
rect 6336 9288 6354 9306
rect 6336 9306 6354 9324
rect 6336 9324 6354 9342
rect 6336 9342 6354 9360
rect 6336 9360 6354 9378
rect 6336 9378 6354 9396
rect 6336 9396 6354 9414
rect 6336 9414 6354 9432
rect 6336 9432 6354 9450
rect 6336 9450 6354 9468
rect 6336 9468 6354 9486
rect 6336 9486 6354 9504
rect 6336 9504 6354 9522
rect 6336 9522 6354 9540
rect 6336 9540 6354 9558
rect 6336 9558 6354 9576
rect 6336 9576 6354 9594
rect 6336 9594 6354 9612
rect 6336 9612 6354 9630
rect 6336 9630 6354 9648
rect 6336 9648 6354 9666
rect 6354 1404 6372 1422
rect 6354 1422 6372 1440
rect 6354 1440 6372 1458
rect 6354 1458 6372 1476
rect 6354 1476 6372 1494
rect 6354 1494 6372 1512
rect 6354 1512 6372 1530
rect 6354 1530 6372 1548
rect 6354 1548 6372 1566
rect 6354 1566 6372 1584
rect 6354 1584 6372 1602
rect 6354 1602 6372 1620
rect 6354 1620 6372 1638
rect 6354 1638 6372 1656
rect 6354 1656 6372 1674
rect 6354 1674 6372 1692
rect 6354 1692 6372 1710
rect 6354 1710 6372 1728
rect 6354 1728 6372 1746
rect 6354 1746 6372 1764
rect 6354 1764 6372 1782
rect 6354 1782 6372 1800
rect 6354 1800 6372 1818
rect 6354 1818 6372 1836
rect 6354 1836 6372 1854
rect 6354 1854 6372 1872
rect 6354 1872 6372 1890
rect 6354 1890 6372 1908
rect 6354 1908 6372 1926
rect 6354 1926 6372 1944
rect 6354 1944 6372 1962
rect 6354 1962 6372 1980
rect 6354 1980 6372 1998
rect 6354 1998 6372 2016
rect 6354 2016 6372 2034
rect 6354 2034 6372 2052
rect 6354 2052 6372 2070
rect 6354 2070 6372 2088
rect 6354 2088 6372 2106
rect 6354 2106 6372 2124
rect 6354 2124 6372 2142
rect 6354 2142 6372 2160
rect 6354 2160 6372 2178
rect 6354 2178 6372 2196
rect 6354 2196 6372 2214
rect 6354 2214 6372 2232
rect 6354 2232 6372 2250
rect 6354 2250 6372 2268
rect 6354 2268 6372 2286
rect 6354 2286 6372 2304
rect 6354 2304 6372 2322
rect 6354 2322 6372 2340
rect 6354 2340 6372 2358
rect 6354 2358 6372 2376
rect 6354 2376 6372 2394
rect 6354 2394 6372 2412
rect 6354 2412 6372 2430
rect 6354 2430 6372 2448
rect 6354 2448 6372 2466
rect 6354 2466 6372 2484
rect 6354 2484 6372 2502
rect 6354 2502 6372 2520
rect 6354 2520 6372 2538
rect 6354 2538 6372 2556
rect 6354 2556 6372 2574
rect 6354 2574 6372 2592
rect 6354 2592 6372 2610
rect 6354 2610 6372 2628
rect 6354 2628 6372 2646
rect 6354 2646 6372 2664
rect 6354 2664 6372 2682
rect 6354 2682 6372 2700
rect 6354 2700 6372 2718
rect 6354 2718 6372 2736
rect 6354 2736 6372 2754
rect 6354 2754 6372 2772
rect 6354 2772 6372 2790
rect 6354 2790 6372 2808
rect 6354 2808 6372 2826
rect 6354 2826 6372 2844
rect 6354 2844 6372 2862
rect 6354 2862 6372 2880
rect 6354 3240 6372 3258
rect 6354 3258 6372 3276
rect 6354 3276 6372 3294
rect 6354 3294 6372 3312
rect 6354 3312 6372 3330
rect 6354 3330 6372 3348
rect 6354 3348 6372 3366
rect 6354 3366 6372 3384
rect 6354 3384 6372 3402
rect 6354 3402 6372 3420
rect 6354 3420 6372 3438
rect 6354 3438 6372 3456
rect 6354 3456 6372 3474
rect 6354 3474 6372 3492
rect 6354 3492 6372 3510
rect 6354 3510 6372 3528
rect 6354 3528 6372 3546
rect 6354 3546 6372 3564
rect 6354 3564 6372 3582
rect 6354 3582 6372 3600
rect 6354 3600 6372 3618
rect 6354 3618 6372 3636
rect 6354 3636 6372 3654
rect 6354 3654 6372 3672
rect 6354 3672 6372 3690
rect 6354 3690 6372 3708
rect 6354 3708 6372 3726
rect 6354 3726 6372 3744
rect 6354 3744 6372 3762
rect 6354 3762 6372 3780
rect 6354 3780 6372 3798
rect 6354 3798 6372 3816
rect 6354 3816 6372 3834
rect 6354 3834 6372 3852
rect 6354 3852 6372 3870
rect 6354 3870 6372 3888
rect 6354 3888 6372 3906
rect 6354 3906 6372 3924
rect 6354 3924 6372 3942
rect 6354 3942 6372 3960
rect 6354 3960 6372 3978
rect 6354 3978 6372 3996
rect 6354 3996 6372 4014
rect 6354 4014 6372 4032
rect 6354 4032 6372 4050
rect 6354 4050 6372 4068
rect 6354 4068 6372 4086
rect 6354 4086 6372 4104
rect 6354 4104 6372 4122
rect 6354 4122 6372 4140
rect 6354 4140 6372 4158
rect 6354 4158 6372 4176
rect 6354 4176 6372 4194
rect 6354 4194 6372 4212
rect 6354 4212 6372 4230
rect 6354 4230 6372 4248
rect 6354 4248 6372 4266
rect 6354 4266 6372 4284
rect 6354 4284 6372 4302
rect 6354 4302 6372 4320
rect 6354 4320 6372 4338
rect 6354 4338 6372 4356
rect 6354 4356 6372 4374
rect 6354 4374 6372 4392
rect 6354 4392 6372 4410
rect 6354 4410 6372 4428
rect 6354 4428 6372 4446
rect 6354 4446 6372 4464
rect 6354 4464 6372 4482
rect 6354 4482 6372 4500
rect 6354 4500 6372 4518
rect 6354 4518 6372 4536
rect 6354 4536 6372 4554
rect 6354 4554 6372 4572
rect 6354 4572 6372 4590
rect 6354 4590 6372 4608
rect 6354 4608 6372 4626
rect 6354 4626 6372 4644
rect 6354 4644 6372 4662
rect 6354 4662 6372 4680
rect 6354 4680 6372 4698
rect 6354 4698 6372 4716
rect 6354 4716 6372 4734
rect 6354 4734 6372 4752
rect 6354 4752 6372 4770
rect 6354 4770 6372 4788
rect 6354 4788 6372 4806
rect 6354 4806 6372 4824
rect 6354 4824 6372 4842
rect 6354 4842 6372 4860
rect 6354 4860 6372 4878
rect 6354 4878 6372 4896
rect 6354 4896 6372 4914
rect 6354 4914 6372 4932
rect 6354 4932 6372 4950
rect 6354 4950 6372 4968
rect 6354 4968 6372 4986
rect 6354 4986 6372 5004
rect 6354 5004 6372 5022
rect 6354 5022 6372 5040
rect 6354 5040 6372 5058
rect 6354 5058 6372 5076
rect 6354 5076 6372 5094
rect 6354 5094 6372 5112
rect 6354 5112 6372 5130
rect 6354 5130 6372 5148
rect 6354 5148 6372 5166
rect 6354 5166 6372 5184
rect 6354 5184 6372 5202
rect 6354 5202 6372 5220
rect 6354 5220 6372 5238
rect 6354 5238 6372 5256
rect 6354 5256 6372 5274
rect 6354 5274 6372 5292
rect 6354 5292 6372 5310
rect 6354 5310 6372 5328
rect 6354 5328 6372 5346
rect 6354 5346 6372 5364
rect 6354 5364 6372 5382
rect 6354 5382 6372 5400
rect 6354 5400 6372 5418
rect 6354 5418 6372 5436
rect 6354 5436 6372 5454
rect 6354 5454 6372 5472
rect 6354 5472 6372 5490
rect 6354 5490 6372 5508
rect 6354 5508 6372 5526
rect 6354 5526 6372 5544
rect 6354 5544 6372 5562
rect 6354 5562 6372 5580
rect 6354 5580 6372 5598
rect 6354 5598 6372 5616
rect 6354 5616 6372 5634
rect 6354 5634 6372 5652
rect 6354 5652 6372 5670
rect 6354 5670 6372 5688
rect 6354 5688 6372 5706
rect 6354 6246 6372 6264
rect 6354 6264 6372 6282
rect 6354 6282 6372 6300
rect 6354 6300 6372 6318
rect 6354 6318 6372 6336
rect 6354 6336 6372 6354
rect 6354 6354 6372 6372
rect 6354 6372 6372 6390
rect 6354 6390 6372 6408
rect 6354 6408 6372 6426
rect 6354 6426 6372 6444
rect 6354 6444 6372 6462
rect 6354 6462 6372 6480
rect 6354 6480 6372 6498
rect 6354 6498 6372 6516
rect 6354 6516 6372 6534
rect 6354 6534 6372 6552
rect 6354 6552 6372 6570
rect 6354 6570 6372 6588
rect 6354 6588 6372 6606
rect 6354 6606 6372 6624
rect 6354 6624 6372 6642
rect 6354 6642 6372 6660
rect 6354 6660 6372 6678
rect 6354 6678 6372 6696
rect 6354 6696 6372 6714
rect 6354 6714 6372 6732
rect 6354 6732 6372 6750
rect 6354 6750 6372 6768
rect 6354 6768 6372 6786
rect 6354 6786 6372 6804
rect 6354 6804 6372 6822
rect 6354 6822 6372 6840
rect 6354 6840 6372 6858
rect 6354 6858 6372 6876
rect 6354 6876 6372 6894
rect 6354 6894 6372 6912
rect 6354 6912 6372 6930
rect 6354 6930 6372 6948
rect 6354 6948 6372 6966
rect 6354 6966 6372 6984
rect 6354 6984 6372 7002
rect 6354 7002 6372 7020
rect 6354 7020 6372 7038
rect 6354 7038 6372 7056
rect 6354 7056 6372 7074
rect 6354 7074 6372 7092
rect 6354 7092 6372 7110
rect 6354 7110 6372 7128
rect 6354 7128 6372 7146
rect 6354 7146 6372 7164
rect 6354 7164 6372 7182
rect 6354 7182 6372 7200
rect 6354 7200 6372 7218
rect 6354 7218 6372 7236
rect 6354 7236 6372 7254
rect 6354 7254 6372 7272
rect 6354 7272 6372 7290
rect 6354 7290 6372 7308
rect 6354 7308 6372 7326
rect 6354 7326 6372 7344
rect 6354 7344 6372 7362
rect 6354 7362 6372 7380
rect 6354 7380 6372 7398
rect 6354 7398 6372 7416
rect 6354 7416 6372 7434
rect 6354 7434 6372 7452
rect 6354 7452 6372 7470
rect 6354 7470 6372 7488
rect 6354 7488 6372 7506
rect 6354 7506 6372 7524
rect 6354 7524 6372 7542
rect 6354 7542 6372 7560
rect 6354 7560 6372 7578
rect 6354 7578 6372 7596
rect 6354 7596 6372 7614
rect 6354 7614 6372 7632
rect 6354 7632 6372 7650
rect 6354 7650 6372 7668
rect 6354 7668 6372 7686
rect 6354 7686 6372 7704
rect 6354 7704 6372 7722
rect 6354 7722 6372 7740
rect 6354 7740 6372 7758
rect 6354 7758 6372 7776
rect 6354 7776 6372 7794
rect 6354 7794 6372 7812
rect 6354 7812 6372 7830
rect 6354 7830 6372 7848
rect 6354 7848 6372 7866
rect 6354 7866 6372 7884
rect 6354 7884 6372 7902
rect 6354 7902 6372 7920
rect 6354 7920 6372 7938
rect 6354 7938 6372 7956
rect 6354 7956 6372 7974
rect 6354 7974 6372 7992
rect 6354 7992 6372 8010
rect 6354 8010 6372 8028
rect 6354 8028 6372 8046
rect 6354 8046 6372 8064
rect 6354 8064 6372 8082
rect 6354 8082 6372 8100
rect 6354 8100 6372 8118
rect 6354 8118 6372 8136
rect 6354 8136 6372 8154
rect 6354 8154 6372 8172
rect 6354 8172 6372 8190
rect 6354 8190 6372 8208
rect 6354 8208 6372 8226
rect 6354 8226 6372 8244
rect 6354 8244 6372 8262
rect 6354 8262 6372 8280
rect 6354 8280 6372 8298
rect 6354 8298 6372 8316
rect 6354 8316 6372 8334
rect 6354 8334 6372 8352
rect 6354 8352 6372 8370
rect 6354 8370 6372 8388
rect 6354 8388 6372 8406
rect 6354 8406 6372 8424
rect 6354 8424 6372 8442
rect 6354 8442 6372 8460
rect 6354 8460 6372 8478
rect 6354 8478 6372 8496
rect 6354 8496 6372 8514
rect 6354 8514 6372 8532
rect 6354 8532 6372 8550
rect 6354 8550 6372 8568
rect 6354 8568 6372 8586
rect 6354 8586 6372 8604
rect 6354 8604 6372 8622
rect 6354 8622 6372 8640
rect 6354 8640 6372 8658
rect 6354 8658 6372 8676
rect 6354 8676 6372 8694
rect 6354 8694 6372 8712
rect 6354 8712 6372 8730
rect 6354 8730 6372 8748
rect 6354 8748 6372 8766
rect 6354 8766 6372 8784
rect 6354 8784 6372 8802
rect 6354 8802 6372 8820
rect 6354 8820 6372 8838
rect 6354 8838 6372 8856
rect 6354 8856 6372 8874
rect 6354 8874 6372 8892
rect 6354 8892 6372 8910
rect 6354 8910 6372 8928
rect 6354 8928 6372 8946
rect 6354 8946 6372 8964
rect 6354 8964 6372 8982
rect 6354 8982 6372 9000
rect 6354 9000 6372 9018
rect 6354 9018 6372 9036
rect 6354 9036 6372 9054
rect 6354 9054 6372 9072
rect 6354 9072 6372 9090
rect 6354 9090 6372 9108
rect 6354 9108 6372 9126
rect 6354 9126 6372 9144
rect 6354 9144 6372 9162
rect 6354 9162 6372 9180
rect 6354 9180 6372 9198
rect 6354 9198 6372 9216
rect 6354 9216 6372 9234
rect 6354 9234 6372 9252
rect 6354 9252 6372 9270
rect 6354 9270 6372 9288
rect 6354 9288 6372 9306
rect 6354 9306 6372 9324
rect 6354 9324 6372 9342
rect 6354 9342 6372 9360
rect 6354 9360 6372 9378
rect 6354 9378 6372 9396
rect 6354 9396 6372 9414
rect 6354 9414 6372 9432
rect 6354 9432 6372 9450
rect 6354 9450 6372 9468
rect 6354 9468 6372 9486
rect 6354 9486 6372 9504
rect 6354 9504 6372 9522
rect 6354 9522 6372 9540
rect 6354 9540 6372 9558
rect 6354 9558 6372 9576
rect 6354 9576 6372 9594
rect 6354 9594 6372 9612
rect 6354 9612 6372 9630
rect 6354 9630 6372 9648
rect 6354 9648 6372 9666
rect 6354 9666 6372 9684
rect 6372 1404 6390 1422
rect 6372 1422 6390 1440
rect 6372 1440 6390 1458
rect 6372 1458 6390 1476
rect 6372 1476 6390 1494
rect 6372 1494 6390 1512
rect 6372 1512 6390 1530
rect 6372 1530 6390 1548
rect 6372 1548 6390 1566
rect 6372 1566 6390 1584
rect 6372 1584 6390 1602
rect 6372 1602 6390 1620
rect 6372 1620 6390 1638
rect 6372 1638 6390 1656
rect 6372 1656 6390 1674
rect 6372 1674 6390 1692
rect 6372 1692 6390 1710
rect 6372 1710 6390 1728
rect 6372 1728 6390 1746
rect 6372 1746 6390 1764
rect 6372 1764 6390 1782
rect 6372 1782 6390 1800
rect 6372 1800 6390 1818
rect 6372 1818 6390 1836
rect 6372 1836 6390 1854
rect 6372 1854 6390 1872
rect 6372 1872 6390 1890
rect 6372 1890 6390 1908
rect 6372 1908 6390 1926
rect 6372 1926 6390 1944
rect 6372 1944 6390 1962
rect 6372 1962 6390 1980
rect 6372 1980 6390 1998
rect 6372 1998 6390 2016
rect 6372 2016 6390 2034
rect 6372 2034 6390 2052
rect 6372 2052 6390 2070
rect 6372 2070 6390 2088
rect 6372 2088 6390 2106
rect 6372 2106 6390 2124
rect 6372 2124 6390 2142
rect 6372 2142 6390 2160
rect 6372 2160 6390 2178
rect 6372 2178 6390 2196
rect 6372 2196 6390 2214
rect 6372 2214 6390 2232
rect 6372 2232 6390 2250
rect 6372 2250 6390 2268
rect 6372 2268 6390 2286
rect 6372 2286 6390 2304
rect 6372 2304 6390 2322
rect 6372 2322 6390 2340
rect 6372 2340 6390 2358
rect 6372 2358 6390 2376
rect 6372 2376 6390 2394
rect 6372 2394 6390 2412
rect 6372 2412 6390 2430
rect 6372 2430 6390 2448
rect 6372 2448 6390 2466
rect 6372 2466 6390 2484
rect 6372 2484 6390 2502
rect 6372 2502 6390 2520
rect 6372 2520 6390 2538
rect 6372 2538 6390 2556
rect 6372 2556 6390 2574
rect 6372 2574 6390 2592
rect 6372 2592 6390 2610
rect 6372 2610 6390 2628
rect 6372 2628 6390 2646
rect 6372 2646 6390 2664
rect 6372 2664 6390 2682
rect 6372 2682 6390 2700
rect 6372 2700 6390 2718
rect 6372 2718 6390 2736
rect 6372 2736 6390 2754
rect 6372 2754 6390 2772
rect 6372 2772 6390 2790
rect 6372 2790 6390 2808
rect 6372 2808 6390 2826
rect 6372 2826 6390 2844
rect 6372 2844 6390 2862
rect 6372 2862 6390 2880
rect 6372 2880 6390 2898
rect 6372 3258 6390 3276
rect 6372 3276 6390 3294
rect 6372 3294 6390 3312
rect 6372 3312 6390 3330
rect 6372 3330 6390 3348
rect 6372 3348 6390 3366
rect 6372 3366 6390 3384
rect 6372 3384 6390 3402
rect 6372 3402 6390 3420
rect 6372 3420 6390 3438
rect 6372 3438 6390 3456
rect 6372 3456 6390 3474
rect 6372 3474 6390 3492
rect 6372 3492 6390 3510
rect 6372 3510 6390 3528
rect 6372 3528 6390 3546
rect 6372 3546 6390 3564
rect 6372 3564 6390 3582
rect 6372 3582 6390 3600
rect 6372 3600 6390 3618
rect 6372 3618 6390 3636
rect 6372 3636 6390 3654
rect 6372 3654 6390 3672
rect 6372 3672 6390 3690
rect 6372 3690 6390 3708
rect 6372 3708 6390 3726
rect 6372 3726 6390 3744
rect 6372 3744 6390 3762
rect 6372 3762 6390 3780
rect 6372 3780 6390 3798
rect 6372 3798 6390 3816
rect 6372 3816 6390 3834
rect 6372 3834 6390 3852
rect 6372 3852 6390 3870
rect 6372 3870 6390 3888
rect 6372 3888 6390 3906
rect 6372 3906 6390 3924
rect 6372 3924 6390 3942
rect 6372 3942 6390 3960
rect 6372 3960 6390 3978
rect 6372 3978 6390 3996
rect 6372 3996 6390 4014
rect 6372 4014 6390 4032
rect 6372 4032 6390 4050
rect 6372 4050 6390 4068
rect 6372 4068 6390 4086
rect 6372 4086 6390 4104
rect 6372 4104 6390 4122
rect 6372 4122 6390 4140
rect 6372 4140 6390 4158
rect 6372 4158 6390 4176
rect 6372 4176 6390 4194
rect 6372 4194 6390 4212
rect 6372 4212 6390 4230
rect 6372 4230 6390 4248
rect 6372 4248 6390 4266
rect 6372 4266 6390 4284
rect 6372 4284 6390 4302
rect 6372 4302 6390 4320
rect 6372 4320 6390 4338
rect 6372 4338 6390 4356
rect 6372 4356 6390 4374
rect 6372 4374 6390 4392
rect 6372 4392 6390 4410
rect 6372 4410 6390 4428
rect 6372 4428 6390 4446
rect 6372 4446 6390 4464
rect 6372 4464 6390 4482
rect 6372 4482 6390 4500
rect 6372 4500 6390 4518
rect 6372 4518 6390 4536
rect 6372 4536 6390 4554
rect 6372 4554 6390 4572
rect 6372 4572 6390 4590
rect 6372 4590 6390 4608
rect 6372 4608 6390 4626
rect 6372 4626 6390 4644
rect 6372 4644 6390 4662
rect 6372 4662 6390 4680
rect 6372 4680 6390 4698
rect 6372 4698 6390 4716
rect 6372 4716 6390 4734
rect 6372 4734 6390 4752
rect 6372 4752 6390 4770
rect 6372 4770 6390 4788
rect 6372 4788 6390 4806
rect 6372 4806 6390 4824
rect 6372 4824 6390 4842
rect 6372 4842 6390 4860
rect 6372 4860 6390 4878
rect 6372 4878 6390 4896
rect 6372 4896 6390 4914
rect 6372 4914 6390 4932
rect 6372 4932 6390 4950
rect 6372 4950 6390 4968
rect 6372 4968 6390 4986
rect 6372 4986 6390 5004
rect 6372 5004 6390 5022
rect 6372 5022 6390 5040
rect 6372 5040 6390 5058
rect 6372 5058 6390 5076
rect 6372 5076 6390 5094
rect 6372 5094 6390 5112
rect 6372 5112 6390 5130
rect 6372 5130 6390 5148
rect 6372 5148 6390 5166
rect 6372 5166 6390 5184
rect 6372 5184 6390 5202
rect 6372 5202 6390 5220
rect 6372 5220 6390 5238
rect 6372 5238 6390 5256
rect 6372 5256 6390 5274
rect 6372 5274 6390 5292
rect 6372 5292 6390 5310
rect 6372 5310 6390 5328
rect 6372 5328 6390 5346
rect 6372 5346 6390 5364
rect 6372 5364 6390 5382
rect 6372 5382 6390 5400
rect 6372 5400 6390 5418
rect 6372 5418 6390 5436
rect 6372 5436 6390 5454
rect 6372 5454 6390 5472
rect 6372 5472 6390 5490
rect 6372 5490 6390 5508
rect 6372 5508 6390 5526
rect 6372 5526 6390 5544
rect 6372 5544 6390 5562
rect 6372 5562 6390 5580
rect 6372 5580 6390 5598
rect 6372 5598 6390 5616
rect 6372 5616 6390 5634
rect 6372 5634 6390 5652
rect 6372 5652 6390 5670
rect 6372 5670 6390 5688
rect 6372 5688 6390 5706
rect 6372 5706 6390 5724
rect 6372 6282 6390 6300
rect 6372 6300 6390 6318
rect 6372 6318 6390 6336
rect 6372 6336 6390 6354
rect 6372 6354 6390 6372
rect 6372 6372 6390 6390
rect 6372 6390 6390 6408
rect 6372 6408 6390 6426
rect 6372 6426 6390 6444
rect 6372 6444 6390 6462
rect 6372 6462 6390 6480
rect 6372 6480 6390 6498
rect 6372 6498 6390 6516
rect 6372 6516 6390 6534
rect 6372 6534 6390 6552
rect 6372 6552 6390 6570
rect 6372 6570 6390 6588
rect 6372 6588 6390 6606
rect 6372 6606 6390 6624
rect 6372 6624 6390 6642
rect 6372 6642 6390 6660
rect 6372 6660 6390 6678
rect 6372 6678 6390 6696
rect 6372 6696 6390 6714
rect 6372 6714 6390 6732
rect 6372 6732 6390 6750
rect 6372 6750 6390 6768
rect 6372 6768 6390 6786
rect 6372 6786 6390 6804
rect 6372 6804 6390 6822
rect 6372 6822 6390 6840
rect 6372 6840 6390 6858
rect 6372 6858 6390 6876
rect 6372 6876 6390 6894
rect 6372 6894 6390 6912
rect 6372 6912 6390 6930
rect 6372 6930 6390 6948
rect 6372 6948 6390 6966
rect 6372 6966 6390 6984
rect 6372 6984 6390 7002
rect 6372 7002 6390 7020
rect 6372 7020 6390 7038
rect 6372 7038 6390 7056
rect 6372 7056 6390 7074
rect 6372 7074 6390 7092
rect 6372 7092 6390 7110
rect 6372 7110 6390 7128
rect 6372 7128 6390 7146
rect 6372 7146 6390 7164
rect 6372 7164 6390 7182
rect 6372 7182 6390 7200
rect 6372 7200 6390 7218
rect 6372 7218 6390 7236
rect 6372 7236 6390 7254
rect 6372 7254 6390 7272
rect 6372 7272 6390 7290
rect 6372 7290 6390 7308
rect 6372 7308 6390 7326
rect 6372 7326 6390 7344
rect 6372 7344 6390 7362
rect 6372 7362 6390 7380
rect 6372 7380 6390 7398
rect 6372 7398 6390 7416
rect 6372 7416 6390 7434
rect 6372 7434 6390 7452
rect 6372 7452 6390 7470
rect 6372 7470 6390 7488
rect 6372 7488 6390 7506
rect 6372 7506 6390 7524
rect 6372 7524 6390 7542
rect 6372 7542 6390 7560
rect 6372 7560 6390 7578
rect 6372 7578 6390 7596
rect 6372 7596 6390 7614
rect 6372 7614 6390 7632
rect 6372 7632 6390 7650
rect 6372 7650 6390 7668
rect 6372 7668 6390 7686
rect 6372 7686 6390 7704
rect 6372 7704 6390 7722
rect 6372 7722 6390 7740
rect 6372 7740 6390 7758
rect 6372 7758 6390 7776
rect 6372 7776 6390 7794
rect 6372 7794 6390 7812
rect 6372 7812 6390 7830
rect 6372 7830 6390 7848
rect 6372 7848 6390 7866
rect 6372 7866 6390 7884
rect 6372 7884 6390 7902
rect 6372 7902 6390 7920
rect 6372 7920 6390 7938
rect 6372 7938 6390 7956
rect 6372 7956 6390 7974
rect 6372 7974 6390 7992
rect 6372 7992 6390 8010
rect 6372 8010 6390 8028
rect 6372 8028 6390 8046
rect 6372 8046 6390 8064
rect 6372 8064 6390 8082
rect 6372 8082 6390 8100
rect 6372 8100 6390 8118
rect 6372 8118 6390 8136
rect 6372 8136 6390 8154
rect 6372 8154 6390 8172
rect 6372 8172 6390 8190
rect 6372 8190 6390 8208
rect 6372 8208 6390 8226
rect 6372 8226 6390 8244
rect 6372 8244 6390 8262
rect 6372 8262 6390 8280
rect 6372 8280 6390 8298
rect 6372 8298 6390 8316
rect 6372 8316 6390 8334
rect 6372 8334 6390 8352
rect 6372 8352 6390 8370
rect 6372 8370 6390 8388
rect 6372 8388 6390 8406
rect 6372 8406 6390 8424
rect 6372 8424 6390 8442
rect 6372 8442 6390 8460
rect 6372 8460 6390 8478
rect 6372 8478 6390 8496
rect 6372 8496 6390 8514
rect 6372 8514 6390 8532
rect 6372 8532 6390 8550
rect 6372 8550 6390 8568
rect 6372 8568 6390 8586
rect 6372 8586 6390 8604
rect 6372 8604 6390 8622
rect 6372 8622 6390 8640
rect 6372 8640 6390 8658
rect 6372 8658 6390 8676
rect 6372 8676 6390 8694
rect 6372 8694 6390 8712
rect 6372 8712 6390 8730
rect 6372 8730 6390 8748
rect 6372 8748 6390 8766
rect 6372 8766 6390 8784
rect 6372 8784 6390 8802
rect 6372 8802 6390 8820
rect 6372 8820 6390 8838
rect 6372 8838 6390 8856
rect 6372 8856 6390 8874
rect 6372 8874 6390 8892
rect 6372 8892 6390 8910
rect 6372 8910 6390 8928
rect 6372 8928 6390 8946
rect 6372 8946 6390 8964
rect 6372 8964 6390 8982
rect 6372 8982 6390 9000
rect 6372 9000 6390 9018
rect 6372 9018 6390 9036
rect 6372 9036 6390 9054
rect 6372 9054 6390 9072
rect 6372 9072 6390 9090
rect 6372 9090 6390 9108
rect 6372 9108 6390 9126
rect 6372 9126 6390 9144
rect 6372 9144 6390 9162
rect 6372 9162 6390 9180
rect 6372 9180 6390 9198
rect 6372 9198 6390 9216
rect 6372 9216 6390 9234
rect 6372 9234 6390 9252
rect 6372 9252 6390 9270
rect 6372 9270 6390 9288
rect 6372 9288 6390 9306
rect 6372 9306 6390 9324
rect 6372 9324 6390 9342
rect 6372 9342 6390 9360
rect 6372 9360 6390 9378
rect 6372 9378 6390 9396
rect 6372 9396 6390 9414
rect 6372 9414 6390 9432
rect 6372 9432 6390 9450
rect 6372 9450 6390 9468
rect 6372 9468 6390 9486
rect 6372 9486 6390 9504
rect 6372 9504 6390 9522
rect 6372 9522 6390 9540
rect 6372 9540 6390 9558
rect 6372 9558 6390 9576
rect 6372 9576 6390 9594
rect 6372 9594 6390 9612
rect 6372 9612 6390 9630
rect 6372 9630 6390 9648
rect 6372 9648 6390 9666
rect 6372 9666 6390 9684
rect 6372 9684 6390 9702
rect 6390 1422 6408 1440
rect 6390 1440 6408 1458
rect 6390 1458 6408 1476
rect 6390 1476 6408 1494
rect 6390 1494 6408 1512
rect 6390 1512 6408 1530
rect 6390 1530 6408 1548
rect 6390 1548 6408 1566
rect 6390 1566 6408 1584
rect 6390 1584 6408 1602
rect 6390 1602 6408 1620
rect 6390 1620 6408 1638
rect 6390 1638 6408 1656
rect 6390 1656 6408 1674
rect 6390 1674 6408 1692
rect 6390 1692 6408 1710
rect 6390 1710 6408 1728
rect 6390 1728 6408 1746
rect 6390 1746 6408 1764
rect 6390 1764 6408 1782
rect 6390 1782 6408 1800
rect 6390 1800 6408 1818
rect 6390 1818 6408 1836
rect 6390 1836 6408 1854
rect 6390 1854 6408 1872
rect 6390 1872 6408 1890
rect 6390 1890 6408 1908
rect 6390 1908 6408 1926
rect 6390 1926 6408 1944
rect 6390 1944 6408 1962
rect 6390 1962 6408 1980
rect 6390 1980 6408 1998
rect 6390 1998 6408 2016
rect 6390 2016 6408 2034
rect 6390 2034 6408 2052
rect 6390 2052 6408 2070
rect 6390 2070 6408 2088
rect 6390 2088 6408 2106
rect 6390 2106 6408 2124
rect 6390 2124 6408 2142
rect 6390 2142 6408 2160
rect 6390 2160 6408 2178
rect 6390 2178 6408 2196
rect 6390 2196 6408 2214
rect 6390 2214 6408 2232
rect 6390 2232 6408 2250
rect 6390 2250 6408 2268
rect 6390 2268 6408 2286
rect 6390 2286 6408 2304
rect 6390 2304 6408 2322
rect 6390 2322 6408 2340
rect 6390 2340 6408 2358
rect 6390 2358 6408 2376
rect 6390 2376 6408 2394
rect 6390 2394 6408 2412
rect 6390 2412 6408 2430
rect 6390 2430 6408 2448
rect 6390 2448 6408 2466
rect 6390 2466 6408 2484
rect 6390 2484 6408 2502
rect 6390 2502 6408 2520
rect 6390 2520 6408 2538
rect 6390 2538 6408 2556
rect 6390 2556 6408 2574
rect 6390 2574 6408 2592
rect 6390 2592 6408 2610
rect 6390 2610 6408 2628
rect 6390 2628 6408 2646
rect 6390 2646 6408 2664
rect 6390 2664 6408 2682
rect 6390 2682 6408 2700
rect 6390 2700 6408 2718
rect 6390 2718 6408 2736
rect 6390 2736 6408 2754
rect 6390 2754 6408 2772
rect 6390 2772 6408 2790
rect 6390 2790 6408 2808
rect 6390 2808 6408 2826
rect 6390 2826 6408 2844
rect 6390 2844 6408 2862
rect 6390 2862 6408 2880
rect 6390 2880 6408 2898
rect 6390 3276 6408 3294
rect 6390 3294 6408 3312
rect 6390 3312 6408 3330
rect 6390 3330 6408 3348
rect 6390 3348 6408 3366
rect 6390 3366 6408 3384
rect 6390 3384 6408 3402
rect 6390 3402 6408 3420
rect 6390 3420 6408 3438
rect 6390 3438 6408 3456
rect 6390 3456 6408 3474
rect 6390 3474 6408 3492
rect 6390 3492 6408 3510
rect 6390 3510 6408 3528
rect 6390 3528 6408 3546
rect 6390 3546 6408 3564
rect 6390 3564 6408 3582
rect 6390 3582 6408 3600
rect 6390 3600 6408 3618
rect 6390 3618 6408 3636
rect 6390 3636 6408 3654
rect 6390 3654 6408 3672
rect 6390 3672 6408 3690
rect 6390 3690 6408 3708
rect 6390 3708 6408 3726
rect 6390 3726 6408 3744
rect 6390 3744 6408 3762
rect 6390 3762 6408 3780
rect 6390 3780 6408 3798
rect 6390 3798 6408 3816
rect 6390 3816 6408 3834
rect 6390 3834 6408 3852
rect 6390 3852 6408 3870
rect 6390 3870 6408 3888
rect 6390 3888 6408 3906
rect 6390 3906 6408 3924
rect 6390 3924 6408 3942
rect 6390 3942 6408 3960
rect 6390 3960 6408 3978
rect 6390 3978 6408 3996
rect 6390 3996 6408 4014
rect 6390 4014 6408 4032
rect 6390 4032 6408 4050
rect 6390 4050 6408 4068
rect 6390 4068 6408 4086
rect 6390 4086 6408 4104
rect 6390 4104 6408 4122
rect 6390 4122 6408 4140
rect 6390 4140 6408 4158
rect 6390 4158 6408 4176
rect 6390 4176 6408 4194
rect 6390 4194 6408 4212
rect 6390 4212 6408 4230
rect 6390 4230 6408 4248
rect 6390 4248 6408 4266
rect 6390 4266 6408 4284
rect 6390 4284 6408 4302
rect 6390 4302 6408 4320
rect 6390 4320 6408 4338
rect 6390 4338 6408 4356
rect 6390 4356 6408 4374
rect 6390 4374 6408 4392
rect 6390 4392 6408 4410
rect 6390 4410 6408 4428
rect 6390 4428 6408 4446
rect 6390 4446 6408 4464
rect 6390 4464 6408 4482
rect 6390 4482 6408 4500
rect 6390 4500 6408 4518
rect 6390 4518 6408 4536
rect 6390 4536 6408 4554
rect 6390 4554 6408 4572
rect 6390 4572 6408 4590
rect 6390 4590 6408 4608
rect 6390 4608 6408 4626
rect 6390 4626 6408 4644
rect 6390 4644 6408 4662
rect 6390 4662 6408 4680
rect 6390 4680 6408 4698
rect 6390 4698 6408 4716
rect 6390 4716 6408 4734
rect 6390 4734 6408 4752
rect 6390 4752 6408 4770
rect 6390 4770 6408 4788
rect 6390 4788 6408 4806
rect 6390 4806 6408 4824
rect 6390 4824 6408 4842
rect 6390 4842 6408 4860
rect 6390 4860 6408 4878
rect 6390 4878 6408 4896
rect 6390 4896 6408 4914
rect 6390 4914 6408 4932
rect 6390 4932 6408 4950
rect 6390 4950 6408 4968
rect 6390 4968 6408 4986
rect 6390 4986 6408 5004
rect 6390 5004 6408 5022
rect 6390 5022 6408 5040
rect 6390 5040 6408 5058
rect 6390 5058 6408 5076
rect 6390 5076 6408 5094
rect 6390 5094 6408 5112
rect 6390 5112 6408 5130
rect 6390 5130 6408 5148
rect 6390 5148 6408 5166
rect 6390 5166 6408 5184
rect 6390 5184 6408 5202
rect 6390 5202 6408 5220
rect 6390 5220 6408 5238
rect 6390 5238 6408 5256
rect 6390 5256 6408 5274
rect 6390 5274 6408 5292
rect 6390 5292 6408 5310
rect 6390 5310 6408 5328
rect 6390 5328 6408 5346
rect 6390 5346 6408 5364
rect 6390 5364 6408 5382
rect 6390 5382 6408 5400
rect 6390 5400 6408 5418
rect 6390 5418 6408 5436
rect 6390 5436 6408 5454
rect 6390 5454 6408 5472
rect 6390 5472 6408 5490
rect 6390 5490 6408 5508
rect 6390 5508 6408 5526
rect 6390 5526 6408 5544
rect 6390 5544 6408 5562
rect 6390 5562 6408 5580
rect 6390 5580 6408 5598
rect 6390 5598 6408 5616
rect 6390 5616 6408 5634
rect 6390 5634 6408 5652
rect 6390 5652 6408 5670
rect 6390 5670 6408 5688
rect 6390 5688 6408 5706
rect 6390 5706 6408 5724
rect 6390 5724 6408 5742
rect 6390 6336 6408 6354
rect 6390 6354 6408 6372
rect 6390 6372 6408 6390
rect 6390 6390 6408 6408
rect 6390 6408 6408 6426
rect 6390 6426 6408 6444
rect 6390 6444 6408 6462
rect 6390 6462 6408 6480
rect 6390 6480 6408 6498
rect 6390 6498 6408 6516
rect 6390 6516 6408 6534
rect 6390 6534 6408 6552
rect 6390 6552 6408 6570
rect 6390 6570 6408 6588
rect 6390 6588 6408 6606
rect 6390 6606 6408 6624
rect 6390 6624 6408 6642
rect 6390 6642 6408 6660
rect 6390 6660 6408 6678
rect 6390 6678 6408 6696
rect 6390 6696 6408 6714
rect 6390 6714 6408 6732
rect 6390 6732 6408 6750
rect 6390 6750 6408 6768
rect 6390 6768 6408 6786
rect 6390 6786 6408 6804
rect 6390 6804 6408 6822
rect 6390 6822 6408 6840
rect 6390 6840 6408 6858
rect 6390 6858 6408 6876
rect 6390 6876 6408 6894
rect 6390 6894 6408 6912
rect 6390 6912 6408 6930
rect 6390 6930 6408 6948
rect 6390 6948 6408 6966
rect 6390 6966 6408 6984
rect 6390 6984 6408 7002
rect 6390 7002 6408 7020
rect 6390 7020 6408 7038
rect 6390 7038 6408 7056
rect 6390 7056 6408 7074
rect 6390 7074 6408 7092
rect 6390 7092 6408 7110
rect 6390 7110 6408 7128
rect 6390 7128 6408 7146
rect 6390 7146 6408 7164
rect 6390 7164 6408 7182
rect 6390 7182 6408 7200
rect 6390 7200 6408 7218
rect 6390 7218 6408 7236
rect 6390 7236 6408 7254
rect 6390 7254 6408 7272
rect 6390 7272 6408 7290
rect 6390 7290 6408 7308
rect 6390 7308 6408 7326
rect 6390 7326 6408 7344
rect 6390 7344 6408 7362
rect 6390 7362 6408 7380
rect 6390 7380 6408 7398
rect 6390 7398 6408 7416
rect 6390 7416 6408 7434
rect 6390 7434 6408 7452
rect 6390 7452 6408 7470
rect 6390 7470 6408 7488
rect 6390 7488 6408 7506
rect 6390 7506 6408 7524
rect 6390 7524 6408 7542
rect 6390 7542 6408 7560
rect 6390 7560 6408 7578
rect 6390 7578 6408 7596
rect 6390 7596 6408 7614
rect 6390 7614 6408 7632
rect 6390 7632 6408 7650
rect 6390 7650 6408 7668
rect 6390 7668 6408 7686
rect 6390 7686 6408 7704
rect 6390 7704 6408 7722
rect 6390 7722 6408 7740
rect 6390 7740 6408 7758
rect 6390 7758 6408 7776
rect 6390 7776 6408 7794
rect 6390 7794 6408 7812
rect 6390 7812 6408 7830
rect 6390 7830 6408 7848
rect 6390 7848 6408 7866
rect 6390 7866 6408 7884
rect 6390 7884 6408 7902
rect 6390 7902 6408 7920
rect 6390 7920 6408 7938
rect 6390 7938 6408 7956
rect 6390 7956 6408 7974
rect 6390 7974 6408 7992
rect 6390 7992 6408 8010
rect 6390 8010 6408 8028
rect 6390 8028 6408 8046
rect 6390 8046 6408 8064
rect 6390 8064 6408 8082
rect 6390 8082 6408 8100
rect 6390 8100 6408 8118
rect 6390 8118 6408 8136
rect 6390 8136 6408 8154
rect 6390 8154 6408 8172
rect 6390 8172 6408 8190
rect 6390 8190 6408 8208
rect 6390 8208 6408 8226
rect 6390 8226 6408 8244
rect 6390 8244 6408 8262
rect 6390 8262 6408 8280
rect 6390 8280 6408 8298
rect 6390 8298 6408 8316
rect 6390 8316 6408 8334
rect 6390 8334 6408 8352
rect 6390 8352 6408 8370
rect 6390 8370 6408 8388
rect 6390 8388 6408 8406
rect 6390 8406 6408 8424
rect 6390 8424 6408 8442
rect 6390 8442 6408 8460
rect 6390 8460 6408 8478
rect 6390 8478 6408 8496
rect 6390 8496 6408 8514
rect 6390 8514 6408 8532
rect 6390 8532 6408 8550
rect 6390 8550 6408 8568
rect 6390 8568 6408 8586
rect 6390 8586 6408 8604
rect 6390 8604 6408 8622
rect 6390 8622 6408 8640
rect 6390 8640 6408 8658
rect 6390 8658 6408 8676
rect 6390 8676 6408 8694
rect 6390 8694 6408 8712
rect 6390 8712 6408 8730
rect 6390 8730 6408 8748
rect 6390 8748 6408 8766
rect 6390 8766 6408 8784
rect 6390 8784 6408 8802
rect 6390 8802 6408 8820
rect 6390 8820 6408 8838
rect 6390 8838 6408 8856
rect 6390 8856 6408 8874
rect 6390 8874 6408 8892
rect 6390 8892 6408 8910
rect 6390 8910 6408 8928
rect 6390 8928 6408 8946
rect 6390 8946 6408 8964
rect 6390 8964 6408 8982
rect 6390 8982 6408 9000
rect 6390 9000 6408 9018
rect 6390 9018 6408 9036
rect 6390 9036 6408 9054
rect 6390 9054 6408 9072
rect 6390 9072 6408 9090
rect 6390 9090 6408 9108
rect 6390 9108 6408 9126
rect 6390 9126 6408 9144
rect 6390 9144 6408 9162
rect 6390 9162 6408 9180
rect 6390 9180 6408 9198
rect 6390 9198 6408 9216
rect 6390 9216 6408 9234
rect 6390 9234 6408 9252
rect 6390 9252 6408 9270
rect 6390 9270 6408 9288
rect 6390 9288 6408 9306
rect 6390 9306 6408 9324
rect 6390 9324 6408 9342
rect 6390 9342 6408 9360
rect 6390 9360 6408 9378
rect 6390 9378 6408 9396
rect 6390 9396 6408 9414
rect 6390 9414 6408 9432
rect 6390 9432 6408 9450
rect 6390 9450 6408 9468
rect 6390 9468 6408 9486
rect 6390 9486 6408 9504
rect 6390 9504 6408 9522
rect 6390 9522 6408 9540
rect 6390 9540 6408 9558
rect 6390 9558 6408 9576
rect 6390 9576 6408 9594
rect 6390 9594 6408 9612
rect 6390 9612 6408 9630
rect 6390 9630 6408 9648
rect 6390 9648 6408 9666
rect 6390 9666 6408 9684
rect 6390 9684 6408 9702
rect 6390 9702 6408 9720
rect 6408 1422 6426 1440
rect 6408 1440 6426 1458
rect 6408 1458 6426 1476
rect 6408 1476 6426 1494
rect 6408 1494 6426 1512
rect 6408 1512 6426 1530
rect 6408 1530 6426 1548
rect 6408 1548 6426 1566
rect 6408 1566 6426 1584
rect 6408 1584 6426 1602
rect 6408 1602 6426 1620
rect 6408 1620 6426 1638
rect 6408 1638 6426 1656
rect 6408 1656 6426 1674
rect 6408 1674 6426 1692
rect 6408 1692 6426 1710
rect 6408 1710 6426 1728
rect 6408 1728 6426 1746
rect 6408 1746 6426 1764
rect 6408 1764 6426 1782
rect 6408 1782 6426 1800
rect 6408 1800 6426 1818
rect 6408 1818 6426 1836
rect 6408 1836 6426 1854
rect 6408 1854 6426 1872
rect 6408 1872 6426 1890
rect 6408 1890 6426 1908
rect 6408 1908 6426 1926
rect 6408 1926 6426 1944
rect 6408 1944 6426 1962
rect 6408 1962 6426 1980
rect 6408 1980 6426 1998
rect 6408 1998 6426 2016
rect 6408 2016 6426 2034
rect 6408 2034 6426 2052
rect 6408 2052 6426 2070
rect 6408 2070 6426 2088
rect 6408 2088 6426 2106
rect 6408 2106 6426 2124
rect 6408 2124 6426 2142
rect 6408 2142 6426 2160
rect 6408 2160 6426 2178
rect 6408 2178 6426 2196
rect 6408 2196 6426 2214
rect 6408 2214 6426 2232
rect 6408 2232 6426 2250
rect 6408 2250 6426 2268
rect 6408 2268 6426 2286
rect 6408 2286 6426 2304
rect 6408 2304 6426 2322
rect 6408 2322 6426 2340
rect 6408 2340 6426 2358
rect 6408 2358 6426 2376
rect 6408 2376 6426 2394
rect 6408 2394 6426 2412
rect 6408 2412 6426 2430
rect 6408 2430 6426 2448
rect 6408 2448 6426 2466
rect 6408 2466 6426 2484
rect 6408 2484 6426 2502
rect 6408 2502 6426 2520
rect 6408 2520 6426 2538
rect 6408 2538 6426 2556
rect 6408 2556 6426 2574
rect 6408 2574 6426 2592
rect 6408 2592 6426 2610
rect 6408 2610 6426 2628
rect 6408 2628 6426 2646
rect 6408 2646 6426 2664
rect 6408 2664 6426 2682
rect 6408 2682 6426 2700
rect 6408 2700 6426 2718
rect 6408 2718 6426 2736
rect 6408 2736 6426 2754
rect 6408 2754 6426 2772
rect 6408 2772 6426 2790
rect 6408 2790 6426 2808
rect 6408 2808 6426 2826
rect 6408 2826 6426 2844
rect 6408 2844 6426 2862
rect 6408 2862 6426 2880
rect 6408 2880 6426 2898
rect 6408 3294 6426 3312
rect 6408 3312 6426 3330
rect 6408 3330 6426 3348
rect 6408 3348 6426 3366
rect 6408 3366 6426 3384
rect 6408 3384 6426 3402
rect 6408 3402 6426 3420
rect 6408 3420 6426 3438
rect 6408 3438 6426 3456
rect 6408 3456 6426 3474
rect 6408 3474 6426 3492
rect 6408 3492 6426 3510
rect 6408 3510 6426 3528
rect 6408 3528 6426 3546
rect 6408 3546 6426 3564
rect 6408 3564 6426 3582
rect 6408 3582 6426 3600
rect 6408 3600 6426 3618
rect 6408 3618 6426 3636
rect 6408 3636 6426 3654
rect 6408 3654 6426 3672
rect 6408 3672 6426 3690
rect 6408 3690 6426 3708
rect 6408 3708 6426 3726
rect 6408 3726 6426 3744
rect 6408 3744 6426 3762
rect 6408 3762 6426 3780
rect 6408 3780 6426 3798
rect 6408 3798 6426 3816
rect 6408 3816 6426 3834
rect 6408 3834 6426 3852
rect 6408 3852 6426 3870
rect 6408 3870 6426 3888
rect 6408 3888 6426 3906
rect 6408 3906 6426 3924
rect 6408 3924 6426 3942
rect 6408 3942 6426 3960
rect 6408 3960 6426 3978
rect 6408 3978 6426 3996
rect 6408 3996 6426 4014
rect 6408 4014 6426 4032
rect 6408 4032 6426 4050
rect 6408 4050 6426 4068
rect 6408 4068 6426 4086
rect 6408 4086 6426 4104
rect 6408 4104 6426 4122
rect 6408 4122 6426 4140
rect 6408 4140 6426 4158
rect 6408 4158 6426 4176
rect 6408 4176 6426 4194
rect 6408 4194 6426 4212
rect 6408 4212 6426 4230
rect 6408 4230 6426 4248
rect 6408 4248 6426 4266
rect 6408 4266 6426 4284
rect 6408 4284 6426 4302
rect 6408 4302 6426 4320
rect 6408 4320 6426 4338
rect 6408 4338 6426 4356
rect 6408 4356 6426 4374
rect 6408 4374 6426 4392
rect 6408 4392 6426 4410
rect 6408 4410 6426 4428
rect 6408 4428 6426 4446
rect 6408 4446 6426 4464
rect 6408 4464 6426 4482
rect 6408 4482 6426 4500
rect 6408 4500 6426 4518
rect 6408 4518 6426 4536
rect 6408 4536 6426 4554
rect 6408 4554 6426 4572
rect 6408 4572 6426 4590
rect 6408 4590 6426 4608
rect 6408 4608 6426 4626
rect 6408 4626 6426 4644
rect 6408 4644 6426 4662
rect 6408 4662 6426 4680
rect 6408 4680 6426 4698
rect 6408 4698 6426 4716
rect 6408 4716 6426 4734
rect 6408 4734 6426 4752
rect 6408 4752 6426 4770
rect 6408 4770 6426 4788
rect 6408 4788 6426 4806
rect 6408 4806 6426 4824
rect 6408 4824 6426 4842
rect 6408 4842 6426 4860
rect 6408 4860 6426 4878
rect 6408 4878 6426 4896
rect 6408 4896 6426 4914
rect 6408 4914 6426 4932
rect 6408 4932 6426 4950
rect 6408 4950 6426 4968
rect 6408 4968 6426 4986
rect 6408 4986 6426 5004
rect 6408 5004 6426 5022
rect 6408 5022 6426 5040
rect 6408 5040 6426 5058
rect 6408 5058 6426 5076
rect 6408 5076 6426 5094
rect 6408 5094 6426 5112
rect 6408 5112 6426 5130
rect 6408 5130 6426 5148
rect 6408 5148 6426 5166
rect 6408 5166 6426 5184
rect 6408 5184 6426 5202
rect 6408 5202 6426 5220
rect 6408 5220 6426 5238
rect 6408 5238 6426 5256
rect 6408 5256 6426 5274
rect 6408 5274 6426 5292
rect 6408 5292 6426 5310
rect 6408 5310 6426 5328
rect 6408 5328 6426 5346
rect 6408 5346 6426 5364
rect 6408 5364 6426 5382
rect 6408 5382 6426 5400
rect 6408 5400 6426 5418
rect 6408 5418 6426 5436
rect 6408 5436 6426 5454
rect 6408 5454 6426 5472
rect 6408 5472 6426 5490
rect 6408 5490 6426 5508
rect 6408 5508 6426 5526
rect 6408 5526 6426 5544
rect 6408 5544 6426 5562
rect 6408 5562 6426 5580
rect 6408 5580 6426 5598
rect 6408 5598 6426 5616
rect 6408 5616 6426 5634
rect 6408 5634 6426 5652
rect 6408 5652 6426 5670
rect 6408 5670 6426 5688
rect 6408 5688 6426 5706
rect 6408 5706 6426 5724
rect 6408 5724 6426 5742
rect 6408 5742 6426 5760
rect 6408 6372 6426 6390
rect 6408 6390 6426 6408
rect 6408 6408 6426 6426
rect 6408 6426 6426 6444
rect 6408 6444 6426 6462
rect 6408 6462 6426 6480
rect 6408 6480 6426 6498
rect 6408 6498 6426 6516
rect 6408 6516 6426 6534
rect 6408 6534 6426 6552
rect 6408 6552 6426 6570
rect 6408 6570 6426 6588
rect 6408 6588 6426 6606
rect 6408 6606 6426 6624
rect 6408 6624 6426 6642
rect 6408 6642 6426 6660
rect 6408 6660 6426 6678
rect 6408 6678 6426 6696
rect 6408 6696 6426 6714
rect 6408 6714 6426 6732
rect 6408 6732 6426 6750
rect 6408 6750 6426 6768
rect 6408 6768 6426 6786
rect 6408 6786 6426 6804
rect 6408 6804 6426 6822
rect 6408 6822 6426 6840
rect 6408 6840 6426 6858
rect 6408 6858 6426 6876
rect 6408 6876 6426 6894
rect 6408 6894 6426 6912
rect 6408 6912 6426 6930
rect 6408 6930 6426 6948
rect 6408 6948 6426 6966
rect 6408 6966 6426 6984
rect 6408 6984 6426 7002
rect 6408 7002 6426 7020
rect 6408 7020 6426 7038
rect 6408 7038 6426 7056
rect 6408 7056 6426 7074
rect 6408 7074 6426 7092
rect 6408 7092 6426 7110
rect 6408 7110 6426 7128
rect 6408 7128 6426 7146
rect 6408 7146 6426 7164
rect 6408 7164 6426 7182
rect 6408 7182 6426 7200
rect 6408 7200 6426 7218
rect 6408 7218 6426 7236
rect 6408 7236 6426 7254
rect 6408 7254 6426 7272
rect 6408 7272 6426 7290
rect 6408 7290 6426 7308
rect 6408 7308 6426 7326
rect 6408 7326 6426 7344
rect 6408 7344 6426 7362
rect 6408 7362 6426 7380
rect 6408 7380 6426 7398
rect 6408 7398 6426 7416
rect 6408 7416 6426 7434
rect 6408 7434 6426 7452
rect 6408 7452 6426 7470
rect 6408 7470 6426 7488
rect 6408 7488 6426 7506
rect 6408 7506 6426 7524
rect 6408 7524 6426 7542
rect 6408 7542 6426 7560
rect 6408 7560 6426 7578
rect 6408 7578 6426 7596
rect 6408 7596 6426 7614
rect 6408 7614 6426 7632
rect 6408 7632 6426 7650
rect 6408 7650 6426 7668
rect 6408 7668 6426 7686
rect 6408 7686 6426 7704
rect 6408 7704 6426 7722
rect 6408 7722 6426 7740
rect 6408 7740 6426 7758
rect 6408 7758 6426 7776
rect 6408 7776 6426 7794
rect 6408 7794 6426 7812
rect 6408 7812 6426 7830
rect 6408 7830 6426 7848
rect 6408 7848 6426 7866
rect 6408 7866 6426 7884
rect 6408 7884 6426 7902
rect 6408 7902 6426 7920
rect 6408 7920 6426 7938
rect 6408 7938 6426 7956
rect 6408 7956 6426 7974
rect 6408 7974 6426 7992
rect 6408 7992 6426 8010
rect 6408 8010 6426 8028
rect 6408 8028 6426 8046
rect 6408 8046 6426 8064
rect 6408 8064 6426 8082
rect 6408 8082 6426 8100
rect 6408 8100 6426 8118
rect 6408 8118 6426 8136
rect 6408 8136 6426 8154
rect 6408 8154 6426 8172
rect 6408 8172 6426 8190
rect 6408 8190 6426 8208
rect 6408 8208 6426 8226
rect 6408 8226 6426 8244
rect 6408 8244 6426 8262
rect 6408 8262 6426 8280
rect 6408 8280 6426 8298
rect 6408 8298 6426 8316
rect 6408 8316 6426 8334
rect 6408 8334 6426 8352
rect 6408 8352 6426 8370
rect 6408 8370 6426 8388
rect 6408 8388 6426 8406
rect 6408 8406 6426 8424
rect 6408 8424 6426 8442
rect 6408 8442 6426 8460
rect 6408 8460 6426 8478
rect 6408 8478 6426 8496
rect 6408 8496 6426 8514
rect 6408 8514 6426 8532
rect 6408 8532 6426 8550
rect 6408 8550 6426 8568
rect 6408 8568 6426 8586
rect 6408 8586 6426 8604
rect 6408 8604 6426 8622
rect 6408 8622 6426 8640
rect 6408 8640 6426 8658
rect 6408 8658 6426 8676
rect 6408 8676 6426 8694
rect 6408 8694 6426 8712
rect 6408 8712 6426 8730
rect 6408 8730 6426 8748
rect 6408 8748 6426 8766
rect 6408 8766 6426 8784
rect 6408 8784 6426 8802
rect 6408 8802 6426 8820
rect 6408 8820 6426 8838
rect 6408 8838 6426 8856
rect 6408 8856 6426 8874
rect 6408 8874 6426 8892
rect 6408 8892 6426 8910
rect 6408 8910 6426 8928
rect 6408 8928 6426 8946
rect 6408 8946 6426 8964
rect 6408 8964 6426 8982
rect 6408 8982 6426 9000
rect 6408 9000 6426 9018
rect 6408 9018 6426 9036
rect 6408 9036 6426 9054
rect 6408 9054 6426 9072
rect 6408 9072 6426 9090
rect 6408 9090 6426 9108
rect 6408 9108 6426 9126
rect 6408 9126 6426 9144
rect 6408 9144 6426 9162
rect 6408 9162 6426 9180
rect 6408 9180 6426 9198
rect 6408 9198 6426 9216
rect 6408 9216 6426 9234
rect 6408 9234 6426 9252
rect 6408 9252 6426 9270
rect 6408 9270 6426 9288
rect 6408 9288 6426 9306
rect 6408 9306 6426 9324
rect 6408 9324 6426 9342
rect 6408 9342 6426 9360
rect 6408 9360 6426 9378
rect 6408 9378 6426 9396
rect 6408 9396 6426 9414
rect 6408 9414 6426 9432
rect 6408 9432 6426 9450
rect 6408 9450 6426 9468
rect 6408 9468 6426 9486
rect 6408 9486 6426 9504
rect 6408 9504 6426 9522
rect 6408 9522 6426 9540
rect 6408 9540 6426 9558
rect 6408 9558 6426 9576
rect 6408 9576 6426 9594
rect 6408 9594 6426 9612
rect 6408 9612 6426 9630
rect 6408 9630 6426 9648
rect 6408 9648 6426 9666
rect 6408 9666 6426 9684
rect 6408 9684 6426 9702
rect 6408 9702 6426 9720
rect 6408 9720 6426 9738
rect 6408 9738 6426 9756
rect 6426 1440 6444 1458
rect 6426 1458 6444 1476
rect 6426 1476 6444 1494
rect 6426 1494 6444 1512
rect 6426 1512 6444 1530
rect 6426 1530 6444 1548
rect 6426 1548 6444 1566
rect 6426 1566 6444 1584
rect 6426 1584 6444 1602
rect 6426 1602 6444 1620
rect 6426 1620 6444 1638
rect 6426 1638 6444 1656
rect 6426 1656 6444 1674
rect 6426 1674 6444 1692
rect 6426 1692 6444 1710
rect 6426 1710 6444 1728
rect 6426 1728 6444 1746
rect 6426 1746 6444 1764
rect 6426 1764 6444 1782
rect 6426 1782 6444 1800
rect 6426 1800 6444 1818
rect 6426 1818 6444 1836
rect 6426 1836 6444 1854
rect 6426 1854 6444 1872
rect 6426 1872 6444 1890
rect 6426 1890 6444 1908
rect 6426 1908 6444 1926
rect 6426 1926 6444 1944
rect 6426 1944 6444 1962
rect 6426 1962 6444 1980
rect 6426 1980 6444 1998
rect 6426 1998 6444 2016
rect 6426 2016 6444 2034
rect 6426 2034 6444 2052
rect 6426 2052 6444 2070
rect 6426 2070 6444 2088
rect 6426 2088 6444 2106
rect 6426 2106 6444 2124
rect 6426 2124 6444 2142
rect 6426 2142 6444 2160
rect 6426 2160 6444 2178
rect 6426 2178 6444 2196
rect 6426 2196 6444 2214
rect 6426 2214 6444 2232
rect 6426 2232 6444 2250
rect 6426 2250 6444 2268
rect 6426 2268 6444 2286
rect 6426 2286 6444 2304
rect 6426 2304 6444 2322
rect 6426 2322 6444 2340
rect 6426 2340 6444 2358
rect 6426 2358 6444 2376
rect 6426 2376 6444 2394
rect 6426 2394 6444 2412
rect 6426 2412 6444 2430
rect 6426 2430 6444 2448
rect 6426 2448 6444 2466
rect 6426 2466 6444 2484
rect 6426 2484 6444 2502
rect 6426 2502 6444 2520
rect 6426 2520 6444 2538
rect 6426 2538 6444 2556
rect 6426 2556 6444 2574
rect 6426 2574 6444 2592
rect 6426 2592 6444 2610
rect 6426 2610 6444 2628
rect 6426 2628 6444 2646
rect 6426 2646 6444 2664
rect 6426 2664 6444 2682
rect 6426 2682 6444 2700
rect 6426 2700 6444 2718
rect 6426 2718 6444 2736
rect 6426 2736 6444 2754
rect 6426 2754 6444 2772
rect 6426 2772 6444 2790
rect 6426 2790 6444 2808
rect 6426 2808 6444 2826
rect 6426 2826 6444 2844
rect 6426 2844 6444 2862
rect 6426 2862 6444 2880
rect 6426 2880 6444 2898
rect 6426 2898 6444 2916
rect 6426 3330 6444 3348
rect 6426 3348 6444 3366
rect 6426 3366 6444 3384
rect 6426 3384 6444 3402
rect 6426 3402 6444 3420
rect 6426 3420 6444 3438
rect 6426 3438 6444 3456
rect 6426 3456 6444 3474
rect 6426 3474 6444 3492
rect 6426 3492 6444 3510
rect 6426 3510 6444 3528
rect 6426 3528 6444 3546
rect 6426 3546 6444 3564
rect 6426 3564 6444 3582
rect 6426 3582 6444 3600
rect 6426 3600 6444 3618
rect 6426 3618 6444 3636
rect 6426 3636 6444 3654
rect 6426 3654 6444 3672
rect 6426 3672 6444 3690
rect 6426 3690 6444 3708
rect 6426 3708 6444 3726
rect 6426 3726 6444 3744
rect 6426 3744 6444 3762
rect 6426 3762 6444 3780
rect 6426 3780 6444 3798
rect 6426 3798 6444 3816
rect 6426 3816 6444 3834
rect 6426 3834 6444 3852
rect 6426 3852 6444 3870
rect 6426 3870 6444 3888
rect 6426 3888 6444 3906
rect 6426 3906 6444 3924
rect 6426 3924 6444 3942
rect 6426 3942 6444 3960
rect 6426 3960 6444 3978
rect 6426 3978 6444 3996
rect 6426 3996 6444 4014
rect 6426 4014 6444 4032
rect 6426 4032 6444 4050
rect 6426 4050 6444 4068
rect 6426 4068 6444 4086
rect 6426 4086 6444 4104
rect 6426 4104 6444 4122
rect 6426 4122 6444 4140
rect 6426 4140 6444 4158
rect 6426 4158 6444 4176
rect 6426 4176 6444 4194
rect 6426 4194 6444 4212
rect 6426 4212 6444 4230
rect 6426 4230 6444 4248
rect 6426 4248 6444 4266
rect 6426 4266 6444 4284
rect 6426 4284 6444 4302
rect 6426 4302 6444 4320
rect 6426 4320 6444 4338
rect 6426 4338 6444 4356
rect 6426 4356 6444 4374
rect 6426 4374 6444 4392
rect 6426 4392 6444 4410
rect 6426 4410 6444 4428
rect 6426 4428 6444 4446
rect 6426 4446 6444 4464
rect 6426 4464 6444 4482
rect 6426 4482 6444 4500
rect 6426 4500 6444 4518
rect 6426 4518 6444 4536
rect 6426 4536 6444 4554
rect 6426 4554 6444 4572
rect 6426 4572 6444 4590
rect 6426 4590 6444 4608
rect 6426 4608 6444 4626
rect 6426 4626 6444 4644
rect 6426 4644 6444 4662
rect 6426 4662 6444 4680
rect 6426 4680 6444 4698
rect 6426 4698 6444 4716
rect 6426 4716 6444 4734
rect 6426 4734 6444 4752
rect 6426 4752 6444 4770
rect 6426 4770 6444 4788
rect 6426 4788 6444 4806
rect 6426 4806 6444 4824
rect 6426 4824 6444 4842
rect 6426 4842 6444 4860
rect 6426 4860 6444 4878
rect 6426 4878 6444 4896
rect 6426 4896 6444 4914
rect 6426 4914 6444 4932
rect 6426 4932 6444 4950
rect 6426 4950 6444 4968
rect 6426 4968 6444 4986
rect 6426 4986 6444 5004
rect 6426 5004 6444 5022
rect 6426 5022 6444 5040
rect 6426 5040 6444 5058
rect 6426 5058 6444 5076
rect 6426 5076 6444 5094
rect 6426 5094 6444 5112
rect 6426 5112 6444 5130
rect 6426 5130 6444 5148
rect 6426 5148 6444 5166
rect 6426 5166 6444 5184
rect 6426 5184 6444 5202
rect 6426 5202 6444 5220
rect 6426 5220 6444 5238
rect 6426 5238 6444 5256
rect 6426 5256 6444 5274
rect 6426 5274 6444 5292
rect 6426 5292 6444 5310
rect 6426 5310 6444 5328
rect 6426 5328 6444 5346
rect 6426 5346 6444 5364
rect 6426 5364 6444 5382
rect 6426 5382 6444 5400
rect 6426 5400 6444 5418
rect 6426 5418 6444 5436
rect 6426 5436 6444 5454
rect 6426 5454 6444 5472
rect 6426 5472 6444 5490
rect 6426 5490 6444 5508
rect 6426 5508 6444 5526
rect 6426 5526 6444 5544
rect 6426 5544 6444 5562
rect 6426 5562 6444 5580
rect 6426 5580 6444 5598
rect 6426 5598 6444 5616
rect 6426 5616 6444 5634
rect 6426 5634 6444 5652
rect 6426 5652 6444 5670
rect 6426 5670 6444 5688
rect 6426 5688 6444 5706
rect 6426 5706 6444 5724
rect 6426 5724 6444 5742
rect 6426 5742 6444 5760
rect 6426 5760 6444 5778
rect 6426 6408 6444 6426
rect 6426 6426 6444 6444
rect 6426 6444 6444 6462
rect 6426 6462 6444 6480
rect 6426 6480 6444 6498
rect 6426 6498 6444 6516
rect 6426 6516 6444 6534
rect 6426 6534 6444 6552
rect 6426 6552 6444 6570
rect 6426 6570 6444 6588
rect 6426 6588 6444 6606
rect 6426 6606 6444 6624
rect 6426 6624 6444 6642
rect 6426 6642 6444 6660
rect 6426 6660 6444 6678
rect 6426 6678 6444 6696
rect 6426 6696 6444 6714
rect 6426 6714 6444 6732
rect 6426 6732 6444 6750
rect 6426 6750 6444 6768
rect 6426 6768 6444 6786
rect 6426 6786 6444 6804
rect 6426 6804 6444 6822
rect 6426 6822 6444 6840
rect 6426 6840 6444 6858
rect 6426 6858 6444 6876
rect 6426 6876 6444 6894
rect 6426 6894 6444 6912
rect 6426 6912 6444 6930
rect 6426 6930 6444 6948
rect 6426 6948 6444 6966
rect 6426 6966 6444 6984
rect 6426 6984 6444 7002
rect 6426 7002 6444 7020
rect 6426 7020 6444 7038
rect 6426 7038 6444 7056
rect 6426 7056 6444 7074
rect 6426 7074 6444 7092
rect 6426 7092 6444 7110
rect 6426 7110 6444 7128
rect 6426 7128 6444 7146
rect 6426 7146 6444 7164
rect 6426 7164 6444 7182
rect 6426 7182 6444 7200
rect 6426 7200 6444 7218
rect 6426 7218 6444 7236
rect 6426 7236 6444 7254
rect 6426 7254 6444 7272
rect 6426 7272 6444 7290
rect 6426 7290 6444 7308
rect 6426 7308 6444 7326
rect 6426 7326 6444 7344
rect 6426 7344 6444 7362
rect 6426 7362 6444 7380
rect 6426 7380 6444 7398
rect 6426 7398 6444 7416
rect 6426 7416 6444 7434
rect 6426 7434 6444 7452
rect 6426 7452 6444 7470
rect 6426 7470 6444 7488
rect 6426 7488 6444 7506
rect 6426 7506 6444 7524
rect 6426 7524 6444 7542
rect 6426 7542 6444 7560
rect 6426 7560 6444 7578
rect 6426 7578 6444 7596
rect 6426 7596 6444 7614
rect 6426 7614 6444 7632
rect 6426 7632 6444 7650
rect 6426 7650 6444 7668
rect 6426 7668 6444 7686
rect 6426 7686 6444 7704
rect 6426 7704 6444 7722
rect 6426 7722 6444 7740
rect 6426 7740 6444 7758
rect 6426 7758 6444 7776
rect 6426 7776 6444 7794
rect 6426 7794 6444 7812
rect 6426 7812 6444 7830
rect 6426 7830 6444 7848
rect 6426 7848 6444 7866
rect 6426 7866 6444 7884
rect 6426 7884 6444 7902
rect 6426 7902 6444 7920
rect 6426 7920 6444 7938
rect 6426 7938 6444 7956
rect 6426 7956 6444 7974
rect 6426 7974 6444 7992
rect 6426 7992 6444 8010
rect 6426 8010 6444 8028
rect 6426 8028 6444 8046
rect 6426 8046 6444 8064
rect 6426 8064 6444 8082
rect 6426 8082 6444 8100
rect 6426 8100 6444 8118
rect 6426 8118 6444 8136
rect 6426 8136 6444 8154
rect 6426 8154 6444 8172
rect 6426 8172 6444 8190
rect 6426 8190 6444 8208
rect 6426 8208 6444 8226
rect 6426 8226 6444 8244
rect 6426 8244 6444 8262
rect 6426 8262 6444 8280
rect 6426 8280 6444 8298
rect 6426 8298 6444 8316
rect 6426 8316 6444 8334
rect 6426 8334 6444 8352
rect 6426 8352 6444 8370
rect 6426 8370 6444 8388
rect 6426 8388 6444 8406
rect 6426 8406 6444 8424
rect 6426 8424 6444 8442
rect 6426 8442 6444 8460
rect 6426 8460 6444 8478
rect 6426 8478 6444 8496
rect 6426 8496 6444 8514
rect 6426 8514 6444 8532
rect 6426 8532 6444 8550
rect 6426 8550 6444 8568
rect 6426 8568 6444 8586
rect 6426 8586 6444 8604
rect 6426 8604 6444 8622
rect 6426 8622 6444 8640
rect 6426 8640 6444 8658
rect 6426 8658 6444 8676
rect 6426 8676 6444 8694
rect 6426 8694 6444 8712
rect 6426 8712 6444 8730
rect 6426 8730 6444 8748
rect 6426 8748 6444 8766
rect 6426 8766 6444 8784
rect 6426 8784 6444 8802
rect 6426 8802 6444 8820
rect 6426 8820 6444 8838
rect 6426 8838 6444 8856
rect 6426 8856 6444 8874
rect 6426 8874 6444 8892
rect 6426 8892 6444 8910
rect 6426 8910 6444 8928
rect 6426 8928 6444 8946
rect 6426 8946 6444 8964
rect 6426 8964 6444 8982
rect 6426 8982 6444 9000
rect 6426 9000 6444 9018
rect 6426 9018 6444 9036
rect 6426 9036 6444 9054
rect 6426 9054 6444 9072
rect 6426 9072 6444 9090
rect 6426 9090 6444 9108
rect 6426 9108 6444 9126
rect 6426 9126 6444 9144
rect 6426 9144 6444 9162
rect 6426 9162 6444 9180
rect 6426 9180 6444 9198
rect 6426 9198 6444 9216
rect 6426 9216 6444 9234
rect 6426 9234 6444 9252
rect 6426 9252 6444 9270
rect 6426 9270 6444 9288
rect 6426 9288 6444 9306
rect 6426 9306 6444 9324
rect 6426 9324 6444 9342
rect 6426 9342 6444 9360
rect 6426 9360 6444 9378
rect 6426 9378 6444 9396
rect 6426 9396 6444 9414
rect 6426 9414 6444 9432
rect 6426 9432 6444 9450
rect 6426 9450 6444 9468
rect 6426 9468 6444 9486
rect 6426 9486 6444 9504
rect 6426 9504 6444 9522
rect 6426 9522 6444 9540
rect 6426 9540 6444 9558
rect 6426 9558 6444 9576
rect 6426 9576 6444 9594
rect 6426 9594 6444 9612
rect 6426 9612 6444 9630
rect 6426 9630 6444 9648
rect 6426 9648 6444 9666
rect 6426 9666 6444 9684
rect 6426 9684 6444 9702
rect 6426 9702 6444 9720
rect 6426 9720 6444 9738
rect 6426 9738 6444 9756
rect 6426 9756 6444 9774
rect 6444 1458 6462 1476
rect 6444 1476 6462 1494
rect 6444 1494 6462 1512
rect 6444 1512 6462 1530
rect 6444 1530 6462 1548
rect 6444 1548 6462 1566
rect 6444 1566 6462 1584
rect 6444 1584 6462 1602
rect 6444 1602 6462 1620
rect 6444 1620 6462 1638
rect 6444 1638 6462 1656
rect 6444 1656 6462 1674
rect 6444 1674 6462 1692
rect 6444 1692 6462 1710
rect 6444 1710 6462 1728
rect 6444 1728 6462 1746
rect 6444 1746 6462 1764
rect 6444 1764 6462 1782
rect 6444 1782 6462 1800
rect 6444 1800 6462 1818
rect 6444 1818 6462 1836
rect 6444 1836 6462 1854
rect 6444 1854 6462 1872
rect 6444 1872 6462 1890
rect 6444 1890 6462 1908
rect 6444 1908 6462 1926
rect 6444 1926 6462 1944
rect 6444 1944 6462 1962
rect 6444 1962 6462 1980
rect 6444 1980 6462 1998
rect 6444 1998 6462 2016
rect 6444 2016 6462 2034
rect 6444 2034 6462 2052
rect 6444 2052 6462 2070
rect 6444 2070 6462 2088
rect 6444 2088 6462 2106
rect 6444 2106 6462 2124
rect 6444 2124 6462 2142
rect 6444 2142 6462 2160
rect 6444 2160 6462 2178
rect 6444 2178 6462 2196
rect 6444 2196 6462 2214
rect 6444 2214 6462 2232
rect 6444 2232 6462 2250
rect 6444 2250 6462 2268
rect 6444 2268 6462 2286
rect 6444 2286 6462 2304
rect 6444 2304 6462 2322
rect 6444 2322 6462 2340
rect 6444 2340 6462 2358
rect 6444 2358 6462 2376
rect 6444 2376 6462 2394
rect 6444 2394 6462 2412
rect 6444 2412 6462 2430
rect 6444 2430 6462 2448
rect 6444 2448 6462 2466
rect 6444 2466 6462 2484
rect 6444 2484 6462 2502
rect 6444 2502 6462 2520
rect 6444 2520 6462 2538
rect 6444 2538 6462 2556
rect 6444 2556 6462 2574
rect 6444 2574 6462 2592
rect 6444 2592 6462 2610
rect 6444 2610 6462 2628
rect 6444 2628 6462 2646
rect 6444 2646 6462 2664
rect 6444 2664 6462 2682
rect 6444 2682 6462 2700
rect 6444 2700 6462 2718
rect 6444 2718 6462 2736
rect 6444 2736 6462 2754
rect 6444 2754 6462 2772
rect 6444 2772 6462 2790
rect 6444 2790 6462 2808
rect 6444 2808 6462 2826
rect 6444 2826 6462 2844
rect 6444 2844 6462 2862
rect 6444 2862 6462 2880
rect 6444 2880 6462 2898
rect 6444 2898 6462 2916
rect 6444 3348 6462 3366
rect 6444 3366 6462 3384
rect 6444 3384 6462 3402
rect 6444 3402 6462 3420
rect 6444 3420 6462 3438
rect 6444 3438 6462 3456
rect 6444 3456 6462 3474
rect 6444 3474 6462 3492
rect 6444 3492 6462 3510
rect 6444 3510 6462 3528
rect 6444 3528 6462 3546
rect 6444 3546 6462 3564
rect 6444 3564 6462 3582
rect 6444 3582 6462 3600
rect 6444 3600 6462 3618
rect 6444 3618 6462 3636
rect 6444 3636 6462 3654
rect 6444 3654 6462 3672
rect 6444 3672 6462 3690
rect 6444 3690 6462 3708
rect 6444 3708 6462 3726
rect 6444 3726 6462 3744
rect 6444 3744 6462 3762
rect 6444 3762 6462 3780
rect 6444 3780 6462 3798
rect 6444 3798 6462 3816
rect 6444 3816 6462 3834
rect 6444 3834 6462 3852
rect 6444 3852 6462 3870
rect 6444 3870 6462 3888
rect 6444 3888 6462 3906
rect 6444 3906 6462 3924
rect 6444 3924 6462 3942
rect 6444 3942 6462 3960
rect 6444 3960 6462 3978
rect 6444 3978 6462 3996
rect 6444 3996 6462 4014
rect 6444 4014 6462 4032
rect 6444 4032 6462 4050
rect 6444 4050 6462 4068
rect 6444 4068 6462 4086
rect 6444 4086 6462 4104
rect 6444 4104 6462 4122
rect 6444 4122 6462 4140
rect 6444 4140 6462 4158
rect 6444 4158 6462 4176
rect 6444 4176 6462 4194
rect 6444 4194 6462 4212
rect 6444 4212 6462 4230
rect 6444 4230 6462 4248
rect 6444 4248 6462 4266
rect 6444 4266 6462 4284
rect 6444 4284 6462 4302
rect 6444 4302 6462 4320
rect 6444 4320 6462 4338
rect 6444 4338 6462 4356
rect 6444 4356 6462 4374
rect 6444 4374 6462 4392
rect 6444 4392 6462 4410
rect 6444 4410 6462 4428
rect 6444 4428 6462 4446
rect 6444 4446 6462 4464
rect 6444 4464 6462 4482
rect 6444 4482 6462 4500
rect 6444 4500 6462 4518
rect 6444 4518 6462 4536
rect 6444 4536 6462 4554
rect 6444 4554 6462 4572
rect 6444 4572 6462 4590
rect 6444 4590 6462 4608
rect 6444 4608 6462 4626
rect 6444 4626 6462 4644
rect 6444 4644 6462 4662
rect 6444 4662 6462 4680
rect 6444 4680 6462 4698
rect 6444 4698 6462 4716
rect 6444 4716 6462 4734
rect 6444 4734 6462 4752
rect 6444 4752 6462 4770
rect 6444 4770 6462 4788
rect 6444 4788 6462 4806
rect 6444 4806 6462 4824
rect 6444 4824 6462 4842
rect 6444 4842 6462 4860
rect 6444 4860 6462 4878
rect 6444 4878 6462 4896
rect 6444 4896 6462 4914
rect 6444 4914 6462 4932
rect 6444 4932 6462 4950
rect 6444 4950 6462 4968
rect 6444 4968 6462 4986
rect 6444 4986 6462 5004
rect 6444 5004 6462 5022
rect 6444 5022 6462 5040
rect 6444 5040 6462 5058
rect 6444 5058 6462 5076
rect 6444 5076 6462 5094
rect 6444 5094 6462 5112
rect 6444 5112 6462 5130
rect 6444 5130 6462 5148
rect 6444 5148 6462 5166
rect 6444 5166 6462 5184
rect 6444 5184 6462 5202
rect 6444 5202 6462 5220
rect 6444 5220 6462 5238
rect 6444 5238 6462 5256
rect 6444 5256 6462 5274
rect 6444 5274 6462 5292
rect 6444 5292 6462 5310
rect 6444 5310 6462 5328
rect 6444 5328 6462 5346
rect 6444 5346 6462 5364
rect 6444 5364 6462 5382
rect 6444 5382 6462 5400
rect 6444 5400 6462 5418
rect 6444 5418 6462 5436
rect 6444 5436 6462 5454
rect 6444 5454 6462 5472
rect 6444 5472 6462 5490
rect 6444 5490 6462 5508
rect 6444 5508 6462 5526
rect 6444 5526 6462 5544
rect 6444 5544 6462 5562
rect 6444 5562 6462 5580
rect 6444 5580 6462 5598
rect 6444 5598 6462 5616
rect 6444 5616 6462 5634
rect 6444 5634 6462 5652
rect 6444 5652 6462 5670
rect 6444 5670 6462 5688
rect 6444 5688 6462 5706
rect 6444 5706 6462 5724
rect 6444 5724 6462 5742
rect 6444 5742 6462 5760
rect 6444 5760 6462 5778
rect 6444 5778 6462 5796
rect 6444 6462 6462 6480
rect 6444 6480 6462 6498
rect 6444 6498 6462 6516
rect 6444 6516 6462 6534
rect 6444 6534 6462 6552
rect 6444 6552 6462 6570
rect 6444 6570 6462 6588
rect 6444 6588 6462 6606
rect 6444 6606 6462 6624
rect 6444 6624 6462 6642
rect 6444 6642 6462 6660
rect 6444 6660 6462 6678
rect 6444 6678 6462 6696
rect 6444 6696 6462 6714
rect 6444 6714 6462 6732
rect 6444 6732 6462 6750
rect 6444 6750 6462 6768
rect 6444 6768 6462 6786
rect 6444 6786 6462 6804
rect 6444 6804 6462 6822
rect 6444 6822 6462 6840
rect 6444 6840 6462 6858
rect 6444 6858 6462 6876
rect 6444 6876 6462 6894
rect 6444 6894 6462 6912
rect 6444 6912 6462 6930
rect 6444 6930 6462 6948
rect 6444 6948 6462 6966
rect 6444 6966 6462 6984
rect 6444 6984 6462 7002
rect 6444 7002 6462 7020
rect 6444 7020 6462 7038
rect 6444 7038 6462 7056
rect 6444 7056 6462 7074
rect 6444 7074 6462 7092
rect 6444 7092 6462 7110
rect 6444 7110 6462 7128
rect 6444 7128 6462 7146
rect 6444 7146 6462 7164
rect 6444 7164 6462 7182
rect 6444 7182 6462 7200
rect 6444 7200 6462 7218
rect 6444 7218 6462 7236
rect 6444 7236 6462 7254
rect 6444 7254 6462 7272
rect 6444 7272 6462 7290
rect 6444 7290 6462 7308
rect 6444 7308 6462 7326
rect 6444 7326 6462 7344
rect 6444 7344 6462 7362
rect 6444 7362 6462 7380
rect 6444 7380 6462 7398
rect 6444 7398 6462 7416
rect 6444 7416 6462 7434
rect 6444 7434 6462 7452
rect 6444 7452 6462 7470
rect 6444 7470 6462 7488
rect 6444 7488 6462 7506
rect 6444 7506 6462 7524
rect 6444 7524 6462 7542
rect 6444 7542 6462 7560
rect 6444 7560 6462 7578
rect 6444 7578 6462 7596
rect 6444 7596 6462 7614
rect 6444 7614 6462 7632
rect 6444 7632 6462 7650
rect 6444 7650 6462 7668
rect 6444 7668 6462 7686
rect 6444 7686 6462 7704
rect 6444 7704 6462 7722
rect 6444 7722 6462 7740
rect 6444 7740 6462 7758
rect 6444 7758 6462 7776
rect 6444 7776 6462 7794
rect 6444 7794 6462 7812
rect 6444 7812 6462 7830
rect 6444 7830 6462 7848
rect 6444 7848 6462 7866
rect 6444 7866 6462 7884
rect 6444 7884 6462 7902
rect 6444 7902 6462 7920
rect 6444 7920 6462 7938
rect 6444 7938 6462 7956
rect 6444 7956 6462 7974
rect 6444 7974 6462 7992
rect 6444 7992 6462 8010
rect 6444 8010 6462 8028
rect 6444 8028 6462 8046
rect 6444 8046 6462 8064
rect 6444 8064 6462 8082
rect 6444 8082 6462 8100
rect 6444 8100 6462 8118
rect 6444 8118 6462 8136
rect 6444 8136 6462 8154
rect 6444 8154 6462 8172
rect 6444 8172 6462 8190
rect 6444 8190 6462 8208
rect 6444 8208 6462 8226
rect 6444 8226 6462 8244
rect 6444 8244 6462 8262
rect 6444 8262 6462 8280
rect 6444 8280 6462 8298
rect 6444 8298 6462 8316
rect 6444 8316 6462 8334
rect 6444 8334 6462 8352
rect 6444 8352 6462 8370
rect 6444 8370 6462 8388
rect 6444 8388 6462 8406
rect 6444 8406 6462 8424
rect 6444 8424 6462 8442
rect 6444 8442 6462 8460
rect 6444 8460 6462 8478
rect 6444 8478 6462 8496
rect 6444 8496 6462 8514
rect 6444 8514 6462 8532
rect 6444 8532 6462 8550
rect 6444 8550 6462 8568
rect 6444 8568 6462 8586
rect 6444 8586 6462 8604
rect 6444 8604 6462 8622
rect 6444 8622 6462 8640
rect 6444 8640 6462 8658
rect 6444 8658 6462 8676
rect 6444 8676 6462 8694
rect 6444 8694 6462 8712
rect 6444 8712 6462 8730
rect 6444 8730 6462 8748
rect 6444 8748 6462 8766
rect 6444 8766 6462 8784
rect 6444 8784 6462 8802
rect 6444 8802 6462 8820
rect 6444 8820 6462 8838
rect 6444 8838 6462 8856
rect 6444 8856 6462 8874
rect 6444 8874 6462 8892
rect 6444 8892 6462 8910
rect 6444 8910 6462 8928
rect 6444 8928 6462 8946
rect 6444 8946 6462 8964
rect 6444 8964 6462 8982
rect 6444 8982 6462 9000
rect 6444 9000 6462 9018
rect 6444 9018 6462 9036
rect 6444 9036 6462 9054
rect 6444 9054 6462 9072
rect 6444 9072 6462 9090
rect 6444 9090 6462 9108
rect 6444 9108 6462 9126
rect 6444 9126 6462 9144
rect 6444 9144 6462 9162
rect 6444 9162 6462 9180
rect 6444 9180 6462 9198
rect 6444 9198 6462 9216
rect 6444 9216 6462 9234
rect 6444 9234 6462 9252
rect 6444 9252 6462 9270
rect 6444 9270 6462 9288
rect 6444 9288 6462 9306
rect 6444 9306 6462 9324
rect 6444 9324 6462 9342
rect 6444 9342 6462 9360
rect 6444 9360 6462 9378
rect 6444 9378 6462 9396
rect 6444 9396 6462 9414
rect 6444 9414 6462 9432
rect 6444 9432 6462 9450
rect 6444 9450 6462 9468
rect 6444 9468 6462 9486
rect 6444 9486 6462 9504
rect 6444 9504 6462 9522
rect 6444 9522 6462 9540
rect 6444 9540 6462 9558
rect 6444 9558 6462 9576
rect 6444 9576 6462 9594
rect 6444 9594 6462 9612
rect 6444 9612 6462 9630
rect 6444 9630 6462 9648
rect 6444 9648 6462 9666
rect 6444 9666 6462 9684
rect 6444 9684 6462 9702
rect 6444 9702 6462 9720
rect 6444 9720 6462 9738
rect 6444 9738 6462 9756
rect 6444 9756 6462 9774
rect 6444 9774 6462 9792
rect 6462 1458 6480 1476
rect 6462 1476 6480 1494
rect 6462 1494 6480 1512
rect 6462 1512 6480 1530
rect 6462 1530 6480 1548
rect 6462 1548 6480 1566
rect 6462 1566 6480 1584
rect 6462 1584 6480 1602
rect 6462 1602 6480 1620
rect 6462 1620 6480 1638
rect 6462 1638 6480 1656
rect 6462 1656 6480 1674
rect 6462 1674 6480 1692
rect 6462 1692 6480 1710
rect 6462 1710 6480 1728
rect 6462 1728 6480 1746
rect 6462 1746 6480 1764
rect 6462 1764 6480 1782
rect 6462 1782 6480 1800
rect 6462 1800 6480 1818
rect 6462 1818 6480 1836
rect 6462 1836 6480 1854
rect 6462 1854 6480 1872
rect 6462 1872 6480 1890
rect 6462 1890 6480 1908
rect 6462 1908 6480 1926
rect 6462 1926 6480 1944
rect 6462 1944 6480 1962
rect 6462 1962 6480 1980
rect 6462 1980 6480 1998
rect 6462 1998 6480 2016
rect 6462 2016 6480 2034
rect 6462 2034 6480 2052
rect 6462 2052 6480 2070
rect 6462 2070 6480 2088
rect 6462 2088 6480 2106
rect 6462 2106 6480 2124
rect 6462 2124 6480 2142
rect 6462 2142 6480 2160
rect 6462 2160 6480 2178
rect 6462 2178 6480 2196
rect 6462 2196 6480 2214
rect 6462 2214 6480 2232
rect 6462 2232 6480 2250
rect 6462 2250 6480 2268
rect 6462 2268 6480 2286
rect 6462 2286 6480 2304
rect 6462 2304 6480 2322
rect 6462 2322 6480 2340
rect 6462 2340 6480 2358
rect 6462 2358 6480 2376
rect 6462 2376 6480 2394
rect 6462 2394 6480 2412
rect 6462 2412 6480 2430
rect 6462 2430 6480 2448
rect 6462 2448 6480 2466
rect 6462 2466 6480 2484
rect 6462 2484 6480 2502
rect 6462 2502 6480 2520
rect 6462 2520 6480 2538
rect 6462 2538 6480 2556
rect 6462 2556 6480 2574
rect 6462 2574 6480 2592
rect 6462 2592 6480 2610
rect 6462 2610 6480 2628
rect 6462 2628 6480 2646
rect 6462 2646 6480 2664
rect 6462 2664 6480 2682
rect 6462 2682 6480 2700
rect 6462 2700 6480 2718
rect 6462 2718 6480 2736
rect 6462 2736 6480 2754
rect 6462 2754 6480 2772
rect 6462 2772 6480 2790
rect 6462 2790 6480 2808
rect 6462 2808 6480 2826
rect 6462 2826 6480 2844
rect 6462 2844 6480 2862
rect 6462 2862 6480 2880
rect 6462 2880 6480 2898
rect 6462 2898 6480 2916
rect 6462 3366 6480 3384
rect 6462 3384 6480 3402
rect 6462 3402 6480 3420
rect 6462 3420 6480 3438
rect 6462 3438 6480 3456
rect 6462 3456 6480 3474
rect 6462 3474 6480 3492
rect 6462 3492 6480 3510
rect 6462 3510 6480 3528
rect 6462 3528 6480 3546
rect 6462 3546 6480 3564
rect 6462 3564 6480 3582
rect 6462 3582 6480 3600
rect 6462 3600 6480 3618
rect 6462 3618 6480 3636
rect 6462 3636 6480 3654
rect 6462 3654 6480 3672
rect 6462 3672 6480 3690
rect 6462 3690 6480 3708
rect 6462 3708 6480 3726
rect 6462 3726 6480 3744
rect 6462 3744 6480 3762
rect 6462 3762 6480 3780
rect 6462 3780 6480 3798
rect 6462 3798 6480 3816
rect 6462 3816 6480 3834
rect 6462 3834 6480 3852
rect 6462 3852 6480 3870
rect 6462 3870 6480 3888
rect 6462 3888 6480 3906
rect 6462 3906 6480 3924
rect 6462 3924 6480 3942
rect 6462 3942 6480 3960
rect 6462 3960 6480 3978
rect 6462 3978 6480 3996
rect 6462 3996 6480 4014
rect 6462 4014 6480 4032
rect 6462 4032 6480 4050
rect 6462 4050 6480 4068
rect 6462 4068 6480 4086
rect 6462 4086 6480 4104
rect 6462 4104 6480 4122
rect 6462 4122 6480 4140
rect 6462 4140 6480 4158
rect 6462 4158 6480 4176
rect 6462 4176 6480 4194
rect 6462 4194 6480 4212
rect 6462 4212 6480 4230
rect 6462 4230 6480 4248
rect 6462 4248 6480 4266
rect 6462 4266 6480 4284
rect 6462 4284 6480 4302
rect 6462 4302 6480 4320
rect 6462 4320 6480 4338
rect 6462 4338 6480 4356
rect 6462 4356 6480 4374
rect 6462 4374 6480 4392
rect 6462 4392 6480 4410
rect 6462 4410 6480 4428
rect 6462 4428 6480 4446
rect 6462 4446 6480 4464
rect 6462 4464 6480 4482
rect 6462 4482 6480 4500
rect 6462 4500 6480 4518
rect 6462 4518 6480 4536
rect 6462 4536 6480 4554
rect 6462 4554 6480 4572
rect 6462 4572 6480 4590
rect 6462 4590 6480 4608
rect 6462 4608 6480 4626
rect 6462 4626 6480 4644
rect 6462 4644 6480 4662
rect 6462 4662 6480 4680
rect 6462 4680 6480 4698
rect 6462 4698 6480 4716
rect 6462 4716 6480 4734
rect 6462 4734 6480 4752
rect 6462 4752 6480 4770
rect 6462 4770 6480 4788
rect 6462 4788 6480 4806
rect 6462 4806 6480 4824
rect 6462 4824 6480 4842
rect 6462 4842 6480 4860
rect 6462 4860 6480 4878
rect 6462 4878 6480 4896
rect 6462 4896 6480 4914
rect 6462 4914 6480 4932
rect 6462 4932 6480 4950
rect 6462 4950 6480 4968
rect 6462 4968 6480 4986
rect 6462 4986 6480 5004
rect 6462 5004 6480 5022
rect 6462 5022 6480 5040
rect 6462 5040 6480 5058
rect 6462 5058 6480 5076
rect 6462 5076 6480 5094
rect 6462 5094 6480 5112
rect 6462 5112 6480 5130
rect 6462 5130 6480 5148
rect 6462 5148 6480 5166
rect 6462 5166 6480 5184
rect 6462 5184 6480 5202
rect 6462 5202 6480 5220
rect 6462 5220 6480 5238
rect 6462 5238 6480 5256
rect 6462 5256 6480 5274
rect 6462 5274 6480 5292
rect 6462 5292 6480 5310
rect 6462 5310 6480 5328
rect 6462 5328 6480 5346
rect 6462 5346 6480 5364
rect 6462 5364 6480 5382
rect 6462 5382 6480 5400
rect 6462 5400 6480 5418
rect 6462 5418 6480 5436
rect 6462 5436 6480 5454
rect 6462 5454 6480 5472
rect 6462 5472 6480 5490
rect 6462 5490 6480 5508
rect 6462 5508 6480 5526
rect 6462 5526 6480 5544
rect 6462 5544 6480 5562
rect 6462 5562 6480 5580
rect 6462 5580 6480 5598
rect 6462 5598 6480 5616
rect 6462 5616 6480 5634
rect 6462 5634 6480 5652
rect 6462 5652 6480 5670
rect 6462 5670 6480 5688
rect 6462 5688 6480 5706
rect 6462 5706 6480 5724
rect 6462 5724 6480 5742
rect 6462 5742 6480 5760
rect 6462 5760 6480 5778
rect 6462 5778 6480 5796
rect 6462 6498 6480 6516
rect 6462 6516 6480 6534
rect 6462 6534 6480 6552
rect 6462 6552 6480 6570
rect 6462 6570 6480 6588
rect 6462 6588 6480 6606
rect 6462 6606 6480 6624
rect 6462 6624 6480 6642
rect 6462 6642 6480 6660
rect 6462 6660 6480 6678
rect 6462 6678 6480 6696
rect 6462 6696 6480 6714
rect 6462 6714 6480 6732
rect 6462 6732 6480 6750
rect 6462 6750 6480 6768
rect 6462 6768 6480 6786
rect 6462 6786 6480 6804
rect 6462 6804 6480 6822
rect 6462 6822 6480 6840
rect 6462 6840 6480 6858
rect 6462 6858 6480 6876
rect 6462 6876 6480 6894
rect 6462 6894 6480 6912
rect 6462 6912 6480 6930
rect 6462 6930 6480 6948
rect 6462 6948 6480 6966
rect 6462 6966 6480 6984
rect 6462 6984 6480 7002
rect 6462 7002 6480 7020
rect 6462 7020 6480 7038
rect 6462 7038 6480 7056
rect 6462 7056 6480 7074
rect 6462 7074 6480 7092
rect 6462 7092 6480 7110
rect 6462 7110 6480 7128
rect 6462 7128 6480 7146
rect 6462 7146 6480 7164
rect 6462 7164 6480 7182
rect 6462 7182 6480 7200
rect 6462 7200 6480 7218
rect 6462 7218 6480 7236
rect 6462 7236 6480 7254
rect 6462 7254 6480 7272
rect 6462 7272 6480 7290
rect 6462 7290 6480 7308
rect 6462 7308 6480 7326
rect 6462 7326 6480 7344
rect 6462 7344 6480 7362
rect 6462 7362 6480 7380
rect 6462 7380 6480 7398
rect 6462 7398 6480 7416
rect 6462 7416 6480 7434
rect 6462 7434 6480 7452
rect 6462 7452 6480 7470
rect 6462 7470 6480 7488
rect 6462 7488 6480 7506
rect 6462 7506 6480 7524
rect 6462 7524 6480 7542
rect 6462 7542 6480 7560
rect 6462 7560 6480 7578
rect 6462 7578 6480 7596
rect 6462 7596 6480 7614
rect 6462 7614 6480 7632
rect 6462 7632 6480 7650
rect 6462 7650 6480 7668
rect 6462 7668 6480 7686
rect 6462 7686 6480 7704
rect 6462 7704 6480 7722
rect 6462 7722 6480 7740
rect 6462 7740 6480 7758
rect 6462 7758 6480 7776
rect 6462 7776 6480 7794
rect 6462 7794 6480 7812
rect 6462 7812 6480 7830
rect 6462 7830 6480 7848
rect 6462 7848 6480 7866
rect 6462 7866 6480 7884
rect 6462 7884 6480 7902
rect 6462 7902 6480 7920
rect 6462 7920 6480 7938
rect 6462 7938 6480 7956
rect 6462 7956 6480 7974
rect 6462 7974 6480 7992
rect 6462 7992 6480 8010
rect 6462 8010 6480 8028
rect 6462 8028 6480 8046
rect 6462 8046 6480 8064
rect 6462 8064 6480 8082
rect 6462 8082 6480 8100
rect 6462 8100 6480 8118
rect 6462 8118 6480 8136
rect 6462 8136 6480 8154
rect 6462 8154 6480 8172
rect 6462 8172 6480 8190
rect 6462 8190 6480 8208
rect 6462 8208 6480 8226
rect 6462 8226 6480 8244
rect 6462 8244 6480 8262
rect 6462 8262 6480 8280
rect 6462 8280 6480 8298
rect 6462 8298 6480 8316
rect 6462 8316 6480 8334
rect 6462 8334 6480 8352
rect 6462 8352 6480 8370
rect 6462 8370 6480 8388
rect 6462 8388 6480 8406
rect 6462 8406 6480 8424
rect 6462 8424 6480 8442
rect 6462 8442 6480 8460
rect 6462 8460 6480 8478
rect 6462 8478 6480 8496
rect 6462 8496 6480 8514
rect 6462 8514 6480 8532
rect 6462 8532 6480 8550
rect 6462 8550 6480 8568
rect 6462 8568 6480 8586
rect 6462 8586 6480 8604
rect 6462 8604 6480 8622
rect 6462 8622 6480 8640
rect 6462 8640 6480 8658
rect 6462 8658 6480 8676
rect 6462 8676 6480 8694
rect 6462 8694 6480 8712
rect 6462 8712 6480 8730
rect 6462 8730 6480 8748
rect 6462 8748 6480 8766
rect 6462 8766 6480 8784
rect 6462 8784 6480 8802
rect 6462 8802 6480 8820
rect 6462 8820 6480 8838
rect 6462 8838 6480 8856
rect 6462 8856 6480 8874
rect 6462 8874 6480 8892
rect 6462 8892 6480 8910
rect 6462 8910 6480 8928
rect 6462 8928 6480 8946
rect 6462 8946 6480 8964
rect 6462 8964 6480 8982
rect 6462 8982 6480 9000
rect 6462 9000 6480 9018
rect 6462 9018 6480 9036
rect 6462 9036 6480 9054
rect 6462 9054 6480 9072
rect 6462 9072 6480 9090
rect 6462 9090 6480 9108
rect 6462 9108 6480 9126
rect 6462 9126 6480 9144
rect 6462 9144 6480 9162
rect 6462 9162 6480 9180
rect 6462 9180 6480 9198
rect 6462 9198 6480 9216
rect 6462 9216 6480 9234
rect 6462 9234 6480 9252
rect 6462 9252 6480 9270
rect 6462 9270 6480 9288
rect 6462 9288 6480 9306
rect 6462 9306 6480 9324
rect 6462 9324 6480 9342
rect 6462 9342 6480 9360
rect 6462 9360 6480 9378
rect 6462 9378 6480 9396
rect 6462 9396 6480 9414
rect 6462 9414 6480 9432
rect 6462 9432 6480 9450
rect 6462 9450 6480 9468
rect 6462 9468 6480 9486
rect 6462 9486 6480 9504
rect 6462 9504 6480 9522
rect 6462 9522 6480 9540
rect 6462 9540 6480 9558
rect 6462 9558 6480 9576
rect 6462 9576 6480 9594
rect 6462 9594 6480 9612
rect 6462 9612 6480 9630
rect 6462 9630 6480 9648
rect 6462 9648 6480 9666
rect 6462 9666 6480 9684
rect 6462 9684 6480 9702
rect 6462 9702 6480 9720
rect 6462 9720 6480 9738
rect 6462 9738 6480 9756
rect 6462 9756 6480 9774
rect 6462 9774 6480 9792
rect 6462 9792 6480 9810
rect 6480 1476 6498 1494
rect 6480 1494 6498 1512
rect 6480 1512 6498 1530
rect 6480 1530 6498 1548
rect 6480 1548 6498 1566
rect 6480 1566 6498 1584
rect 6480 1584 6498 1602
rect 6480 1602 6498 1620
rect 6480 1620 6498 1638
rect 6480 1638 6498 1656
rect 6480 1656 6498 1674
rect 6480 1674 6498 1692
rect 6480 1692 6498 1710
rect 6480 1710 6498 1728
rect 6480 1728 6498 1746
rect 6480 1746 6498 1764
rect 6480 1764 6498 1782
rect 6480 1782 6498 1800
rect 6480 1800 6498 1818
rect 6480 1818 6498 1836
rect 6480 1836 6498 1854
rect 6480 1854 6498 1872
rect 6480 1872 6498 1890
rect 6480 1890 6498 1908
rect 6480 1908 6498 1926
rect 6480 1926 6498 1944
rect 6480 1944 6498 1962
rect 6480 1962 6498 1980
rect 6480 1980 6498 1998
rect 6480 1998 6498 2016
rect 6480 2016 6498 2034
rect 6480 2034 6498 2052
rect 6480 2052 6498 2070
rect 6480 2070 6498 2088
rect 6480 2088 6498 2106
rect 6480 2106 6498 2124
rect 6480 2124 6498 2142
rect 6480 2142 6498 2160
rect 6480 2160 6498 2178
rect 6480 2178 6498 2196
rect 6480 2196 6498 2214
rect 6480 2214 6498 2232
rect 6480 2232 6498 2250
rect 6480 2250 6498 2268
rect 6480 2268 6498 2286
rect 6480 2286 6498 2304
rect 6480 2304 6498 2322
rect 6480 2322 6498 2340
rect 6480 2340 6498 2358
rect 6480 2358 6498 2376
rect 6480 2376 6498 2394
rect 6480 2394 6498 2412
rect 6480 2412 6498 2430
rect 6480 2430 6498 2448
rect 6480 2448 6498 2466
rect 6480 2466 6498 2484
rect 6480 2484 6498 2502
rect 6480 2502 6498 2520
rect 6480 2520 6498 2538
rect 6480 2538 6498 2556
rect 6480 2556 6498 2574
rect 6480 2574 6498 2592
rect 6480 2592 6498 2610
rect 6480 2610 6498 2628
rect 6480 2628 6498 2646
rect 6480 2646 6498 2664
rect 6480 2664 6498 2682
rect 6480 2682 6498 2700
rect 6480 2700 6498 2718
rect 6480 2718 6498 2736
rect 6480 2736 6498 2754
rect 6480 2754 6498 2772
rect 6480 2772 6498 2790
rect 6480 2790 6498 2808
rect 6480 2808 6498 2826
rect 6480 2826 6498 2844
rect 6480 2844 6498 2862
rect 6480 2862 6498 2880
rect 6480 2880 6498 2898
rect 6480 2898 6498 2916
rect 6480 2916 6498 2934
rect 6480 3384 6498 3402
rect 6480 3402 6498 3420
rect 6480 3420 6498 3438
rect 6480 3438 6498 3456
rect 6480 3456 6498 3474
rect 6480 3474 6498 3492
rect 6480 3492 6498 3510
rect 6480 3510 6498 3528
rect 6480 3528 6498 3546
rect 6480 3546 6498 3564
rect 6480 3564 6498 3582
rect 6480 3582 6498 3600
rect 6480 3600 6498 3618
rect 6480 3618 6498 3636
rect 6480 3636 6498 3654
rect 6480 3654 6498 3672
rect 6480 3672 6498 3690
rect 6480 3690 6498 3708
rect 6480 3708 6498 3726
rect 6480 3726 6498 3744
rect 6480 3744 6498 3762
rect 6480 3762 6498 3780
rect 6480 3780 6498 3798
rect 6480 3798 6498 3816
rect 6480 3816 6498 3834
rect 6480 3834 6498 3852
rect 6480 3852 6498 3870
rect 6480 3870 6498 3888
rect 6480 3888 6498 3906
rect 6480 3906 6498 3924
rect 6480 3924 6498 3942
rect 6480 3942 6498 3960
rect 6480 3960 6498 3978
rect 6480 3978 6498 3996
rect 6480 3996 6498 4014
rect 6480 4014 6498 4032
rect 6480 4032 6498 4050
rect 6480 4050 6498 4068
rect 6480 4068 6498 4086
rect 6480 4086 6498 4104
rect 6480 4104 6498 4122
rect 6480 4122 6498 4140
rect 6480 4140 6498 4158
rect 6480 4158 6498 4176
rect 6480 4176 6498 4194
rect 6480 4194 6498 4212
rect 6480 4212 6498 4230
rect 6480 4230 6498 4248
rect 6480 4248 6498 4266
rect 6480 4266 6498 4284
rect 6480 4284 6498 4302
rect 6480 4302 6498 4320
rect 6480 4320 6498 4338
rect 6480 4338 6498 4356
rect 6480 4356 6498 4374
rect 6480 4374 6498 4392
rect 6480 4392 6498 4410
rect 6480 4410 6498 4428
rect 6480 4428 6498 4446
rect 6480 4446 6498 4464
rect 6480 4464 6498 4482
rect 6480 4482 6498 4500
rect 6480 4500 6498 4518
rect 6480 4518 6498 4536
rect 6480 4536 6498 4554
rect 6480 4554 6498 4572
rect 6480 4572 6498 4590
rect 6480 4590 6498 4608
rect 6480 4608 6498 4626
rect 6480 4626 6498 4644
rect 6480 4644 6498 4662
rect 6480 4662 6498 4680
rect 6480 4680 6498 4698
rect 6480 4698 6498 4716
rect 6480 4716 6498 4734
rect 6480 4734 6498 4752
rect 6480 4752 6498 4770
rect 6480 4770 6498 4788
rect 6480 4788 6498 4806
rect 6480 4806 6498 4824
rect 6480 4824 6498 4842
rect 6480 4842 6498 4860
rect 6480 4860 6498 4878
rect 6480 4878 6498 4896
rect 6480 4896 6498 4914
rect 6480 4914 6498 4932
rect 6480 4932 6498 4950
rect 6480 4950 6498 4968
rect 6480 4968 6498 4986
rect 6480 4986 6498 5004
rect 6480 5004 6498 5022
rect 6480 5022 6498 5040
rect 6480 5040 6498 5058
rect 6480 5058 6498 5076
rect 6480 5076 6498 5094
rect 6480 5094 6498 5112
rect 6480 5112 6498 5130
rect 6480 5130 6498 5148
rect 6480 5148 6498 5166
rect 6480 5166 6498 5184
rect 6480 5184 6498 5202
rect 6480 5202 6498 5220
rect 6480 5220 6498 5238
rect 6480 5238 6498 5256
rect 6480 5256 6498 5274
rect 6480 5274 6498 5292
rect 6480 5292 6498 5310
rect 6480 5310 6498 5328
rect 6480 5328 6498 5346
rect 6480 5346 6498 5364
rect 6480 5364 6498 5382
rect 6480 5382 6498 5400
rect 6480 5400 6498 5418
rect 6480 5418 6498 5436
rect 6480 5436 6498 5454
rect 6480 5454 6498 5472
rect 6480 5472 6498 5490
rect 6480 5490 6498 5508
rect 6480 5508 6498 5526
rect 6480 5526 6498 5544
rect 6480 5544 6498 5562
rect 6480 5562 6498 5580
rect 6480 5580 6498 5598
rect 6480 5598 6498 5616
rect 6480 5616 6498 5634
rect 6480 5634 6498 5652
rect 6480 5652 6498 5670
rect 6480 5670 6498 5688
rect 6480 5688 6498 5706
rect 6480 5706 6498 5724
rect 6480 5724 6498 5742
rect 6480 5742 6498 5760
rect 6480 5760 6498 5778
rect 6480 5778 6498 5796
rect 6480 5796 6498 5814
rect 6480 6552 6498 6570
rect 6480 6570 6498 6588
rect 6480 6588 6498 6606
rect 6480 6606 6498 6624
rect 6480 6624 6498 6642
rect 6480 6642 6498 6660
rect 6480 6660 6498 6678
rect 6480 6678 6498 6696
rect 6480 6696 6498 6714
rect 6480 6714 6498 6732
rect 6480 6732 6498 6750
rect 6480 6750 6498 6768
rect 6480 6768 6498 6786
rect 6480 6786 6498 6804
rect 6480 6804 6498 6822
rect 6480 6822 6498 6840
rect 6480 6840 6498 6858
rect 6480 6858 6498 6876
rect 6480 6876 6498 6894
rect 6480 6894 6498 6912
rect 6480 6912 6498 6930
rect 6480 6930 6498 6948
rect 6480 6948 6498 6966
rect 6480 6966 6498 6984
rect 6480 6984 6498 7002
rect 6480 7002 6498 7020
rect 6480 7020 6498 7038
rect 6480 7038 6498 7056
rect 6480 7056 6498 7074
rect 6480 7074 6498 7092
rect 6480 7092 6498 7110
rect 6480 7110 6498 7128
rect 6480 7128 6498 7146
rect 6480 7146 6498 7164
rect 6480 7164 6498 7182
rect 6480 7182 6498 7200
rect 6480 7200 6498 7218
rect 6480 7218 6498 7236
rect 6480 7236 6498 7254
rect 6480 7254 6498 7272
rect 6480 7272 6498 7290
rect 6480 7290 6498 7308
rect 6480 7308 6498 7326
rect 6480 7326 6498 7344
rect 6480 7344 6498 7362
rect 6480 7362 6498 7380
rect 6480 7380 6498 7398
rect 6480 7398 6498 7416
rect 6480 7416 6498 7434
rect 6480 7434 6498 7452
rect 6480 7452 6498 7470
rect 6480 7470 6498 7488
rect 6480 7488 6498 7506
rect 6480 7506 6498 7524
rect 6480 7524 6498 7542
rect 6480 7542 6498 7560
rect 6480 7560 6498 7578
rect 6480 7578 6498 7596
rect 6480 7596 6498 7614
rect 6480 7614 6498 7632
rect 6480 7632 6498 7650
rect 6480 7650 6498 7668
rect 6480 7668 6498 7686
rect 6480 7686 6498 7704
rect 6480 7704 6498 7722
rect 6480 7722 6498 7740
rect 6480 7740 6498 7758
rect 6480 7758 6498 7776
rect 6480 7776 6498 7794
rect 6480 7794 6498 7812
rect 6480 7812 6498 7830
rect 6480 7830 6498 7848
rect 6480 7848 6498 7866
rect 6480 7866 6498 7884
rect 6480 7884 6498 7902
rect 6480 7902 6498 7920
rect 6480 7920 6498 7938
rect 6480 7938 6498 7956
rect 6480 7956 6498 7974
rect 6480 7974 6498 7992
rect 6480 7992 6498 8010
rect 6480 8010 6498 8028
rect 6480 8028 6498 8046
rect 6480 8046 6498 8064
rect 6480 8064 6498 8082
rect 6480 8082 6498 8100
rect 6480 8100 6498 8118
rect 6480 8118 6498 8136
rect 6480 8136 6498 8154
rect 6480 8154 6498 8172
rect 6480 8172 6498 8190
rect 6480 8190 6498 8208
rect 6480 8208 6498 8226
rect 6480 8226 6498 8244
rect 6480 8244 6498 8262
rect 6480 8262 6498 8280
rect 6480 8280 6498 8298
rect 6480 8298 6498 8316
rect 6480 8316 6498 8334
rect 6480 8334 6498 8352
rect 6480 8352 6498 8370
rect 6480 8370 6498 8388
rect 6480 8388 6498 8406
rect 6480 8406 6498 8424
rect 6480 8424 6498 8442
rect 6480 8442 6498 8460
rect 6480 8460 6498 8478
rect 6480 8478 6498 8496
rect 6480 8496 6498 8514
rect 6480 8514 6498 8532
rect 6480 8532 6498 8550
rect 6480 8550 6498 8568
rect 6480 8568 6498 8586
rect 6480 8586 6498 8604
rect 6480 8604 6498 8622
rect 6480 8622 6498 8640
rect 6480 8640 6498 8658
rect 6480 8658 6498 8676
rect 6480 8676 6498 8694
rect 6480 8694 6498 8712
rect 6480 8712 6498 8730
rect 6480 8730 6498 8748
rect 6480 8748 6498 8766
rect 6480 8766 6498 8784
rect 6480 8784 6498 8802
rect 6480 8802 6498 8820
rect 6480 8820 6498 8838
rect 6480 8838 6498 8856
rect 6480 8856 6498 8874
rect 6480 8874 6498 8892
rect 6480 8892 6498 8910
rect 6480 8910 6498 8928
rect 6480 8928 6498 8946
rect 6480 8946 6498 8964
rect 6480 8964 6498 8982
rect 6480 8982 6498 9000
rect 6480 9000 6498 9018
rect 6480 9018 6498 9036
rect 6480 9036 6498 9054
rect 6480 9054 6498 9072
rect 6480 9072 6498 9090
rect 6480 9090 6498 9108
rect 6480 9108 6498 9126
rect 6480 9126 6498 9144
rect 6480 9144 6498 9162
rect 6480 9162 6498 9180
rect 6480 9180 6498 9198
rect 6480 9198 6498 9216
rect 6480 9216 6498 9234
rect 6480 9234 6498 9252
rect 6480 9252 6498 9270
rect 6480 9270 6498 9288
rect 6480 9288 6498 9306
rect 6480 9306 6498 9324
rect 6480 9324 6498 9342
rect 6480 9342 6498 9360
rect 6480 9360 6498 9378
rect 6480 9378 6498 9396
rect 6480 9396 6498 9414
rect 6480 9414 6498 9432
rect 6480 9432 6498 9450
rect 6480 9450 6498 9468
rect 6480 9468 6498 9486
rect 6480 9486 6498 9504
rect 6480 9504 6498 9522
rect 6480 9522 6498 9540
rect 6480 9540 6498 9558
rect 6480 9558 6498 9576
rect 6480 9576 6498 9594
rect 6480 9594 6498 9612
rect 6480 9612 6498 9630
rect 6480 9630 6498 9648
rect 6480 9648 6498 9666
rect 6480 9666 6498 9684
rect 6480 9684 6498 9702
rect 6480 9702 6498 9720
rect 6480 9720 6498 9738
rect 6480 9738 6498 9756
rect 6480 9756 6498 9774
rect 6480 9774 6498 9792
rect 6480 9792 6498 9810
rect 6480 9810 6498 9828
rect 6480 9828 6498 9846
rect 6498 1494 6516 1512
rect 6498 1512 6516 1530
rect 6498 1530 6516 1548
rect 6498 1548 6516 1566
rect 6498 1566 6516 1584
rect 6498 1584 6516 1602
rect 6498 1602 6516 1620
rect 6498 1620 6516 1638
rect 6498 1638 6516 1656
rect 6498 1656 6516 1674
rect 6498 1674 6516 1692
rect 6498 1692 6516 1710
rect 6498 1710 6516 1728
rect 6498 1728 6516 1746
rect 6498 1746 6516 1764
rect 6498 1764 6516 1782
rect 6498 1782 6516 1800
rect 6498 1800 6516 1818
rect 6498 1818 6516 1836
rect 6498 1836 6516 1854
rect 6498 1854 6516 1872
rect 6498 1872 6516 1890
rect 6498 1890 6516 1908
rect 6498 1908 6516 1926
rect 6498 1926 6516 1944
rect 6498 1944 6516 1962
rect 6498 1962 6516 1980
rect 6498 1980 6516 1998
rect 6498 1998 6516 2016
rect 6498 2016 6516 2034
rect 6498 2034 6516 2052
rect 6498 2052 6516 2070
rect 6498 2070 6516 2088
rect 6498 2088 6516 2106
rect 6498 2106 6516 2124
rect 6498 2124 6516 2142
rect 6498 2142 6516 2160
rect 6498 2160 6516 2178
rect 6498 2178 6516 2196
rect 6498 2196 6516 2214
rect 6498 2214 6516 2232
rect 6498 2232 6516 2250
rect 6498 2250 6516 2268
rect 6498 2268 6516 2286
rect 6498 2286 6516 2304
rect 6498 2304 6516 2322
rect 6498 2322 6516 2340
rect 6498 2340 6516 2358
rect 6498 2358 6516 2376
rect 6498 2376 6516 2394
rect 6498 2394 6516 2412
rect 6498 2412 6516 2430
rect 6498 2430 6516 2448
rect 6498 2448 6516 2466
rect 6498 2466 6516 2484
rect 6498 2484 6516 2502
rect 6498 2502 6516 2520
rect 6498 2520 6516 2538
rect 6498 2538 6516 2556
rect 6498 2556 6516 2574
rect 6498 2574 6516 2592
rect 6498 2592 6516 2610
rect 6498 2610 6516 2628
rect 6498 2628 6516 2646
rect 6498 2646 6516 2664
rect 6498 2664 6516 2682
rect 6498 2682 6516 2700
rect 6498 2700 6516 2718
rect 6498 2718 6516 2736
rect 6498 2736 6516 2754
rect 6498 2754 6516 2772
rect 6498 2772 6516 2790
rect 6498 2790 6516 2808
rect 6498 2808 6516 2826
rect 6498 2826 6516 2844
rect 6498 2844 6516 2862
rect 6498 2862 6516 2880
rect 6498 2880 6516 2898
rect 6498 2898 6516 2916
rect 6498 2916 6516 2934
rect 6498 3420 6516 3438
rect 6498 3438 6516 3456
rect 6498 3456 6516 3474
rect 6498 3474 6516 3492
rect 6498 3492 6516 3510
rect 6498 3510 6516 3528
rect 6498 3528 6516 3546
rect 6498 3546 6516 3564
rect 6498 3564 6516 3582
rect 6498 3582 6516 3600
rect 6498 3600 6516 3618
rect 6498 3618 6516 3636
rect 6498 3636 6516 3654
rect 6498 3654 6516 3672
rect 6498 3672 6516 3690
rect 6498 3690 6516 3708
rect 6498 3708 6516 3726
rect 6498 3726 6516 3744
rect 6498 3744 6516 3762
rect 6498 3762 6516 3780
rect 6498 3780 6516 3798
rect 6498 3798 6516 3816
rect 6498 3816 6516 3834
rect 6498 3834 6516 3852
rect 6498 3852 6516 3870
rect 6498 3870 6516 3888
rect 6498 3888 6516 3906
rect 6498 3906 6516 3924
rect 6498 3924 6516 3942
rect 6498 3942 6516 3960
rect 6498 3960 6516 3978
rect 6498 3978 6516 3996
rect 6498 3996 6516 4014
rect 6498 4014 6516 4032
rect 6498 4032 6516 4050
rect 6498 4050 6516 4068
rect 6498 4068 6516 4086
rect 6498 4086 6516 4104
rect 6498 4104 6516 4122
rect 6498 4122 6516 4140
rect 6498 4140 6516 4158
rect 6498 4158 6516 4176
rect 6498 4176 6516 4194
rect 6498 4194 6516 4212
rect 6498 4212 6516 4230
rect 6498 4230 6516 4248
rect 6498 4248 6516 4266
rect 6498 4266 6516 4284
rect 6498 4284 6516 4302
rect 6498 4302 6516 4320
rect 6498 4320 6516 4338
rect 6498 4338 6516 4356
rect 6498 4356 6516 4374
rect 6498 4374 6516 4392
rect 6498 4392 6516 4410
rect 6498 4410 6516 4428
rect 6498 4428 6516 4446
rect 6498 4446 6516 4464
rect 6498 4464 6516 4482
rect 6498 4482 6516 4500
rect 6498 4500 6516 4518
rect 6498 4518 6516 4536
rect 6498 4536 6516 4554
rect 6498 4554 6516 4572
rect 6498 4572 6516 4590
rect 6498 4590 6516 4608
rect 6498 4608 6516 4626
rect 6498 4626 6516 4644
rect 6498 4644 6516 4662
rect 6498 4662 6516 4680
rect 6498 4680 6516 4698
rect 6498 4698 6516 4716
rect 6498 4716 6516 4734
rect 6498 4734 6516 4752
rect 6498 4752 6516 4770
rect 6498 4770 6516 4788
rect 6498 4788 6516 4806
rect 6498 4806 6516 4824
rect 6498 4824 6516 4842
rect 6498 4842 6516 4860
rect 6498 4860 6516 4878
rect 6498 4878 6516 4896
rect 6498 4896 6516 4914
rect 6498 4914 6516 4932
rect 6498 4932 6516 4950
rect 6498 4950 6516 4968
rect 6498 4968 6516 4986
rect 6498 4986 6516 5004
rect 6498 5004 6516 5022
rect 6498 5022 6516 5040
rect 6498 5040 6516 5058
rect 6498 5058 6516 5076
rect 6498 5076 6516 5094
rect 6498 5094 6516 5112
rect 6498 5112 6516 5130
rect 6498 5130 6516 5148
rect 6498 5148 6516 5166
rect 6498 5166 6516 5184
rect 6498 5184 6516 5202
rect 6498 5202 6516 5220
rect 6498 5220 6516 5238
rect 6498 5238 6516 5256
rect 6498 5256 6516 5274
rect 6498 5274 6516 5292
rect 6498 5292 6516 5310
rect 6498 5310 6516 5328
rect 6498 5328 6516 5346
rect 6498 5346 6516 5364
rect 6498 5364 6516 5382
rect 6498 5382 6516 5400
rect 6498 5400 6516 5418
rect 6498 5418 6516 5436
rect 6498 5436 6516 5454
rect 6498 5454 6516 5472
rect 6498 5472 6516 5490
rect 6498 5490 6516 5508
rect 6498 5508 6516 5526
rect 6498 5526 6516 5544
rect 6498 5544 6516 5562
rect 6498 5562 6516 5580
rect 6498 5580 6516 5598
rect 6498 5598 6516 5616
rect 6498 5616 6516 5634
rect 6498 5634 6516 5652
rect 6498 5652 6516 5670
rect 6498 5670 6516 5688
rect 6498 5688 6516 5706
rect 6498 5706 6516 5724
rect 6498 5724 6516 5742
rect 6498 5742 6516 5760
rect 6498 5760 6516 5778
rect 6498 5778 6516 5796
rect 6498 5796 6516 5814
rect 6498 5814 6516 5832
rect 6498 6588 6516 6606
rect 6498 6606 6516 6624
rect 6498 6624 6516 6642
rect 6498 6642 6516 6660
rect 6498 6660 6516 6678
rect 6498 6678 6516 6696
rect 6498 6696 6516 6714
rect 6498 6714 6516 6732
rect 6498 6732 6516 6750
rect 6498 6750 6516 6768
rect 6498 6768 6516 6786
rect 6498 6786 6516 6804
rect 6498 6804 6516 6822
rect 6498 6822 6516 6840
rect 6498 6840 6516 6858
rect 6498 6858 6516 6876
rect 6498 6876 6516 6894
rect 6498 6894 6516 6912
rect 6498 6912 6516 6930
rect 6498 6930 6516 6948
rect 6498 6948 6516 6966
rect 6498 6966 6516 6984
rect 6498 6984 6516 7002
rect 6498 7002 6516 7020
rect 6498 7020 6516 7038
rect 6498 7038 6516 7056
rect 6498 7056 6516 7074
rect 6498 7074 6516 7092
rect 6498 7092 6516 7110
rect 6498 7110 6516 7128
rect 6498 7128 6516 7146
rect 6498 7146 6516 7164
rect 6498 7164 6516 7182
rect 6498 7182 6516 7200
rect 6498 7200 6516 7218
rect 6498 7218 6516 7236
rect 6498 7236 6516 7254
rect 6498 7254 6516 7272
rect 6498 7272 6516 7290
rect 6498 7290 6516 7308
rect 6498 7308 6516 7326
rect 6498 7326 6516 7344
rect 6498 7344 6516 7362
rect 6498 7362 6516 7380
rect 6498 7380 6516 7398
rect 6498 7398 6516 7416
rect 6498 7416 6516 7434
rect 6498 7434 6516 7452
rect 6498 7452 6516 7470
rect 6498 7470 6516 7488
rect 6498 7488 6516 7506
rect 6498 7506 6516 7524
rect 6498 7524 6516 7542
rect 6498 7542 6516 7560
rect 6498 7560 6516 7578
rect 6498 7578 6516 7596
rect 6498 7596 6516 7614
rect 6498 7614 6516 7632
rect 6498 7632 6516 7650
rect 6498 7650 6516 7668
rect 6498 7668 6516 7686
rect 6498 7686 6516 7704
rect 6498 7704 6516 7722
rect 6498 7722 6516 7740
rect 6498 7740 6516 7758
rect 6498 7758 6516 7776
rect 6498 7776 6516 7794
rect 6498 7794 6516 7812
rect 6498 7812 6516 7830
rect 6498 7830 6516 7848
rect 6498 7848 6516 7866
rect 6498 7866 6516 7884
rect 6498 7884 6516 7902
rect 6498 7902 6516 7920
rect 6498 7920 6516 7938
rect 6498 7938 6516 7956
rect 6498 7956 6516 7974
rect 6498 7974 6516 7992
rect 6498 7992 6516 8010
rect 6498 8010 6516 8028
rect 6498 8028 6516 8046
rect 6498 8046 6516 8064
rect 6498 8064 6516 8082
rect 6498 8082 6516 8100
rect 6498 8100 6516 8118
rect 6498 8118 6516 8136
rect 6498 8136 6516 8154
rect 6498 8154 6516 8172
rect 6498 8172 6516 8190
rect 6498 8190 6516 8208
rect 6498 8208 6516 8226
rect 6498 8226 6516 8244
rect 6498 8244 6516 8262
rect 6498 8262 6516 8280
rect 6498 8280 6516 8298
rect 6498 8298 6516 8316
rect 6498 8316 6516 8334
rect 6498 8334 6516 8352
rect 6498 8352 6516 8370
rect 6498 8370 6516 8388
rect 6498 8388 6516 8406
rect 6498 8406 6516 8424
rect 6498 8424 6516 8442
rect 6498 8442 6516 8460
rect 6498 8460 6516 8478
rect 6498 8478 6516 8496
rect 6498 8496 6516 8514
rect 6498 8514 6516 8532
rect 6498 8532 6516 8550
rect 6498 8550 6516 8568
rect 6498 8568 6516 8586
rect 6498 8586 6516 8604
rect 6498 8604 6516 8622
rect 6498 8622 6516 8640
rect 6498 8640 6516 8658
rect 6498 8658 6516 8676
rect 6498 8676 6516 8694
rect 6498 8694 6516 8712
rect 6498 8712 6516 8730
rect 6498 8730 6516 8748
rect 6498 8748 6516 8766
rect 6498 8766 6516 8784
rect 6498 8784 6516 8802
rect 6498 8802 6516 8820
rect 6498 8820 6516 8838
rect 6498 8838 6516 8856
rect 6498 8856 6516 8874
rect 6498 8874 6516 8892
rect 6498 8892 6516 8910
rect 6498 8910 6516 8928
rect 6498 8928 6516 8946
rect 6498 8946 6516 8964
rect 6498 8964 6516 8982
rect 6498 8982 6516 9000
rect 6498 9000 6516 9018
rect 6498 9018 6516 9036
rect 6498 9036 6516 9054
rect 6498 9054 6516 9072
rect 6498 9072 6516 9090
rect 6498 9090 6516 9108
rect 6498 9108 6516 9126
rect 6498 9126 6516 9144
rect 6498 9144 6516 9162
rect 6498 9162 6516 9180
rect 6498 9180 6516 9198
rect 6498 9198 6516 9216
rect 6498 9216 6516 9234
rect 6498 9234 6516 9252
rect 6498 9252 6516 9270
rect 6498 9270 6516 9288
rect 6498 9288 6516 9306
rect 6498 9306 6516 9324
rect 6498 9324 6516 9342
rect 6498 9342 6516 9360
rect 6498 9360 6516 9378
rect 6498 9378 6516 9396
rect 6498 9396 6516 9414
rect 6498 9414 6516 9432
rect 6498 9432 6516 9450
rect 6498 9450 6516 9468
rect 6498 9468 6516 9486
rect 6498 9486 6516 9504
rect 6498 9504 6516 9522
rect 6498 9522 6516 9540
rect 6498 9540 6516 9558
rect 6498 9558 6516 9576
rect 6498 9576 6516 9594
rect 6498 9594 6516 9612
rect 6498 9612 6516 9630
rect 6498 9630 6516 9648
rect 6498 9648 6516 9666
rect 6498 9666 6516 9684
rect 6498 9684 6516 9702
rect 6498 9702 6516 9720
rect 6498 9720 6516 9738
rect 6498 9738 6516 9756
rect 6498 9756 6516 9774
rect 6498 9774 6516 9792
rect 6498 9792 6516 9810
rect 6498 9810 6516 9828
rect 6498 9828 6516 9846
rect 6498 9846 6516 9864
rect 6516 1494 6534 1512
rect 6516 1512 6534 1530
rect 6516 1530 6534 1548
rect 6516 1548 6534 1566
rect 6516 1566 6534 1584
rect 6516 1584 6534 1602
rect 6516 1602 6534 1620
rect 6516 1620 6534 1638
rect 6516 1638 6534 1656
rect 6516 1656 6534 1674
rect 6516 1674 6534 1692
rect 6516 1692 6534 1710
rect 6516 1710 6534 1728
rect 6516 1728 6534 1746
rect 6516 1746 6534 1764
rect 6516 1764 6534 1782
rect 6516 1782 6534 1800
rect 6516 1800 6534 1818
rect 6516 1818 6534 1836
rect 6516 1836 6534 1854
rect 6516 1854 6534 1872
rect 6516 1872 6534 1890
rect 6516 1890 6534 1908
rect 6516 1908 6534 1926
rect 6516 1926 6534 1944
rect 6516 1944 6534 1962
rect 6516 1962 6534 1980
rect 6516 1980 6534 1998
rect 6516 1998 6534 2016
rect 6516 2016 6534 2034
rect 6516 2034 6534 2052
rect 6516 2052 6534 2070
rect 6516 2070 6534 2088
rect 6516 2088 6534 2106
rect 6516 2106 6534 2124
rect 6516 2124 6534 2142
rect 6516 2142 6534 2160
rect 6516 2160 6534 2178
rect 6516 2178 6534 2196
rect 6516 2196 6534 2214
rect 6516 2214 6534 2232
rect 6516 2232 6534 2250
rect 6516 2250 6534 2268
rect 6516 2268 6534 2286
rect 6516 2286 6534 2304
rect 6516 2304 6534 2322
rect 6516 2322 6534 2340
rect 6516 2340 6534 2358
rect 6516 2358 6534 2376
rect 6516 2376 6534 2394
rect 6516 2394 6534 2412
rect 6516 2412 6534 2430
rect 6516 2430 6534 2448
rect 6516 2448 6534 2466
rect 6516 2466 6534 2484
rect 6516 2484 6534 2502
rect 6516 2502 6534 2520
rect 6516 2520 6534 2538
rect 6516 2538 6534 2556
rect 6516 2556 6534 2574
rect 6516 2574 6534 2592
rect 6516 2592 6534 2610
rect 6516 2610 6534 2628
rect 6516 2628 6534 2646
rect 6516 2646 6534 2664
rect 6516 2664 6534 2682
rect 6516 2682 6534 2700
rect 6516 2700 6534 2718
rect 6516 2718 6534 2736
rect 6516 2736 6534 2754
rect 6516 2754 6534 2772
rect 6516 2772 6534 2790
rect 6516 2790 6534 2808
rect 6516 2808 6534 2826
rect 6516 2826 6534 2844
rect 6516 2844 6534 2862
rect 6516 2862 6534 2880
rect 6516 2880 6534 2898
rect 6516 2898 6534 2916
rect 6516 2916 6534 2934
rect 6516 3438 6534 3456
rect 6516 3456 6534 3474
rect 6516 3474 6534 3492
rect 6516 3492 6534 3510
rect 6516 3510 6534 3528
rect 6516 3528 6534 3546
rect 6516 3546 6534 3564
rect 6516 3564 6534 3582
rect 6516 3582 6534 3600
rect 6516 3600 6534 3618
rect 6516 3618 6534 3636
rect 6516 3636 6534 3654
rect 6516 3654 6534 3672
rect 6516 3672 6534 3690
rect 6516 3690 6534 3708
rect 6516 3708 6534 3726
rect 6516 3726 6534 3744
rect 6516 3744 6534 3762
rect 6516 3762 6534 3780
rect 6516 3780 6534 3798
rect 6516 3798 6534 3816
rect 6516 3816 6534 3834
rect 6516 3834 6534 3852
rect 6516 3852 6534 3870
rect 6516 3870 6534 3888
rect 6516 3888 6534 3906
rect 6516 3906 6534 3924
rect 6516 3924 6534 3942
rect 6516 3942 6534 3960
rect 6516 3960 6534 3978
rect 6516 3978 6534 3996
rect 6516 3996 6534 4014
rect 6516 4014 6534 4032
rect 6516 4032 6534 4050
rect 6516 4050 6534 4068
rect 6516 4068 6534 4086
rect 6516 4086 6534 4104
rect 6516 4104 6534 4122
rect 6516 4122 6534 4140
rect 6516 4140 6534 4158
rect 6516 4158 6534 4176
rect 6516 4176 6534 4194
rect 6516 4194 6534 4212
rect 6516 4212 6534 4230
rect 6516 4230 6534 4248
rect 6516 4248 6534 4266
rect 6516 4266 6534 4284
rect 6516 4284 6534 4302
rect 6516 4302 6534 4320
rect 6516 4320 6534 4338
rect 6516 4338 6534 4356
rect 6516 4356 6534 4374
rect 6516 4374 6534 4392
rect 6516 4392 6534 4410
rect 6516 4410 6534 4428
rect 6516 4428 6534 4446
rect 6516 4446 6534 4464
rect 6516 4464 6534 4482
rect 6516 4482 6534 4500
rect 6516 4500 6534 4518
rect 6516 4518 6534 4536
rect 6516 4536 6534 4554
rect 6516 4554 6534 4572
rect 6516 4572 6534 4590
rect 6516 4590 6534 4608
rect 6516 4608 6534 4626
rect 6516 4626 6534 4644
rect 6516 4644 6534 4662
rect 6516 4662 6534 4680
rect 6516 4680 6534 4698
rect 6516 4698 6534 4716
rect 6516 4716 6534 4734
rect 6516 4734 6534 4752
rect 6516 4752 6534 4770
rect 6516 4770 6534 4788
rect 6516 4788 6534 4806
rect 6516 4806 6534 4824
rect 6516 4824 6534 4842
rect 6516 4842 6534 4860
rect 6516 4860 6534 4878
rect 6516 4878 6534 4896
rect 6516 4896 6534 4914
rect 6516 4914 6534 4932
rect 6516 4932 6534 4950
rect 6516 4950 6534 4968
rect 6516 4968 6534 4986
rect 6516 4986 6534 5004
rect 6516 5004 6534 5022
rect 6516 5022 6534 5040
rect 6516 5040 6534 5058
rect 6516 5058 6534 5076
rect 6516 5076 6534 5094
rect 6516 5094 6534 5112
rect 6516 5112 6534 5130
rect 6516 5130 6534 5148
rect 6516 5148 6534 5166
rect 6516 5166 6534 5184
rect 6516 5184 6534 5202
rect 6516 5202 6534 5220
rect 6516 5220 6534 5238
rect 6516 5238 6534 5256
rect 6516 5256 6534 5274
rect 6516 5274 6534 5292
rect 6516 5292 6534 5310
rect 6516 5310 6534 5328
rect 6516 5328 6534 5346
rect 6516 5346 6534 5364
rect 6516 5364 6534 5382
rect 6516 5382 6534 5400
rect 6516 5400 6534 5418
rect 6516 5418 6534 5436
rect 6516 5436 6534 5454
rect 6516 5454 6534 5472
rect 6516 5472 6534 5490
rect 6516 5490 6534 5508
rect 6516 5508 6534 5526
rect 6516 5526 6534 5544
rect 6516 5544 6534 5562
rect 6516 5562 6534 5580
rect 6516 5580 6534 5598
rect 6516 5598 6534 5616
rect 6516 5616 6534 5634
rect 6516 5634 6534 5652
rect 6516 5652 6534 5670
rect 6516 5670 6534 5688
rect 6516 5688 6534 5706
rect 6516 5706 6534 5724
rect 6516 5724 6534 5742
rect 6516 5742 6534 5760
rect 6516 5760 6534 5778
rect 6516 5778 6534 5796
rect 6516 5796 6534 5814
rect 6516 5814 6534 5832
rect 6516 5832 6534 5850
rect 6516 6624 6534 6642
rect 6516 6642 6534 6660
rect 6516 6660 6534 6678
rect 6516 6678 6534 6696
rect 6516 6696 6534 6714
rect 6516 6714 6534 6732
rect 6516 6732 6534 6750
rect 6516 6750 6534 6768
rect 6516 6768 6534 6786
rect 6516 6786 6534 6804
rect 6516 6804 6534 6822
rect 6516 6822 6534 6840
rect 6516 6840 6534 6858
rect 6516 6858 6534 6876
rect 6516 6876 6534 6894
rect 6516 6894 6534 6912
rect 6516 6912 6534 6930
rect 6516 6930 6534 6948
rect 6516 6948 6534 6966
rect 6516 6966 6534 6984
rect 6516 6984 6534 7002
rect 6516 7002 6534 7020
rect 6516 7020 6534 7038
rect 6516 7038 6534 7056
rect 6516 7056 6534 7074
rect 6516 7074 6534 7092
rect 6516 7092 6534 7110
rect 6516 7110 6534 7128
rect 6516 7128 6534 7146
rect 6516 7146 6534 7164
rect 6516 7164 6534 7182
rect 6516 7182 6534 7200
rect 6516 7200 6534 7218
rect 6516 7218 6534 7236
rect 6516 7236 6534 7254
rect 6516 7254 6534 7272
rect 6516 7272 6534 7290
rect 6516 7290 6534 7308
rect 6516 7308 6534 7326
rect 6516 7326 6534 7344
rect 6516 7344 6534 7362
rect 6516 7362 6534 7380
rect 6516 7380 6534 7398
rect 6516 7398 6534 7416
rect 6516 7416 6534 7434
rect 6516 7434 6534 7452
rect 6516 7452 6534 7470
rect 6516 7470 6534 7488
rect 6516 7488 6534 7506
rect 6516 7506 6534 7524
rect 6516 7524 6534 7542
rect 6516 7542 6534 7560
rect 6516 7560 6534 7578
rect 6516 7578 6534 7596
rect 6516 7596 6534 7614
rect 6516 7614 6534 7632
rect 6516 7632 6534 7650
rect 6516 7650 6534 7668
rect 6516 7668 6534 7686
rect 6516 7686 6534 7704
rect 6516 7704 6534 7722
rect 6516 7722 6534 7740
rect 6516 7740 6534 7758
rect 6516 7758 6534 7776
rect 6516 7776 6534 7794
rect 6516 7794 6534 7812
rect 6516 7812 6534 7830
rect 6516 7830 6534 7848
rect 6516 7848 6534 7866
rect 6516 7866 6534 7884
rect 6516 7884 6534 7902
rect 6516 7902 6534 7920
rect 6516 7920 6534 7938
rect 6516 7938 6534 7956
rect 6516 7956 6534 7974
rect 6516 7974 6534 7992
rect 6516 7992 6534 8010
rect 6516 8010 6534 8028
rect 6516 8028 6534 8046
rect 6516 8046 6534 8064
rect 6516 8064 6534 8082
rect 6516 8082 6534 8100
rect 6516 8100 6534 8118
rect 6516 8118 6534 8136
rect 6516 8136 6534 8154
rect 6516 8154 6534 8172
rect 6516 8172 6534 8190
rect 6516 8190 6534 8208
rect 6516 8208 6534 8226
rect 6516 8226 6534 8244
rect 6516 8244 6534 8262
rect 6516 8262 6534 8280
rect 6516 8280 6534 8298
rect 6516 8298 6534 8316
rect 6516 8316 6534 8334
rect 6516 8334 6534 8352
rect 6516 8352 6534 8370
rect 6516 8370 6534 8388
rect 6516 8388 6534 8406
rect 6516 8406 6534 8424
rect 6516 8424 6534 8442
rect 6516 8442 6534 8460
rect 6516 8460 6534 8478
rect 6516 8478 6534 8496
rect 6516 8496 6534 8514
rect 6516 8514 6534 8532
rect 6516 8532 6534 8550
rect 6516 8550 6534 8568
rect 6516 8568 6534 8586
rect 6516 8586 6534 8604
rect 6516 8604 6534 8622
rect 6516 8622 6534 8640
rect 6516 8640 6534 8658
rect 6516 8658 6534 8676
rect 6516 8676 6534 8694
rect 6516 8694 6534 8712
rect 6516 8712 6534 8730
rect 6516 8730 6534 8748
rect 6516 8748 6534 8766
rect 6516 8766 6534 8784
rect 6516 8784 6534 8802
rect 6516 8802 6534 8820
rect 6516 8820 6534 8838
rect 6516 8838 6534 8856
rect 6516 8856 6534 8874
rect 6516 8874 6534 8892
rect 6516 8892 6534 8910
rect 6516 8910 6534 8928
rect 6516 8928 6534 8946
rect 6516 8946 6534 8964
rect 6516 8964 6534 8982
rect 6516 8982 6534 9000
rect 6516 9000 6534 9018
rect 6516 9018 6534 9036
rect 6516 9036 6534 9054
rect 6516 9054 6534 9072
rect 6516 9072 6534 9090
rect 6516 9090 6534 9108
rect 6516 9108 6534 9126
rect 6516 9126 6534 9144
rect 6516 9144 6534 9162
rect 6516 9162 6534 9180
rect 6516 9180 6534 9198
rect 6516 9198 6534 9216
rect 6516 9216 6534 9234
rect 6516 9234 6534 9252
rect 6516 9252 6534 9270
rect 6516 9270 6534 9288
rect 6516 9288 6534 9306
rect 6516 9306 6534 9324
rect 6516 9324 6534 9342
rect 6516 9342 6534 9360
rect 6516 9360 6534 9378
rect 6516 9378 6534 9396
rect 6516 9396 6534 9414
rect 6516 9414 6534 9432
rect 6516 9432 6534 9450
rect 6516 9450 6534 9468
rect 6516 9468 6534 9486
rect 6516 9486 6534 9504
rect 6516 9504 6534 9522
rect 6516 9522 6534 9540
rect 6516 9540 6534 9558
rect 6516 9558 6534 9576
rect 6516 9576 6534 9594
rect 6516 9594 6534 9612
rect 6516 9612 6534 9630
rect 6516 9630 6534 9648
rect 6516 9648 6534 9666
rect 6516 9666 6534 9684
rect 6516 9684 6534 9702
rect 6516 9702 6534 9720
rect 6516 9720 6534 9738
rect 6516 9738 6534 9756
rect 6516 9756 6534 9774
rect 6516 9774 6534 9792
rect 6516 9792 6534 9810
rect 6516 9810 6534 9828
rect 6516 9828 6534 9846
rect 6516 9846 6534 9864
rect 6516 9864 6534 9882
rect 6534 1512 6552 1530
rect 6534 1530 6552 1548
rect 6534 1548 6552 1566
rect 6534 1566 6552 1584
rect 6534 1584 6552 1602
rect 6534 1602 6552 1620
rect 6534 1620 6552 1638
rect 6534 1638 6552 1656
rect 6534 1656 6552 1674
rect 6534 1674 6552 1692
rect 6534 1692 6552 1710
rect 6534 1710 6552 1728
rect 6534 1728 6552 1746
rect 6534 1746 6552 1764
rect 6534 1764 6552 1782
rect 6534 1782 6552 1800
rect 6534 1800 6552 1818
rect 6534 1818 6552 1836
rect 6534 1836 6552 1854
rect 6534 1854 6552 1872
rect 6534 1872 6552 1890
rect 6534 1890 6552 1908
rect 6534 1908 6552 1926
rect 6534 1926 6552 1944
rect 6534 1944 6552 1962
rect 6534 1962 6552 1980
rect 6534 1980 6552 1998
rect 6534 1998 6552 2016
rect 6534 2016 6552 2034
rect 6534 2034 6552 2052
rect 6534 2052 6552 2070
rect 6534 2070 6552 2088
rect 6534 2088 6552 2106
rect 6534 2106 6552 2124
rect 6534 2124 6552 2142
rect 6534 2142 6552 2160
rect 6534 2160 6552 2178
rect 6534 2178 6552 2196
rect 6534 2196 6552 2214
rect 6534 2214 6552 2232
rect 6534 2232 6552 2250
rect 6534 2250 6552 2268
rect 6534 2268 6552 2286
rect 6534 2286 6552 2304
rect 6534 2304 6552 2322
rect 6534 2322 6552 2340
rect 6534 2340 6552 2358
rect 6534 2358 6552 2376
rect 6534 2376 6552 2394
rect 6534 2394 6552 2412
rect 6534 2412 6552 2430
rect 6534 2430 6552 2448
rect 6534 2448 6552 2466
rect 6534 2466 6552 2484
rect 6534 2484 6552 2502
rect 6534 2502 6552 2520
rect 6534 2520 6552 2538
rect 6534 2538 6552 2556
rect 6534 2556 6552 2574
rect 6534 2574 6552 2592
rect 6534 2592 6552 2610
rect 6534 2610 6552 2628
rect 6534 2628 6552 2646
rect 6534 2646 6552 2664
rect 6534 2664 6552 2682
rect 6534 2682 6552 2700
rect 6534 2700 6552 2718
rect 6534 2718 6552 2736
rect 6534 2736 6552 2754
rect 6534 2754 6552 2772
rect 6534 2772 6552 2790
rect 6534 2790 6552 2808
rect 6534 2808 6552 2826
rect 6534 2826 6552 2844
rect 6534 2844 6552 2862
rect 6534 2862 6552 2880
rect 6534 2880 6552 2898
rect 6534 2898 6552 2916
rect 6534 2916 6552 2934
rect 6534 2934 6552 2952
rect 6534 3456 6552 3474
rect 6534 3474 6552 3492
rect 6534 3492 6552 3510
rect 6534 3510 6552 3528
rect 6534 3528 6552 3546
rect 6534 3546 6552 3564
rect 6534 3564 6552 3582
rect 6534 3582 6552 3600
rect 6534 3600 6552 3618
rect 6534 3618 6552 3636
rect 6534 3636 6552 3654
rect 6534 3654 6552 3672
rect 6534 3672 6552 3690
rect 6534 3690 6552 3708
rect 6534 3708 6552 3726
rect 6534 3726 6552 3744
rect 6534 3744 6552 3762
rect 6534 3762 6552 3780
rect 6534 3780 6552 3798
rect 6534 3798 6552 3816
rect 6534 3816 6552 3834
rect 6534 3834 6552 3852
rect 6534 3852 6552 3870
rect 6534 3870 6552 3888
rect 6534 3888 6552 3906
rect 6534 3906 6552 3924
rect 6534 3924 6552 3942
rect 6534 3942 6552 3960
rect 6534 3960 6552 3978
rect 6534 3978 6552 3996
rect 6534 3996 6552 4014
rect 6534 4014 6552 4032
rect 6534 4032 6552 4050
rect 6534 4050 6552 4068
rect 6534 4068 6552 4086
rect 6534 4086 6552 4104
rect 6534 4104 6552 4122
rect 6534 4122 6552 4140
rect 6534 4140 6552 4158
rect 6534 4158 6552 4176
rect 6534 4176 6552 4194
rect 6534 4194 6552 4212
rect 6534 4212 6552 4230
rect 6534 4230 6552 4248
rect 6534 4248 6552 4266
rect 6534 4266 6552 4284
rect 6534 4284 6552 4302
rect 6534 4302 6552 4320
rect 6534 4320 6552 4338
rect 6534 4338 6552 4356
rect 6534 4356 6552 4374
rect 6534 4374 6552 4392
rect 6534 4392 6552 4410
rect 6534 4410 6552 4428
rect 6534 4428 6552 4446
rect 6534 4446 6552 4464
rect 6534 4464 6552 4482
rect 6534 4482 6552 4500
rect 6534 4500 6552 4518
rect 6534 4518 6552 4536
rect 6534 4536 6552 4554
rect 6534 4554 6552 4572
rect 6534 4572 6552 4590
rect 6534 4590 6552 4608
rect 6534 4608 6552 4626
rect 6534 4626 6552 4644
rect 6534 4644 6552 4662
rect 6534 4662 6552 4680
rect 6534 4680 6552 4698
rect 6534 4698 6552 4716
rect 6534 4716 6552 4734
rect 6534 4734 6552 4752
rect 6534 4752 6552 4770
rect 6534 4770 6552 4788
rect 6534 4788 6552 4806
rect 6534 4806 6552 4824
rect 6534 4824 6552 4842
rect 6534 4842 6552 4860
rect 6534 4860 6552 4878
rect 6534 4878 6552 4896
rect 6534 4896 6552 4914
rect 6534 4914 6552 4932
rect 6534 4932 6552 4950
rect 6534 4950 6552 4968
rect 6534 4968 6552 4986
rect 6534 4986 6552 5004
rect 6534 5004 6552 5022
rect 6534 5022 6552 5040
rect 6534 5040 6552 5058
rect 6534 5058 6552 5076
rect 6534 5076 6552 5094
rect 6534 5094 6552 5112
rect 6534 5112 6552 5130
rect 6534 5130 6552 5148
rect 6534 5148 6552 5166
rect 6534 5166 6552 5184
rect 6534 5184 6552 5202
rect 6534 5202 6552 5220
rect 6534 5220 6552 5238
rect 6534 5238 6552 5256
rect 6534 5256 6552 5274
rect 6534 5274 6552 5292
rect 6534 5292 6552 5310
rect 6534 5310 6552 5328
rect 6534 5328 6552 5346
rect 6534 5346 6552 5364
rect 6534 5364 6552 5382
rect 6534 5382 6552 5400
rect 6534 5400 6552 5418
rect 6534 5418 6552 5436
rect 6534 5436 6552 5454
rect 6534 5454 6552 5472
rect 6534 5472 6552 5490
rect 6534 5490 6552 5508
rect 6534 5508 6552 5526
rect 6534 5526 6552 5544
rect 6534 5544 6552 5562
rect 6534 5562 6552 5580
rect 6534 5580 6552 5598
rect 6534 5598 6552 5616
rect 6534 5616 6552 5634
rect 6534 5634 6552 5652
rect 6534 5652 6552 5670
rect 6534 5670 6552 5688
rect 6534 5688 6552 5706
rect 6534 5706 6552 5724
rect 6534 5724 6552 5742
rect 6534 5742 6552 5760
rect 6534 5760 6552 5778
rect 6534 5778 6552 5796
rect 6534 5796 6552 5814
rect 6534 5814 6552 5832
rect 6534 5832 6552 5850
rect 6534 5850 6552 5868
rect 6534 6678 6552 6696
rect 6534 6696 6552 6714
rect 6534 6714 6552 6732
rect 6534 6732 6552 6750
rect 6534 6750 6552 6768
rect 6534 6768 6552 6786
rect 6534 6786 6552 6804
rect 6534 6804 6552 6822
rect 6534 6822 6552 6840
rect 6534 6840 6552 6858
rect 6534 6858 6552 6876
rect 6534 6876 6552 6894
rect 6534 6894 6552 6912
rect 6534 6912 6552 6930
rect 6534 6930 6552 6948
rect 6534 6948 6552 6966
rect 6534 6966 6552 6984
rect 6534 6984 6552 7002
rect 6534 7002 6552 7020
rect 6534 7020 6552 7038
rect 6534 7038 6552 7056
rect 6534 7056 6552 7074
rect 6534 7074 6552 7092
rect 6534 7092 6552 7110
rect 6534 7110 6552 7128
rect 6534 7128 6552 7146
rect 6534 7146 6552 7164
rect 6534 7164 6552 7182
rect 6534 7182 6552 7200
rect 6534 7200 6552 7218
rect 6534 7218 6552 7236
rect 6534 7236 6552 7254
rect 6534 7254 6552 7272
rect 6534 7272 6552 7290
rect 6534 7290 6552 7308
rect 6534 7308 6552 7326
rect 6534 7326 6552 7344
rect 6534 7344 6552 7362
rect 6534 7362 6552 7380
rect 6534 7380 6552 7398
rect 6534 7398 6552 7416
rect 6534 7416 6552 7434
rect 6534 7434 6552 7452
rect 6534 7452 6552 7470
rect 6534 7470 6552 7488
rect 6534 7488 6552 7506
rect 6534 7506 6552 7524
rect 6534 7524 6552 7542
rect 6534 7542 6552 7560
rect 6534 7560 6552 7578
rect 6534 7578 6552 7596
rect 6534 7596 6552 7614
rect 6534 7614 6552 7632
rect 6534 7632 6552 7650
rect 6534 7650 6552 7668
rect 6534 7668 6552 7686
rect 6534 7686 6552 7704
rect 6534 7704 6552 7722
rect 6534 7722 6552 7740
rect 6534 7740 6552 7758
rect 6534 7758 6552 7776
rect 6534 7776 6552 7794
rect 6534 7794 6552 7812
rect 6534 7812 6552 7830
rect 6534 7830 6552 7848
rect 6534 7848 6552 7866
rect 6534 7866 6552 7884
rect 6534 7884 6552 7902
rect 6534 7902 6552 7920
rect 6534 7920 6552 7938
rect 6534 7938 6552 7956
rect 6534 7956 6552 7974
rect 6534 7974 6552 7992
rect 6534 7992 6552 8010
rect 6534 8010 6552 8028
rect 6534 8028 6552 8046
rect 6534 8046 6552 8064
rect 6534 8064 6552 8082
rect 6534 8082 6552 8100
rect 6534 8100 6552 8118
rect 6534 8118 6552 8136
rect 6534 8136 6552 8154
rect 6534 8154 6552 8172
rect 6534 8172 6552 8190
rect 6534 8190 6552 8208
rect 6534 8208 6552 8226
rect 6534 8226 6552 8244
rect 6534 8244 6552 8262
rect 6534 8262 6552 8280
rect 6534 8280 6552 8298
rect 6534 8298 6552 8316
rect 6534 8316 6552 8334
rect 6534 8334 6552 8352
rect 6534 8352 6552 8370
rect 6534 8370 6552 8388
rect 6534 8388 6552 8406
rect 6534 8406 6552 8424
rect 6534 8424 6552 8442
rect 6534 8442 6552 8460
rect 6534 8460 6552 8478
rect 6534 8478 6552 8496
rect 6534 8496 6552 8514
rect 6534 8514 6552 8532
rect 6534 8532 6552 8550
rect 6534 8550 6552 8568
rect 6534 8568 6552 8586
rect 6534 8586 6552 8604
rect 6534 8604 6552 8622
rect 6534 8622 6552 8640
rect 6534 8640 6552 8658
rect 6534 8658 6552 8676
rect 6534 8676 6552 8694
rect 6534 8694 6552 8712
rect 6534 8712 6552 8730
rect 6534 8730 6552 8748
rect 6534 8748 6552 8766
rect 6534 8766 6552 8784
rect 6534 8784 6552 8802
rect 6534 8802 6552 8820
rect 6534 8820 6552 8838
rect 6534 8838 6552 8856
rect 6534 8856 6552 8874
rect 6534 8874 6552 8892
rect 6534 8892 6552 8910
rect 6534 8910 6552 8928
rect 6534 8928 6552 8946
rect 6534 8946 6552 8964
rect 6534 8964 6552 8982
rect 6534 8982 6552 9000
rect 6534 9000 6552 9018
rect 6534 9018 6552 9036
rect 6534 9036 6552 9054
rect 6534 9054 6552 9072
rect 6534 9072 6552 9090
rect 6534 9090 6552 9108
rect 6534 9108 6552 9126
rect 6534 9126 6552 9144
rect 6534 9144 6552 9162
rect 6534 9162 6552 9180
rect 6534 9180 6552 9198
rect 6534 9198 6552 9216
rect 6534 9216 6552 9234
rect 6534 9234 6552 9252
rect 6534 9252 6552 9270
rect 6534 9270 6552 9288
rect 6534 9288 6552 9306
rect 6534 9306 6552 9324
rect 6534 9324 6552 9342
rect 6534 9342 6552 9360
rect 6534 9360 6552 9378
rect 6534 9378 6552 9396
rect 6534 9396 6552 9414
rect 6534 9414 6552 9432
rect 6534 9432 6552 9450
rect 6534 9450 6552 9468
rect 6534 9468 6552 9486
rect 6534 9486 6552 9504
rect 6534 9504 6552 9522
rect 6534 9522 6552 9540
rect 6534 9540 6552 9558
rect 6534 9558 6552 9576
rect 6534 9576 6552 9594
rect 6534 9594 6552 9612
rect 6534 9612 6552 9630
rect 6534 9630 6552 9648
rect 6534 9648 6552 9666
rect 6534 9666 6552 9684
rect 6534 9684 6552 9702
rect 6534 9702 6552 9720
rect 6534 9720 6552 9738
rect 6534 9738 6552 9756
rect 6534 9756 6552 9774
rect 6534 9774 6552 9792
rect 6534 9792 6552 9810
rect 6534 9810 6552 9828
rect 6534 9828 6552 9846
rect 6534 9846 6552 9864
rect 6534 9864 6552 9882
rect 6534 9882 6552 9900
rect 6552 1512 6570 1530
rect 6552 1530 6570 1548
rect 6552 1548 6570 1566
rect 6552 1566 6570 1584
rect 6552 1584 6570 1602
rect 6552 1602 6570 1620
rect 6552 1620 6570 1638
rect 6552 1638 6570 1656
rect 6552 1656 6570 1674
rect 6552 1674 6570 1692
rect 6552 1692 6570 1710
rect 6552 1710 6570 1728
rect 6552 1728 6570 1746
rect 6552 1746 6570 1764
rect 6552 1764 6570 1782
rect 6552 1782 6570 1800
rect 6552 1800 6570 1818
rect 6552 1818 6570 1836
rect 6552 1836 6570 1854
rect 6552 1854 6570 1872
rect 6552 1872 6570 1890
rect 6552 1890 6570 1908
rect 6552 1908 6570 1926
rect 6552 1926 6570 1944
rect 6552 1944 6570 1962
rect 6552 1962 6570 1980
rect 6552 1980 6570 1998
rect 6552 1998 6570 2016
rect 6552 2016 6570 2034
rect 6552 2034 6570 2052
rect 6552 2052 6570 2070
rect 6552 2070 6570 2088
rect 6552 2088 6570 2106
rect 6552 2106 6570 2124
rect 6552 2124 6570 2142
rect 6552 2142 6570 2160
rect 6552 2160 6570 2178
rect 6552 2178 6570 2196
rect 6552 2196 6570 2214
rect 6552 2214 6570 2232
rect 6552 2232 6570 2250
rect 6552 2250 6570 2268
rect 6552 2268 6570 2286
rect 6552 2286 6570 2304
rect 6552 2304 6570 2322
rect 6552 2322 6570 2340
rect 6552 2340 6570 2358
rect 6552 2358 6570 2376
rect 6552 2376 6570 2394
rect 6552 2394 6570 2412
rect 6552 2412 6570 2430
rect 6552 2430 6570 2448
rect 6552 2448 6570 2466
rect 6552 2466 6570 2484
rect 6552 2484 6570 2502
rect 6552 2502 6570 2520
rect 6552 2520 6570 2538
rect 6552 2538 6570 2556
rect 6552 2556 6570 2574
rect 6552 2574 6570 2592
rect 6552 2592 6570 2610
rect 6552 2610 6570 2628
rect 6552 2628 6570 2646
rect 6552 2646 6570 2664
rect 6552 2664 6570 2682
rect 6552 2682 6570 2700
rect 6552 2700 6570 2718
rect 6552 2718 6570 2736
rect 6552 2736 6570 2754
rect 6552 2754 6570 2772
rect 6552 2772 6570 2790
rect 6552 2790 6570 2808
rect 6552 2808 6570 2826
rect 6552 2826 6570 2844
rect 6552 2844 6570 2862
rect 6552 2862 6570 2880
rect 6552 2880 6570 2898
rect 6552 2898 6570 2916
rect 6552 2916 6570 2934
rect 6552 2934 6570 2952
rect 6552 3474 6570 3492
rect 6552 3492 6570 3510
rect 6552 3510 6570 3528
rect 6552 3528 6570 3546
rect 6552 3546 6570 3564
rect 6552 3564 6570 3582
rect 6552 3582 6570 3600
rect 6552 3600 6570 3618
rect 6552 3618 6570 3636
rect 6552 3636 6570 3654
rect 6552 3654 6570 3672
rect 6552 3672 6570 3690
rect 6552 3690 6570 3708
rect 6552 3708 6570 3726
rect 6552 3726 6570 3744
rect 6552 3744 6570 3762
rect 6552 3762 6570 3780
rect 6552 3780 6570 3798
rect 6552 3798 6570 3816
rect 6552 3816 6570 3834
rect 6552 3834 6570 3852
rect 6552 3852 6570 3870
rect 6552 3870 6570 3888
rect 6552 3888 6570 3906
rect 6552 3906 6570 3924
rect 6552 3924 6570 3942
rect 6552 3942 6570 3960
rect 6552 3960 6570 3978
rect 6552 3978 6570 3996
rect 6552 3996 6570 4014
rect 6552 4014 6570 4032
rect 6552 4032 6570 4050
rect 6552 4050 6570 4068
rect 6552 4068 6570 4086
rect 6552 4086 6570 4104
rect 6552 4104 6570 4122
rect 6552 4122 6570 4140
rect 6552 4140 6570 4158
rect 6552 4158 6570 4176
rect 6552 4176 6570 4194
rect 6552 4194 6570 4212
rect 6552 4212 6570 4230
rect 6552 4230 6570 4248
rect 6552 4248 6570 4266
rect 6552 4266 6570 4284
rect 6552 4284 6570 4302
rect 6552 4302 6570 4320
rect 6552 4320 6570 4338
rect 6552 4338 6570 4356
rect 6552 4356 6570 4374
rect 6552 4374 6570 4392
rect 6552 4392 6570 4410
rect 6552 4410 6570 4428
rect 6552 4428 6570 4446
rect 6552 4446 6570 4464
rect 6552 4464 6570 4482
rect 6552 4482 6570 4500
rect 6552 4500 6570 4518
rect 6552 4518 6570 4536
rect 6552 4536 6570 4554
rect 6552 4554 6570 4572
rect 6552 4572 6570 4590
rect 6552 4590 6570 4608
rect 6552 4608 6570 4626
rect 6552 4626 6570 4644
rect 6552 4644 6570 4662
rect 6552 4662 6570 4680
rect 6552 4680 6570 4698
rect 6552 4698 6570 4716
rect 6552 4716 6570 4734
rect 6552 4734 6570 4752
rect 6552 4752 6570 4770
rect 6552 4770 6570 4788
rect 6552 4788 6570 4806
rect 6552 4806 6570 4824
rect 6552 4824 6570 4842
rect 6552 4842 6570 4860
rect 6552 4860 6570 4878
rect 6552 4878 6570 4896
rect 6552 4896 6570 4914
rect 6552 4914 6570 4932
rect 6552 4932 6570 4950
rect 6552 4950 6570 4968
rect 6552 4968 6570 4986
rect 6552 4986 6570 5004
rect 6552 5004 6570 5022
rect 6552 5022 6570 5040
rect 6552 5040 6570 5058
rect 6552 5058 6570 5076
rect 6552 5076 6570 5094
rect 6552 5094 6570 5112
rect 6552 5112 6570 5130
rect 6552 5130 6570 5148
rect 6552 5148 6570 5166
rect 6552 5166 6570 5184
rect 6552 5184 6570 5202
rect 6552 5202 6570 5220
rect 6552 5220 6570 5238
rect 6552 5238 6570 5256
rect 6552 5256 6570 5274
rect 6552 5274 6570 5292
rect 6552 5292 6570 5310
rect 6552 5310 6570 5328
rect 6552 5328 6570 5346
rect 6552 5346 6570 5364
rect 6552 5364 6570 5382
rect 6552 5382 6570 5400
rect 6552 5400 6570 5418
rect 6552 5418 6570 5436
rect 6552 5436 6570 5454
rect 6552 5454 6570 5472
rect 6552 5472 6570 5490
rect 6552 5490 6570 5508
rect 6552 5508 6570 5526
rect 6552 5526 6570 5544
rect 6552 5544 6570 5562
rect 6552 5562 6570 5580
rect 6552 5580 6570 5598
rect 6552 5598 6570 5616
rect 6552 5616 6570 5634
rect 6552 5634 6570 5652
rect 6552 5652 6570 5670
rect 6552 5670 6570 5688
rect 6552 5688 6570 5706
rect 6552 5706 6570 5724
rect 6552 5724 6570 5742
rect 6552 5742 6570 5760
rect 6552 5760 6570 5778
rect 6552 5778 6570 5796
rect 6552 5796 6570 5814
rect 6552 5814 6570 5832
rect 6552 5832 6570 5850
rect 6552 5850 6570 5868
rect 6552 5868 6570 5886
rect 6552 6714 6570 6732
rect 6552 6732 6570 6750
rect 6552 6750 6570 6768
rect 6552 6768 6570 6786
rect 6552 6786 6570 6804
rect 6552 6804 6570 6822
rect 6552 6822 6570 6840
rect 6552 6840 6570 6858
rect 6552 6858 6570 6876
rect 6552 6876 6570 6894
rect 6552 6894 6570 6912
rect 6552 6912 6570 6930
rect 6552 6930 6570 6948
rect 6552 6948 6570 6966
rect 6552 6966 6570 6984
rect 6552 6984 6570 7002
rect 6552 7002 6570 7020
rect 6552 7020 6570 7038
rect 6552 7038 6570 7056
rect 6552 7056 6570 7074
rect 6552 7074 6570 7092
rect 6552 7092 6570 7110
rect 6552 7110 6570 7128
rect 6552 7128 6570 7146
rect 6552 7146 6570 7164
rect 6552 7164 6570 7182
rect 6552 7182 6570 7200
rect 6552 7200 6570 7218
rect 6552 7218 6570 7236
rect 6552 7236 6570 7254
rect 6552 7254 6570 7272
rect 6552 7272 6570 7290
rect 6552 7290 6570 7308
rect 6552 7308 6570 7326
rect 6552 7326 6570 7344
rect 6552 7344 6570 7362
rect 6552 7362 6570 7380
rect 6552 7380 6570 7398
rect 6552 7398 6570 7416
rect 6552 7416 6570 7434
rect 6552 7434 6570 7452
rect 6552 7452 6570 7470
rect 6552 7470 6570 7488
rect 6552 7488 6570 7506
rect 6552 7506 6570 7524
rect 6552 7524 6570 7542
rect 6552 7542 6570 7560
rect 6552 7560 6570 7578
rect 6552 7578 6570 7596
rect 6552 7596 6570 7614
rect 6552 7614 6570 7632
rect 6552 7632 6570 7650
rect 6552 7650 6570 7668
rect 6552 7668 6570 7686
rect 6552 7686 6570 7704
rect 6552 7704 6570 7722
rect 6552 7722 6570 7740
rect 6552 7740 6570 7758
rect 6552 7758 6570 7776
rect 6552 7776 6570 7794
rect 6552 7794 6570 7812
rect 6552 7812 6570 7830
rect 6552 7830 6570 7848
rect 6552 7848 6570 7866
rect 6552 7866 6570 7884
rect 6552 7884 6570 7902
rect 6552 7902 6570 7920
rect 6552 7920 6570 7938
rect 6552 7938 6570 7956
rect 6552 7956 6570 7974
rect 6552 7974 6570 7992
rect 6552 7992 6570 8010
rect 6552 8010 6570 8028
rect 6552 8028 6570 8046
rect 6552 8046 6570 8064
rect 6552 8064 6570 8082
rect 6552 8082 6570 8100
rect 6552 8100 6570 8118
rect 6552 8118 6570 8136
rect 6552 8136 6570 8154
rect 6552 8154 6570 8172
rect 6552 8172 6570 8190
rect 6552 8190 6570 8208
rect 6552 8208 6570 8226
rect 6552 8226 6570 8244
rect 6552 8244 6570 8262
rect 6552 8262 6570 8280
rect 6552 8280 6570 8298
rect 6552 8298 6570 8316
rect 6552 8316 6570 8334
rect 6552 8334 6570 8352
rect 6552 8352 6570 8370
rect 6552 8370 6570 8388
rect 6552 8388 6570 8406
rect 6552 8406 6570 8424
rect 6552 8424 6570 8442
rect 6552 8442 6570 8460
rect 6552 8460 6570 8478
rect 6552 8478 6570 8496
rect 6552 8496 6570 8514
rect 6552 8514 6570 8532
rect 6552 8532 6570 8550
rect 6552 8550 6570 8568
rect 6552 8568 6570 8586
rect 6552 8586 6570 8604
rect 6552 8604 6570 8622
rect 6552 8622 6570 8640
rect 6552 8640 6570 8658
rect 6552 8658 6570 8676
rect 6552 8676 6570 8694
rect 6552 8694 6570 8712
rect 6552 8712 6570 8730
rect 6552 8730 6570 8748
rect 6552 8748 6570 8766
rect 6552 8766 6570 8784
rect 6552 8784 6570 8802
rect 6552 8802 6570 8820
rect 6552 8820 6570 8838
rect 6552 8838 6570 8856
rect 6552 8856 6570 8874
rect 6552 8874 6570 8892
rect 6552 8892 6570 8910
rect 6552 8910 6570 8928
rect 6552 8928 6570 8946
rect 6552 8946 6570 8964
rect 6552 8964 6570 8982
rect 6552 8982 6570 9000
rect 6552 9000 6570 9018
rect 6552 9018 6570 9036
rect 6552 9036 6570 9054
rect 6552 9054 6570 9072
rect 6552 9072 6570 9090
rect 6552 9090 6570 9108
rect 6552 9108 6570 9126
rect 6552 9126 6570 9144
rect 6552 9144 6570 9162
rect 6552 9162 6570 9180
rect 6552 9180 6570 9198
rect 6552 9198 6570 9216
rect 6552 9216 6570 9234
rect 6552 9234 6570 9252
rect 6552 9252 6570 9270
rect 6552 9270 6570 9288
rect 6552 9288 6570 9306
rect 6552 9306 6570 9324
rect 6552 9324 6570 9342
rect 6552 9342 6570 9360
rect 6552 9360 6570 9378
rect 6552 9378 6570 9396
rect 6552 9396 6570 9414
rect 6552 9414 6570 9432
rect 6552 9432 6570 9450
rect 6552 9450 6570 9468
rect 6552 9468 6570 9486
rect 6552 9486 6570 9504
rect 6552 9504 6570 9522
rect 6552 9522 6570 9540
rect 6552 9540 6570 9558
rect 6552 9558 6570 9576
rect 6552 9576 6570 9594
rect 6552 9594 6570 9612
rect 6552 9612 6570 9630
rect 6552 9630 6570 9648
rect 6552 9648 6570 9666
rect 6552 9666 6570 9684
rect 6552 9684 6570 9702
rect 6552 9702 6570 9720
rect 6552 9720 6570 9738
rect 6552 9738 6570 9756
rect 6552 9756 6570 9774
rect 6552 9774 6570 9792
rect 6552 9792 6570 9810
rect 6552 9810 6570 9828
rect 6552 9828 6570 9846
rect 6552 9846 6570 9864
rect 6552 9864 6570 9882
rect 6552 9882 6570 9900
rect 6552 9900 6570 9918
rect 6552 9918 6570 9936
rect 6570 1530 6588 1548
rect 6570 1548 6588 1566
rect 6570 1566 6588 1584
rect 6570 1584 6588 1602
rect 6570 1602 6588 1620
rect 6570 1620 6588 1638
rect 6570 1638 6588 1656
rect 6570 1656 6588 1674
rect 6570 1674 6588 1692
rect 6570 1692 6588 1710
rect 6570 1710 6588 1728
rect 6570 1728 6588 1746
rect 6570 1746 6588 1764
rect 6570 1764 6588 1782
rect 6570 1782 6588 1800
rect 6570 1800 6588 1818
rect 6570 1818 6588 1836
rect 6570 1836 6588 1854
rect 6570 1854 6588 1872
rect 6570 1872 6588 1890
rect 6570 1890 6588 1908
rect 6570 1908 6588 1926
rect 6570 1926 6588 1944
rect 6570 1944 6588 1962
rect 6570 1962 6588 1980
rect 6570 1980 6588 1998
rect 6570 1998 6588 2016
rect 6570 2016 6588 2034
rect 6570 2034 6588 2052
rect 6570 2052 6588 2070
rect 6570 2070 6588 2088
rect 6570 2088 6588 2106
rect 6570 2106 6588 2124
rect 6570 2124 6588 2142
rect 6570 2142 6588 2160
rect 6570 2160 6588 2178
rect 6570 2178 6588 2196
rect 6570 2196 6588 2214
rect 6570 2214 6588 2232
rect 6570 2232 6588 2250
rect 6570 2250 6588 2268
rect 6570 2268 6588 2286
rect 6570 2286 6588 2304
rect 6570 2304 6588 2322
rect 6570 2322 6588 2340
rect 6570 2340 6588 2358
rect 6570 2358 6588 2376
rect 6570 2376 6588 2394
rect 6570 2394 6588 2412
rect 6570 2412 6588 2430
rect 6570 2430 6588 2448
rect 6570 2448 6588 2466
rect 6570 2466 6588 2484
rect 6570 2484 6588 2502
rect 6570 2502 6588 2520
rect 6570 2520 6588 2538
rect 6570 2538 6588 2556
rect 6570 2556 6588 2574
rect 6570 2574 6588 2592
rect 6570 2592 6588 2610
rect 6570 2610 6588 2628
rect 6570 2628 6588 2646
rect 6570 2646 6588 2664
rect 6570 2664 6588 2682
rect 6570 2682 6588 2700
rect 6570 2700 6588 2718
rect 6570 2718 6588 2736
rect 6570 2736 6588 2754
rect 6570 2754 6588 2772
rect 6570 2772 6588 2790
rect 6570 2790 6588 2808
rect 6570 2808 6588 2826
rect 6570 2826 6588 2844
rect 6570 2844 6588 2862
rect 6570 2862 6588 2880
rect 6570 2880 6588 2898
rect 6570 2898 6588 2916
rect 6570 2916 6588 2934
rect 6570 2934 6588 2952
rect 6570 3492 6588 3510
rect 6570 3510 6588 3528
rect 6570 3528 6588 3546
rect 6570 3546 6588 3564
rect 6570 3564 6588 3582
rect 6570 3582 6588 3600
rect 6570 3600 6588 3618
rect 6570 3618 6588 3636
rect 6570 3636 6588 3654
rect 6570 3654 6588 3672
rect 6570 3672 6588 3690
rect 6570 3690 6588 3708
rect 6570 3708 6588 3726
rect 6570 3726 6588 3744
rect 6570 3744 6588 3762
rect 6570 3762 6588 3780
rect 6570 3780 6588 3798
rect 6570 3798 6588 3816
rect 6570 3816 6588 3834
rect 6570 3834 6588 3852
rect 6570 3852 6588 3870
rect 6570 3870 6588 3888
rect 6570 3888 6588 3906
rect 6570 3906 6588 3924
rect 6570 3924 6588 3942
rect 6570 3942 6588 3960
rect 6570 3960 6588 3978
rect 6570 3978 6588 3996
rect 6570 3996 6588 4014
rect 6570 4014 6588 4032
rect 6570 4032 6588 4050
rect 6570 4050 6588 4068
rect 6570 4068 6588 4086
rect 6570 4086 6588 4104
rect 6570 4104 6588 4122
rect 6570 4122 6588 4140
rect 6570 4140 6588 4158
rect 6570 4158 6588 4176
rect 6570 4176 6588 4194
rect 6570 4194 6588 4212
rect 6570 4212 6588 4230
rect 6570 4230 6588 4248
rect 6570 4248 6588 4266
rect 6570 4266 6588 4284
rect 6570 4284 6588 4302
rect 6570 4302 6588 4320
rect 6570 4320 6588 4338
rect 6570 4338 6588 4356
rect 6570 4356 6588 4374
rect 6570 4374 6588 4392
rect 6570 4392 6588 4410
rect 6570 4410 6588 4428
rect 6570 4428 6588 4446
rect 6570 4446 6588 4464
rect 6570 4464 6588 4482
rect 6570 4482 6588 4500
rect 6570 4500 6588 4518
rect 6570 4518 6588 4536
rect 6570 4536 6588 4554
rect 6570 4554 6588 4572
rect 6570 4572 6588 4590
rect 6570 4590 6588 4608
rect 6570 4608 6588 4626
rect 6570 4626 6588 4644
rect 6570 4644 6588 4662
rect 6570 4662 6588 4680
rect 6570 4680 6588 4698
rect 6570 4698 6588 4716
rect 6570 4716 6588 4734
rect 6570 4734 6588 4752
rect 6570 4752 6588 4770
rect 6570 4770 6588 4788
rect 6570 4788 6588 4806
rect 6570 4806 6588 4824
rect 6570 4824 6588 4842
rect 6570 4842 6588 4860
rect 6570 4860 6588 4878
rect 6570 4878 6588 4896
rect 6570 4896 6588 4914
rect 6570 4914 6588 4932
rect 6570 4932 6588 4950
rect 6570 4950 6588 4968
rect 6570 4968 6588 4986
rect 6570 4986 6588 5004
rect 6570 5004 6588 5022
rect 6570 5022 6588 5040
rect 6570 5040 6588 5058
rect 6570 5058 6588 5076
rect 6570 5076 6588 5094
rect 6570 5094 6588 5112
rect 6570 5112 6588 5130
rect 6570 5130 6588 5148
rect 6570 5148 6588 5166
rect 6570 5166 6588 5184
rect 6570 5184 6588 5202
rect 6570 5202 6588 5220
rect 6570 5220 6588 5238
rect 6570 5238 6588 5256
rect 6570 5256 6588 5274
rect 6570 5274 6588 5292
rect 6570 5292 6588 5310
rect 6570 5310 6588 5328
rect 6570 5328 6588 5346
rect 6570 5346 6588 5364
rect 6570 5364 6588 5382
rect 6570 5382 6588 5400
rect 6570 5400 6588 5418
rect 6570 5418 6588 5436
rect 6570 5436 6588 5454
rect 6570 5454 6588 5472
rect 6570 5472 6588 5490
rect 6570 5490 6588 5508
rect 6570 5508 6588 5526
rect 6570 5526 6588 5544
rect 6570 5544 6588 5562
rect 6570 5562 6588 5580
rect 6570 5580 6588 5598
rect 6570 5598 6588 5616
rect 6570 5616 6588 5634
rect 6570 5634 6588 5652
rect 6570 5652 6588 5670
rect 6570 5670 6588 5688
rect 6570 5688 6588 5706
rect 6570 5706 6588 5724
rect 6570 5724 6588 5742
rect 6570 5742 6588 5760
rect 6570 5760 6588 5778
rect 6570 5778 6588 5796
rect 6570 5796 6588 5814
rect 6570 5814 6588 5832
rect 6570 5832 6588 5850
rect 6570 5850 6588 5868
rect 6570 5868 6588 5886
rect 6570 5886 6588 5904
rect 6570 6768 6588 6786
rect 6570 6786 6588 6804
rect 6570 6804 6588 6822
rect 6570 6822 6588 6840
rect 6570 6840 6588 6858
rect 6570 6858 6588 6876
rect 6570 6876 6588 6894
rect 6570 6894 6588 6912
rect 6570 6912 6588 6930
rect 6570 6930 6588 6948
rect 6570 6948 6588 6966
rect 6570 6966 6588 6984
rect 6570 6984 6588 7002
rect 6570 7002 6588 7020
rect 6570 7020 6588 7038
rect 6570 7038 6588 7056
rect 6570 7056 6588 7074
rect 6570 7074 6588 7092
rect 6570 7092 6588 7110
rect 6570 7110 6588 7128
rect 6570 7128 6588 7146
rect 6570 7146 6588 7164
rect 6570 7164 6588 7182
rect 6570 7182 6588 7200
rect 6570 7200 6588 7218
rect 6570 7218 6588 7236
rect 6570 7236 6588 7254
rect 6570 7254 6588 7272
rect 6570 7272 6588 7290
rect 6570 7290 6588 7308
rect 6570 7308 6588 7326
rect 6570 7326 6588 7344
rect 6570 7344 6588 7362
rect 6570 7362 6588 7380
rect 6570 7380 6588 7398
rect 6570 7398 6588 7416
rect 6570 7416 6588 7434
rect 6570 7434 6588 7452
rect 6570 7452 6588 7470
rect 6570 7470 6588 7488
rect 6570 7488 6588 7506
rect 6570 7506 6588 7524
rect 6570 7524 6588 7542
rect 6570 7542 6588 7560
rect 6570 7560 6588 7578
rect 6570 7578 6588 7596
rect 6570 7596 6588 7614
rect 6570 7614 6588 7632
rect 6570 7632 6588 7650
rect 6570 7650 6588 7668
rect 6570 7668 6588 7686
rect 6570 7686 6588 7704
rect 6570 7704 6588 7722
rect 6570 7722 6588 7740
rect 6570 7740 6588 7758
rect 6570 7758 6588 7776
rect 6570 7776 6588 7794
rect 6570 7794 6588 7812
rect 6570 7812 6588 7830
rect 6570 7830 6588 7848
rect 6570 7848 6588 7866
rect 6570 7866 6588 7884
rect 6570 7884 6588 7902
rect 6570 7902 6588 7920
rect 6570 7920 6588 7938
rect 6570 7938 6588 7956
rect 6570 7956 6588 7974
rect 6570 7974 6588 7992
rect 6570 7992 6588 8010
rect 6570 8010 6588 8028
rect 6570 8028 6588 8046
rect 6570 8046 6588 8064
rect 6570 8064 6588 8082
rect 6570 8082 6588 8100
rect 6570 8100 6588 8118
rect 6570 8118 6588 8136
rect 6570 8136 6588 8154
rect 6570 8154 6588 8172
rect 6570 8172 6588 8190
rect 6570 8190 6588 8208
rect 6570 8208 6588 8226
rect 6570 8226 6588 8244
rect 6570 8244 6588 8262
rect 6570 8262 6588 8280
rect 6570 8280 6588 8298
rect 6570 8298 6588 8316
rect 6570 8316 6588 8334
rect 6570 8334 6588 8352
rect 6570 8352 6588 8370
rect 6570 8370 6588 8388
rect 6570 8388 6588 8406
rect 6570 8406 6588 8424
rect 6570 8424 6588 8442
rect 6570 8442 6588 8460
rect 6570 8460 6588 8478
rect 6570 8478 6588 8496
rect 6570 8496 6588 8514
rect 6570 8514 6588 8532
rect 6570 8532 6588 8550
rect 6570 8550 6588 8568
rect 6570 8568 6588 8586
rect 6570 8586 6588 8604
rect 6570 8604 6588 8622
rect 6570 8622 6588 8640
rect 6570 8640 6588 8658
rect 6570 8658 6588 8676
rect 6570 8676 6588 8694
rect 6570 8694 6588 8712
rect 6570 8712 6588 8730
rect 6570 8730 6588 8748
rect 6570 8748 6588 8766
rect 6570 8766 6588 8784
rect 6570 8784 6588 8802
rect 6570 8802 6588 8820
rect 6570 8820 6588 8838
rect 6570 8838 6588 8856
rect 6570 8856 6588 8874
rect 6570 8874 6588 8892
rect 6570 8892 6588 8910
rect 6570 8910 6588 8928
rect 6570 8928 6588 8946
rect 6570 8946 6588 8964
rect 6570 8964 6588 8982
rect 6570 8982 6588 9000
rect 6570 9000 6588 9018
rect 6570 9018 6588 9036
rect 6570 9036 6588 9054
rect 6570 9054 6588 9072
rect 6570 9072 6588 9090
rect 6570 9090 6588 9108
rect 6570 9108 6588 9126
rect 6570 9126 6588 9144
rect 6570 9144 6588 9162
rect 6570 9162 6588 9180
rect 6570 9180 6588 9198
rect 6570 9198 6588 9216
rect 6570 9216 6588 9234
rect 6570 9234 6588 9252
rect 6570 9252 6588 9270
rect 6570 9270 6588 9288
rect 6570 9288 6588 9306
rect 6570 9306 6588 9324
rect 6570 9324 6588 9342
rect 6570 9342 6588 9360
rect 6570 9360 6588 9378
rect 6570 9378 6588 9396
rect 6570 9396 6588 9414
rect 6570 9414 6588 9432
rect 6570 9432 6588 9450
rect 6570 9450 6588 9468
rect 6570 9468 6588 9486
rect 6570 9486 6588 9504
rect 6570 9504 6588 9522
rect 6570 9522 6588 9540
rect 6570 9540 6588 9558
rect 6570 9558 6588 9576
rect 6570 9576 6588 9594
rect 6570 9594 6588 9612
rect 6570 9612 6588 9630
rect 6570 9630 6588 9648
rect 6570 9648 6588 9666
rect 6570 9666 6588 9684
rect 6570 9684 6588 9702
rect 6570 9702 6588 9720
rect 6570 9720 6588 9738
rect 6570 9738 6588 9756
rect 6570 9756 6588 9774
rect 6570 9774 6588 9792
rect 6570 9792 6588 9810
rect 6570 9810 6588 9828
rect 6570 9828 6588 9846
rect 6570 9846 6588 9864
rect 6570 9864 6588 9882
rect 6570 9882 6588 9900
rect 6570 9900 6588 9918
rect 6570 9918 6588 9936
rect 6570 9936 6588 9954
rect 6588 1548 6606 1566
rect 6588 1566 6606 1584
rect 6588 1584 6606 1602
rect 6588 1602 6606 1620
rect 6588 1620 6606 1638
rect 6588 1638 6606 1656
rect 6588 1656 6606 1674
rect 6588 1674 6606 1692
rect 6588 1692 6606 1710
rect 6588 1710 6606 1728
rect 6588 1728 6606 1746
rect 6588 1746 6606 1764
rect 6588 1764 6606 1782
rect 6588 1782 6606 1800
rect 6588 1800 6606 1818
rect 6588 1818 6606 1836
rect 6588 1836 6606 1854
rect 6588 1854 6606 1872
rect 6588 1872 6606 1890
rect 6588 1890 6606 1908
rect 6588 1908 6606 1926
rect 6588 1926 6606 1944
rect 6588 1944 6606 1962
rect 6588 1962 6606 1980
rect 6588 1980 6606 1998
rect 6588 1998 6606 2016
rect 6588 2016 6606 2034
rect 6588 2034 6606 2052
rect 6588 2052 6606 2070
rect 6588 2070 6606 2088
rect 6588 2088 6606 2106
rect 6588 2106 6606 2124
rect 6588 2124 6606 2142
rect 6588 2142 6606 2160
rect 6588 2160 6606 2178
rect 6588 2178 6606 2196
rect 6588 2196 6606 2214
rect 6588 2214 6606 2232
rect 6588 2232 6606 2250
rect 6588 2250 6606 2268
rect 6588 2268 6606 2286
rect 6588 2286 6606 2304
rect 6588 2304 6606 2322
rect 6588 2322 6606 2340
rect 6588 2340 6606 2358
rect 6588 2358 6606 2376
rect 6588 2376 6606 2394
rect 6588 2394 6606 2412
rect 6588 2412 6606 2430
rect 6588 2430 6606 2448
rect 6588 2448 6606 2466
rect 6588 2466 6606 2484
rect 6588 2484 6606 2502
rect 6588 2502 6606 2520
rect 6588 2520 6606 2538
rect 6588 2538 6606 2556
rect 6588 2556 6606 2574
rect 6588 2574 6606 2592
rect 6588 2592 6606 2610
rect 6588 2610 6606 2628
rect 6588 2628 6606 2646
rect 6588 2646 6606 2664
rect 6588 2664 6606 2682
rect 6588 2682 6606 2700
rect 6588 2700 6606 2718
rect 6588 2718 6606 2736
rect 6588 2736 6606 2754
rect 6588 2754 6606 2772
rect 6588 2772 6606 2790
rect 6588 2790 6606 2808
rect 6588 2808 6606 2826
rect 6588 2826 6606 2844
rect 6588 2844 6606 2862
rect 6588 2862 6606 2880
rect 6588 2880 6606 2898
rect 6588 2898 6606 2916
rect 6588 2916 6606 2934
rect 6588 2934 6606 2952
rect 6588 2952 6606 2970
rect 6588 3528 6606 3546
rect 6588 3546 6606 3564
rect 6588 3564 6606 3582
rect 6588 3582 6606 3600
rect 6588 3600 6606 3618
rect 6588 3618 6606 3636
rect 6588 3636 6606 3654
rect 6588 3654 6606 3672
rect 6588 3672 6606 3690
rect 6588 3690 6606 3708
rect 6588 3708 6606 3726
rect 6588 3726 6606 3744
rect 6588 3744 6606 3762
rect 6588 3762 6606 3780
rect 6588 3780 6606 3798
rect 6588 3798 6606 3816
rect 6588 3816 6606 3834
rect 6588 3834 6606 3852
rect 6588 3852 6606 3870
rect 6588 3870 6606 3888
rect 6588 3888 6606 3906
rect 6588 3906 6606 3924
rect 6588 3924 6606 3942
rect 6588 3942 6606 3960
rect 6588 3960 6606 3978
rect 6588 3978 6606 3996
rect 6588 3996 6606 4014
rect 6588 4014 6606 4032
rect 6588 4032 6606 4050
rect 6588 4050 6606 4068
rect 6588 4068 6606 4086
rect 6588 4086 6606 4104
rect 6588 4104 6606 4122
rect 6588 4122 6606 4140
rect 6588 4140 6606 4158
rect 6588 4158 6606 4176
rect 6588 4176 6606 4194
rect 6588 4194 6606 4212
rect 6588 4212 6606 4230
rect 6588 4230 6606 4248
rect 6588 4248 6606 4266
rect 6588 4266 6606 4284
rect 6588 4284 6606 4302
rect 6588 4302 6606 4320
rect 6588 4320 6606 4338
rect 6588 4338 6606 4356
rect 6588 4356 6606 4374
rect 6588 4374 6606 4392
rect 6588 4392 6606 4410
rect 6588 4410 6606 4428
rect 6588 4428 6606 4446
rect 6588 4446 6606 4464
rect 6588 4464 6606 4482
rect 6588 4482 6606 4500
rect 6588 4500 6606 4518
rect 6588 4518 6606 4536
rect 6588 4536 6606 4554
rect 6588 4554 6606 4572
rect 6588 4572 6606 4590
rect 6588 4590 6606 4608
rect 6588 4608 6606 4626
rect 6588 4626 6606 4644
rect 6588 4644 6606 4662
rect 6588 4662 6606 4680
rect 6588 4680 6606 4698
rect 6588 4698 6606 4716
rect 6588 4716 6606 4734
rect 6588 4734 6606 4752
rect 6588 4752 6606 4770
rect 6588 4770 6606 4788
rect 6588 4788 6606 4806
rect 6588 4806 6606 4824
rect 6588 4824 6606 4842
rect 6588 4842 6606 4860
rect 6588 4860 6606 4878
rect 6588 4878 6606 4896
rect 6588 4896 6606 4914
rect 6588 4914 6606 4932
rect 6588 4932 6606 4950
rect 6588 4950 6606 4968
rect 6588 4968 6606 4986
rect 6588 4986 6606 5004
rect 6588 5004 6606 5022
rect 6588 5022 6606 5040
rect 6588 5040 6606 5058
rect 6588 5058 6606 5076
rect 6588 5076 6606 5094
rect 6588 5094 6606 5112
rect 6588 5112 6606 5130
rect 6588 5130 6606 5148
rect 6588 5148 6606 5166
rect 6588 5166 6606 5184
rect 6588 5184 6606 5202
rect 6588 5202 6606 5220
rect 6588 5220 6606 5238
rect 6588 5238 6606 5256
rect 6588 5256 6606 5274
rect 6588 5274 6606 5292
rect 6588 5292 6606 5310
rect 6588 5310 6606 5328
rect 6588 5328 6606 5346
rect 6588 5346 6606 5364
rect 6588 5364 6606 5382
rect 6588 5382 6606 5400
rect 6588 5400 6606 5418
rect 6588 5418 6606 5436
rect 6588 5436 6606 5454
rect 6588 5454 6606 5472
rect 6588 5472 6606 5490
rect 6588 5490 6606 5508
rect 6588 5508 6606 5526
rect 6588 5526 6606 5544
rect 6588 5544 6606 5562
rect 6588 5562 6606 5580
rect 6588 5580 6606 5598
rect 6588 5598 6606 5616
rect 6588 5616 6606 5634
rect 6588 5634 6606 5652
rect 6588 5652 6606 5670
rect 6588 5670 6606 5688
rect 6588 5688 6606 5706
rect 6588 5706 6606 5724
rect 6588 5724 6606 5742
rect 6588 5742 6606 5760
rect 6588 5760 6606 5778
rect 6588 5778 6606 5796
rect 6588 5796 6606 5814
rect 6588 5814 6606 5832
rect 6588 5832 6606 5850
rect 6588 5850 6606 5868
rect 6588 5868 6606 5886
rect 6588 5886 6606 5904
rect 6588 5904 6606 5922
rect 6588 6804 6606 6822
rect 6588 6822 6606 6840
rect 6588 6840 6606 6858
rect 6588 6858 6606 6876
rect 6588 6876 6606 6894
rect 6588 6894 6606 6912
rect 6588 6912 6606 6930
rect 6588 6930 6606 6948
rect 6588 6948 6606 6966
rect 6588 6966 6606 6984
rect 6588 6984 6606 7002
rect 6588 7002 6606 7020
rect 6588 7020 6606 7038
rect 6588 7038 6606 7056
rect 6588 7056 6606 7074
rect 6588 7074 6606 7092
rect 6588 7092 6606 7110
rect 6588 7110 6606 7128
rect 6588 7128 6606 7146
rect 6588 7146 6606 7164
rect 6588 7164 6606 7182
rect 6588 7182 6606 7200
rect 6588 7200 6606 7218
rect 6588 7218 6606 7236
rect 6588 7236 6606 7254
rect 6588 7254 6606 7272
rect 6588 7272 6606 7290
rect 6588 7290 6606 7308
rect 6588 7308 6606 7326
rect 6588 7326 6606 7344
rect 6588 7344 6606 7362
rect 6588 7362 6606 7380
rect 6588 7380 6606 7398
rect 6588 7398 6606 7416
rect 6588 7416 6606 7434
rect 6588 7434 6606 7452
rect 6588 7452 6606 7470
rect 6588 7470 6606 7488
rect 6588 7488 6606 7506
rect 6588 7506 6606 7524
rect 6588 7524 6606 7542
rect 6588 7542 6606 7560
rect 6588 7560 6606 7578
rect 6588 7578 6606 7596
rect 6588 7596 6606 7614
rect 6588 7614 6606 7632
rect 6588 7632 6606 7650
rect 6588 7650 6606 7668
rect 6588 7668 6606 7686
rect 6588 7686 6606 7704
rect 6588 7704 6606 7722
rect 6588 7722 6606 7740
rect 6588 7740 6606 7758
rect 6588 7758 6606 7776
rect 6588 7776 6606 7794
rect 6588 7794 6606 7812
rect 6588 7812 6606 7830
rect 6588 7830 6606 7848
rect 6588 7848 6606 7866
rect 6588 7866 6606 7884
rect 6588 7884 6606 7902
rect 6588 7902 6606 7920
rect 6588 7920 6606 7938
rect 6588 7938 6606 7956
rect 6588 7956 6606 7974
rect 6588 7974 6606 7992
rect 6588 7992 6606 8010
rect 6588 8010 6606 8028
rect 6588 8028 6606 8046
rect 6588 8046 6606 8064
rect 6588 8064 6606 8082
rect 6588 8082 6606 8100
rect 6588 8100 6606 8118
rect 6588 8118 6606 8136
rect 6588 8136 6606 8154
rect 6588 8154 6606 8172
rect 6588 8172 6606 8190
rect 6588 8190 6606 8208
rect 6588 8208 6606 8226
rect 6588 8226 6606 8244
rect 6588 8244 6606 8262
rect 6588 8262 6606 8280
rect 6588 8280 6606 8298
rect 6588 8298 6606 8316
rect 6588 8316 6606 8334
rect 6588 8334 6606 8352
rect 6588 8352 6606 8370
rect 6588 8370 6606 8388
rect 6588 8388 6606 8406
rect 6588 8406 6606 8424
rect 6588 8424 6606 8442
rect 6588 8442 6606 8460
rect 6588 8460 6606 8478
rect 6588 8478 6606 8496
rect 6588 8496 6606 8514
rect 6588 8514 6606 8532
rect 6588 8532 6606 8550
rect 6588 8550 6606 8568
rect 6588 8568 6606 8586
rect 6588 8586 6606 8604
rect 6588 8604 6606 8622
rect 6588 8622 6606 8640
rect 6588 8640 6606 8658
rect 6588 8658 6606 8676
rect 6588 8676 6606 8694
rect 6588 8694 6606 8712
rect 6588 8712 6606 8730
rect 6588 8730 6606 8748
rect 6588 8748 6606 8766
rect 6588 8766 6606 8784
rect 6588 8784 6606 8802
rect 6588 8802 6606 8820
rect 6588 8820 6606 8838
rect 6588 8838 6606 8856
rect 6588 8856 6606 8874
rect 6588 8874 6606 8892
rect 6588 8892 6606 8910
rect 6588 8910 6606 8928
rect 6588 8928 6606 8946
rect 6588 8946 6606 8964
rect 6588 8964 6606 8982
rect 6588 8982 6606 9000
rect 6588 9000 6606 9018
rect 6588 9018 6606 9036
rect 6588 9036 6606 9054
rect 6588 9054 6606 9072
rect 6588 9072 6606 9090
rect 6588 9090 6606 9108
rect 6588 9108 6606 9126
rect 6588 9126 6606 9144
rect 6588 9144 6606 9162
rect 6588 9162 6606 9180
rect 6588 9180 6606 9198
rect 6588 9198 6606 9216
rect 6588 9216 6606 9234
rect 6588 9234 6606 9252
rect 6588 9252 6606 9270
rect 6588 9270 6606 9288
rect 6588 9288 6606 9306
rect 6588 9306 6606 9324
rect 6588 9324 6606 9342
rect 6588 9342 6606 9360
rect 6588 9360 6606 9378
rect 6588 9378 6606 9396
rect 6588 9396 6606 9414
rect 6588 9414 6606 9432
rect 6588 9432 6606 9450
rect 6588 9450 6606 9468
rect 6588 9468 6606 9486
rect 6588 9486 6606 9504
rect 6588 9504 6606 9522
rect 6588 9522 6606 9540
rect 6588 9540 6606 9558
rect 6588 9558 6606 9576
rect 6588 9576 6606 9594
rect 6588 9594 6606 9612
rect 6588 9612 6606 9630
rect 6588 9630 6606 9648
rect 6588 9648 6606 9666
rect 6588 9666 6606 9684
rect 6588 9684 6606 9702
rect 6588 9702 6606 9720
rect 6588 9720 6606 9738
rect 6588 9738 6606 9756
rect 6588 9756 6606 9774
rect 6588 9774 6606 9792
rect 6588 9792 6606 9810
rect 6588 9810 6606 9828
rect 6588 9828 6606 9846
rect 6588 9846 6606 9864
rect 6588 9864 6606 9882
rect 6588 9882 6606 9900
rect 6588 9900 6606 9918
rect 6588 9918 6606 9936
rect 6588 9936 6606 9954
rect 6588 9954 6606 9972
rect 6606 1548 6624 1566
rect 6606 1566 6624 1584
rect 6606 1584 6624 1602
rect 6606 1602 6624 1620
rect 6606 1620 6624 1638
rect 6606 1638 6624 1656
rect 6606 1656 6624 1674
rect 6606 1674 6624 1692
rect 6606 1692 6624 1710
rect 6606 1710 6624 1728
rect 6606 1728 6624 1746
rect 6606 1746 6624 1764
rect 6606 1764 6624 1782
rect 6606 1782 6624 1800
rect 6606 1800 6624 1818
rect 6606 1818 6624 1836
rect 6606 1836 6624 1854
rect 6606 1854 6624 1872
rect 6606 1872 6624 1890
rect 6606 1890 6624 1908
rect 6606 1908 6624 1926
rect 6606 1926 6624 1944
rect 6606 1944 6624 1962
rect 6606 1962 6624 1980
rect 6606 1980 6624 1998
rect 6606 1998 6624 2016
rect 6606 2016 6624 2034
rect 6606 2034 6624 2052
rect 6606 2052 6624 2070
rect 6606 2070 6624 2088
rect 6606 2088 6624 2106
rect 6606 2106 6624 2124
rect 6606 2124 6624 2142
rect 6606 2142 6624 2160
rect 6606 2160 6624 2178
rect 6606 2178 6624 2196
rect 6606 2196 6624 2214
rect 6606 2214 6624 2232
rect 6606 2232 6624 2250
rect 6606 2250 6624 2268
rect 6606 2268 6624 2286
rect 6606 2286 6624 2304
rect 6606 2304 6624 2322
rect 6606 2322 6624 2340
rect 6606 2340 6624 2358
rect 6606 2358 6624 2376
rect 6606 2376 6624 2394
rect 6606 2394 6624 2412
rect 6606 2412 6624 2430
rect 6606 2430 6624 2448
rect 6606 2448 6624 2466
rect 6606 2466 6624 2484
rect 6606 2484 6624 2502
rect 6606 2502 6624 2520
rect 6606 2520 6624 2538
rect 6606 2538 6624 2556
rect 6606 2556 6624 2574
rect 6606 2574 6624 2592
rect 6606 2592 6624 2610
rect 6606 2610 6624 2628
rect 6606 2628 6624 2646
rect 6606 2646 6624 2664
rect 6606 2664 6624 2682
rect 6606 2682 6624 2700
rect 6606 2700 6624 2718
rect 6606 2718 6624 2736
rect 6606 2736 6624 2754
rect 6606 2754 6624 2772
rect 6606 2772 6624 2790
rect 6606 2790 6624 2808
rect 6606 2808 6624 2826
rect 6606 2826 6624 2844
rect 6606 2844 6624 2862
rect 6606 2862 6624 2880
rect 6606 2880 6624 2898
rect 6606 2898 6624 2916
rect 6606 2916 6624 2934
rect 6606 2934 6624 2952
rect 6606 2952 6624 2970
rect 6606 3132 6624 3150
rect 6606 3546 6624 3564
rect 6606 3564 6624 3582
rect 6606 3582 6624 3600
rect 6606 3600 6624 3618
rect 6606 3618 6624 3636
rect 6606 3636 6624 3654
rect 6606 3654 6624 3672
rect 6606 3672 6624 3690
rect 6606 3690 6624 3708
rect 6606 3708 6624 3726
rect 6606 3726 6624 3744
rect 6606 3744 6624 3762
rect 6606 3762 6624 3780
rect 6606 3780 6624 3798
rect 6606 3798 6624 3816
rect 6606 3816 6624 3834
rect 6606 3834 6624 3852
rect 6606 3852 6624 3870
rect 6606 3870 6624 3888
rect 6606 3888 6624 3906
rect 6606 3906 6624 3924
rect 6606 3924 6624 3942
rect 6606 3942 6624 3960
rect 6606 3960 6624 3978
rect 6606 3978 6624 3996
rect 6606 3996 6624 4014
rect 6606 4014 6624 4032
rect 6606 4032 6624 4050
rect 6606 4050 6624 4068
rect 6606 4068 6624 4086
rect 6606 4086 6624 4104
rect 6606 4104 6624 4122
rect 6606 4122 6624 4140
rect 6606 4140 6624 4158
rect 6606 4158 6624 4176
rect 6606 4176 6624 4194
rect 6606 4194 6624 4212
rect 6606 4212 6624 4230
rect 6606 4230 6624 4248
rect 6606 4248 6624 4266
rect 6606 4266 6624 4284
rect 6606 4284 6624 4302
rect 6606 4302 6624 4320
rect 6606 4320 6624 4338
rect 6606 4338 6624 4356
rect 6606 4356 6624 4374
rect 6606 4374 6624 4392
rect 6606 4392 6624 4410
rect 6606 4410 6624 4428
rect 6606 4428 6624 4446
rect 6606 4446 6624 4464
rect 6606 4464 6624 4482
rect 6606 4482 6624 4500
rect 6606 4500 6624 4518
rect 6606 4518 6624 4536
rect 6606 4536 6624 4554
rect 6606 4554 6624 4572
rect 6606 4572 6624 4590
rect 6606 4590 6624 4608
rect 6606 4608 6624 4626
rect 6606 4626 6624 4644
rect 6606 4644 6624 4662
rect 6606 4662 6624 4680
rect 6606 4680 6624 4698
rect 6606 4698 6624 4716
rect 6606 4716 6624 4734
rect 6606 4734 6624 4752
rect 6606 4752 6624 4770
rect 6606 4770 6624 4788
rect 6606 4788 6624 4806
rect 6606 4806 6624 4824
rect 6606 4824 6624 4842
rect 6606 4842 6624 4860
rect 6606 4860 6624 4878
rect 6606 4878 6624 4896
rect 6606 4896 6624 4914
rect 6606 4914 6624 4932
rect 6606 4932 6624 4950
rect 6606 4950 6624 4968
rect 6606 4968 6624 4986
rect 6606 4986 6624 5004
rect 6606 5004 6624 5022
rect 6606 5022 6624 5040
rect 6606 5040 6624 5058
rect 6606 5058 6624 5076
rect 6606 5076 6624 5094
rect 6606 5094 6624 5112
rect 6606 5112 6624 5130
rect 6606 5130 6624 5148
rect 6606 5148 6624 5166
rect 6606 5166 6624 5184
rect 6606 5184 6624 5202
rect 6606 5202 6624 5220
rect 6606 5220 6624 5238
rect 6606 5238 6624 5256
rect 6606 5256 6624 5274
rect 6606 5274 6624 5292
rect 6606 5292 6624 5310
rect 6606 5310 6624 5328
rect 6606 5328 6624 5346
rect 6606 5346 6624 5364
rect 6606 5364 6624 5382
rect 6606 5382 6624 5400
rect 6606 5400 6624 5418
rect 6606 5418 6624 5436
rect 6606 5436 6624 5454
rect 6606 5454 6624 5472
rect 6606 5472 6624 5490
rect 6606 5490 6624 5508
rect 6606 5508 6624 5526
rect 6606 5526 6624 5544
rect 6606 5544 6624 5562
rect 6606 5562 6624 5580
rect 6606 5580 6624 5598
rect 6606 5598 6624 5616
rect 6606 5616 6624 5634
rect 6606 5634 6624 5652
rect 6606 5652 6624 5670
rect 6606 5670 6624 5688
rect 6606 5688 6624 5706
rect 6606 5706 6624 5724
rect 6606 5724 6624 5742
rect 6606 5742 6624 5760
rect 6606 5760 6624 5778
rect 6606 5778 6624 5796
rect 6606 5796 6624 5814
rect 6606 5814 6624 5832
rect 6606 5832 6624 5850
rect 6606 5850 6624 5868
rect 6606 5868 6624 5886
rect 6606 5886 6624 5904
rect 6606 5904 6624 5922
rect 6606 5922 6624 5940
rect 6606 6840 6624 6858
rect 6606 6858 6624 6876
rect 6606 6876 6624 6894
rect 6606 6894 6624 6912
rect 6606 6912 6624 6930
rect 6606 6930 6624 6948
rect 6606 6948 6624 6966
rect 6606 6966 6624 6984
rect 6606 6984 6624 7002
rect 6606 7002 6624 7020
rect 6606 7020 6624 7038
rect 6606 7038 6624 7056
rect 6606 7056 6624 7074
rect 6606 7074 6624 7092
rect 6606 7092 6624 7110
rect 6606 7110 6624 7128
rect 6606 7128 6624 7146
rect 6606 7146 6624 7164
rect 6606 7164 6624 7182
rect 6606 7182 6624 7200
rect 6606 7200 6624 7218
rect 6606 7218 6624 7236
rect 6606 7236 6624 7254
rect 6606 7254 6624 7272
rect 6606 7272 6624 7290
rect 6606 7290 6624 7308
rect 6606 7308 6624 7326
rect 6606 7326 6624 7344
rect 6606 7344 6624 7362
rect 6606 7362 6624 7380
rect 6606 7380 6624 7398
rect 6606 7398 6624 7416
rect 6606 7416 6624 7434
rect 6606 7434 6624 7452
rect 6606 7452 6624 7470
rect 6606 7470 6624 7488
rect 6606 7488 6624 7506
rect 6606 7506 6624 7524
rect 6606 7524 6624 7542
rect 6606 7542 6624 7560
rect 6606 7560 6624 7578
rect 6606 7578 6624 7596
rect 6606 7596 6624 7614
rect 6606 7614 6624 7632
rect 6606 7632 6624 7650
rect 6606 7650 6624 7668
rect 6606 7668 6624 7686
rect 6606 7686 6624 7704
rect 6606 7704 6624 7722
rect 6606 7722 6624 7740
rect 6606 7740 6624 7758
rect 6606 7758 6624 7776
rect 6606 7776 6624 7794
rect 6606 7794 6624 7812
rect 6606 7812 6624 7830
rect 6606 7830 6624 7848
rect 6606 7848 6624 7866
rect 6606 7866 6624 7884
rect 6606 7884 6624 7902
rect 6606 7902 6624 7920
rect 6606 7920 6624 7938
rect 6606 7938 6624 7956
rect 6606 7956 6624 7974
rect 6606 7974 6624 7992
rect 6606 7992 6624 8010
rect 6606 8010 6624 8028
rect 6606 8028 6624 8046
rect 6606 8046 6624 8064
rect 6606 8064 6624 8082
rect 6606 8082 6624 8100
rect 6606 8100 6624 8118
rect 6606 8118 6624 8136
rect 6606 8136 6624 8154
rect 6606 8154 6624 8172
rect 6606 8172 6624 8190
rect 6606 8190 6624 8208
rect 6606 8208 6624 8226
rect 6606 8226 6624 8244
rect 6606 8244 6624 8262
rect 6606 8262 6624 8280
rect 6606 8280 6624 8298
rect 6606 8298 6624 8316
rect 6606 8316 6624 8334
rect 6606 8334 6624 8352
rect 6606 8352 6624 8370
rect 6606 8370 6624 8388
rect 6606 8388 6624 8406
rect 6606 8406 6624 8424
rect 6606 8424 6624 8442
rect 6606 8442 6624 8460
rect 6606 8460 6624 8478
rect 6606 8478 6624 8496
rect 6606 8496 6624 8514
rect 6606 8514 6624 8532
rect 6606 8532 6624 8550
rect 6606 8550 6624 8568
rect 6606 8568 6624 8586
rect 6606 8586 6624 8604
rect 6606 8604 6624 8622
rect 6606 8622 6624 8640
rect 6606 8640 6624 8658
rect 6606 8658 6624 8676
rect 6606 8676 6624 8694
rect 6606 8694 6624 8712
rect 6606 8712 6624 8730
rect 6606 8730 6624 8748
rect 6606 8748 6624 8766
rect 6606 8766 6624 8784
rect 6606 8784 6624 8802
rect 6606 8802 6624 8820
rect 6606 8820 6624 8838
rect 6606 8838 6624 8856
rect 6606 8856 6624 8874
rect 6606 8874 6624 8892
rect 6606 8892 6624 8910
rect 6606 8910 6624 8928
rect 6606 8928 6624 8946
rect 6606 8946 6624 8964
rect 6606 8964 6624 8982
rect 6606 8982 6624 9000
rect 6606 9000 6624 9018
rect 6606 9018 6624 9036
rect 6606 9036 6624 9054
rect 6606 9054 6624 9072
rect 6606 9072 6624 9090
rect 6606 9090 6624 9108
rect 6606 9108 6624 9126
rect 6606 9126 6624 9144
rect 6606 9144 6624 9162
rect 6606 9162 6624 9180
rect 6606 9180 6624 9198
rect 6606 9198 6624 9216
rect 6606 9216 6624 9234
rect 6606 9234 6624 9252
rect 6606 9252 6624 9270
rect 6606 9270 6624 9288
rect 6606 9288 6624 9306
rect 6606 9306 6624 9324
rect 6606 9324 6624 9342
rect 6606 9342 6624 9360
rect 6606 9360 6624 9378
rect 6606 9378 6624 9396
rect 6606 9396 6624 9414
rect 6606 9414 6624 9432
rect 6606 9432 6624 9450
rect 6606 9450 6624 9468
rect 6606 9468 6624 9486
rect 6606 9486 6624 9504
rect 6606 9504 6624 9522
rect 6606 9522 6624 9540
rect 6606 9540 6624 9558
rect 6606 9558 6624 9576
rect 6606 9576 6624 9594
rect 6606 9594 6624 9612
rect 6606 9612 6624 9630
rect 6606 9630 6624 9648
rect 6606 9648 6624 9666
rect 6606 9666 6624 9684
rect 6606 9684 6624 9702
rect 6606 9702 6624 9720
rect 6606 9720 6624 9738
rect 6606 9738 6624 9756
rect 6606 9756 6624 9774
rect 6606 9774 6624 9792
rect 6606 9792 6624 9810
rect 6606 9810 6624 9828
rect 6606 9828 6624 9846
rect 6606 9846 6624 9864
rect 6606 9864 6624 9882
rect 6606 9882 6624 9900
rect 6606 9900 6624 9918
rect 6606 9918 6624 9936
rect 6606 9936 6624 9954
rect 6606 9954 6624 9972
rect 6606 9972 6624 9990
rect 6624 1566 6642 1584
rect 6624 1584 6642 1602
rect 6624 1602 6642 1620
rect 6624 1620 6642 1638
rect 6624 1638 6642 1656
rect 6624 1656 6642 1674
rect 6624 1674 6642 1692
rect 6624 1692 6642 1710
rect 6624 1710 6642 1728
rect 6624 1728 6642 1746
rect 6624 1746 6642 1764
rect 6624 1764 6642 1782
rect 6624 1782 6642 1800
rect 6624 1800 6642 1818
rect 6624 1818 6642 1836
rect 6624 1836 6642 1854
rect 6624 1854 6642 1872
rect 6624 1872 6642 1890
rect 6624 1890 6642 1908
rect 6624 1908 6642 1926
rect 6624 1926 6642 1944
rect 6624 1944 6642 1962
rect 6624 1962 6642 1980
rect 6624 1980 6642 1998
rect 6624 1998 6642 2016
rect 6624 2016 6642 2034
rect 6624 2034 6642 2052
rect 6624 2052 6642 2070
rect 6624 2070 6642 2088
rect 6624 2088 6642 2106
rect 6624 2106 6642 2124
rect 6624 2124 6642 2142
rect 6624 2142 6642 2160
rect 6624 2160 6642 2178
rect 6624 2178 6642 2196
rect 6624 2196 6642 2214
rect 6624 2214 6642 2232
rect 6624 2232 6642 2250
rect 6624 2250 6642 2268
rect 6624 2268 6642 2286
rect 6624 2286 6642 2304
rect 6624 2304 6642 2322
rect 6624 2322 6642 2340
rect 6624 2340 6642 2358
rect 6624 2358 6642 2376
rect 6624 2376 6642 2394
rect 6624 2394 6642 2412
rect 6624 2412 6642 2430
rect 6624 2430 6642 2448
rect 6624 2448 6642 2466
rect 6624 2466 6642 2484
rect 6624 2484 6642 2502
rect 6624 2502 6642 2520
rect 6624 2520 6642 2538
rect 6624 2538 6642 2556
rect 6624 2556 6642 2574
rect 6624 2574 6642 2592
rect 6624 2592 6642 2610
rect 6624 2610 6642 2628
rect 6624 2628 6642 2646
rect 6624 2646 6642 2664
rect 6624 2664 6642 2682
rect 6624 2682 6642 2700
rect 6624 2700 6642 2718
rect 6624 2718 6642 2736
rect 6624 2736 6642 2754
rect 6624 2754 6642 2772
rect 6624 2772 6642 2790
rect 6624 2790 6642 2808
rect 6624 2808 6642 2826
rect 6624 2826 6642 2844
rect 6624 2844 6642 2862
rect 6624 2862 6642 2880
rect 6624 2880 6642 2898
rect 6624 2898 6642 2916
rect 6624 2916 6642 2934
rect 6624 2934 6642 2952
rect 6624 2952 6642 2970
rect 6624 3132 6642 3150
rect 6624 3150 6642 3168
rect 6624 3168 6642 3186
rect 6624 3186 6642 3204
rect 6624 3204 6642 3222
rect 6624 3222 6642 3240
rect 6624 3240 6642 3258
rect 6624 3258 6642 3276
rect 6624 3276 6642 3294
rect 6624 3294 6642 3312
rect 6624 3312 6642 3330
rect 6624 3330 6642 3348
rect 6624 3348 6642 3366
rect 6624 3366 6642 3384
rect 6624 3564 6642 3582
rect 6624 3582 6642 3600
rect 6624 3600 6642 3618
rect 6624 3618 6642 3636
rect 6624 3636 6642 3654
rect 6624 3654 6642 3672
rect 6624 3672 6642 3690
rect 6624 3690 6642 3708
rect 6624 3708 6642 3726
rect 6624 3726 6642 3744
rect 6624 3744 6642 3762
rect 6624 3762 6642 3780
rect 6624 3780 6642 3798
rect 6624 3798 6642 3816
rect 6624 3816 6642 3834
rect 6624 3834 6642 3852
rect 6624 3852 6642 3870
rect 6624 3870 6642 3888
rect 6624 3888 6642 3906
rect 6624 3906 6642 3924
rect 6624 3924 6642 3942
rect 6624 3942 6642 3960
rect 6624 3960 6642 3978
rect 6624 3978 6642 3996
rect 6624 3996 6642 4014
rect 6624 4014 6642 4032
rect 6624 4032 6642 4050
rect 6624 4050 6642 4068
rect 6624 4068 6642 4086
rect 6624 4086 6642 4104
rect 6624 4104 6642 4122
rect 6624 4122 6642 4140
rect 6624 4140 6642 4158
rect 6624 4158 6642 4176
rect 6624 4176 6642 4194
rect 6624 4194 6642 4212
rect 6624 4212 6642 4230
rect 6624 4230 6642 4248
rect 6624 4248 6642 4266
rect 6624 4266 6642 4284
rect 6624 4284 6642 4302
rect 6624 4302 6642 4320
rect 6624 4320 6642 4338
rect 6624 4338 6642 4356
rect 6624 4356 6642 4374
rect 6624 4374 6642 4392
rect 6624 4392 6642 4410
rect 6624 4410 6642 4428
rect 6624 4428 6642 4446
rect 6624 4446 6642 4464
rect 6624 4464 6642 4482
rect 6624 4482 6642 4500
rect 6624 4500 6642 4518
rect 6624 4518 6642 4536
rect 6624 4536 6642 4554
rect 6624 4554 6642 4572
rect 6624 4572 6642 4590
rect 6624 4590 6642 4608
rect 6624 4608 6642 4626
rect 6624 4626 6642 4644
rect 6624 4644 6642 4662
rect 6624 4662 6642 4680
rect 6624 4680 6642 4698
rect 6624 4698 6642 4716
rect 6624 4716 6642 4734
rect 6624 4734 6642 4752
rect 6624 4752 6642 4770
rect 6624 4770 6642 4788
rect 6624 4788 6642 4806
rect 6624 4806 6642 4824
rect 6624 4824 6642 4842
rect 6624 4842 6642 4860
rect 6624 4860 6642 4878
rect 6624 4878 6642 4896
rect 6624 4896 6642 4914
rect 6624 4914 6642 4932
rect 6624 4932 6642 4950
rect 6624 4950 6642 4968
rect 6624 4968 6642 4986
rect 6624 4986 6642 5004
rect 6624 5004 6642 5022
rect 6624 5022 6642 5040
rect 6624 5040 6642 5058
rect 6624 5058 6642 5076
rect 6624 5076 6642 5094
rect 6624 5094 6642 5112
rect 6624 5112 6642 5130
rect 6624 5130 6642 5148
rect 6624 5148 6642 5166
rect 6624 5166 6642 5184
rect 6624 5184 6642 5202
rect 6624 5202 6642 5220
rect 6624 5220 6642 5238
rect 6624 5238 6642 5256
rect 6624 5256 6642 5274
rect 6624 5274 6642 5292
rect 6624 5292 6642 5310
rect 6624 5310 6642 5328
rect 6624 5328 6642 5346
rect 6624 5346 6642 5364
rect 6624 5364 6642 5382
rect 6624 5382 6642 5400
rect 6624 5400 6642 5418
rect 6624 5418 6642 5436
rect 6624 5436 6642 5454
rect 6624 5454 6642 5472
rect 6624 5472 6642 5490
rect 6624 5490 6642 5508
rect 6624 5508 6642 5526
rect 6624 5526 6642 5544
rect 6624 5544 6642 5562
rect 6624 5562 6642 5580
rect 6624 5580 6642 5598
rect 6624 5598 6642 5616
rect 6624 5616 6642 5634
rect 6624 5634 6642 5652
rect 6624 5652 6642 5670
rect 6624 5670 6642 5688
rect 6624 5688 6642 5706
rect 6624 5706 6642 5724
rect 6624 5724 6642 5742
rect 6624 5742 6642 5760
rect 6624 5760 6642 5778
rect 6624 5778 6642 5796
rect 6624 5796 6642 5814
rect 6624 5814 6642 5832
rect 6624 5832 6642 5850
rect 6624 5850 6642 5868
rect 6624 5868 6642 5886
rect 6624 5886 6642 5904
rect 6624 5904 6642 5922
rect 6624 5922 6642 5940
rect 6624 6894 6642 6912
rect 6624 6912 6642 6930
rect 6624 6930 6642 6948
rect 6624 6948 6642 6966
rect 6624 6966 6642 6984
rect 6624 6984 6642 7002
rect 6624 7002 6642 7020
rect 6624 7020 6642 7038
rect 6624 7038 6642 7056
rect 6624 7056 6642 7074
rect 6624 7074 6642 7092
rect 6624 7092 6642 7110
rect 6624 7110 6642 7128
rect 6624 7128 6642 7146
rect 6624 7146 6642 7164
rect 6624 7164 6642 7182
rect 6624 7182 6642 7200
rect 6624 7200 6642 7218
rect 6624 7218 6642 7236
rect 6624 7236 6642 7254
rect 6624 7254 6642 7272
rect 6624 7272 6642 7290
rect 6624 7290 6642 7308
rect 6624 7308 6642 7326
rect 6624 7326 6642 7344
rect 6624 7344 6642 7362
rect 6624 7362 6642 7380
rect 6624 7380 6642 7398
rect 6624 7398 6642 7416
rect 6624 7416 6642 7434
rect 6624 7434 6642 7452
rect 6624 7452 6642 7470
rect 6624 7470 6642 7488
rect 6624 7488 6642 7506
rect 6624 7506 6642 7524
rect 6624 7524 6642 7542
rect 6624 7542 6642 7560
rect 6624 7560 6642 7578
rect 6624 7578 6642 7596
rect 6624 7596 6642 7614
rect 6624 7614 6642 7632
rect 6624 7632 6642 7650
rect 6624 7650 6642 7668
rect 6624 7668 6642 7686
rect 6624 7686 6642 7704
rect 6624 7704 6642 7722
rect 6624 7722 6642 7740
rect 6624 7740 6642 7758
rect 6624 7758 6642 7776
rect 6624 7776 6642 7794
rect 6624 7794 6642 7812
rect 6624 7812 6642 7830
rect 6624 7830 6642 7848
rect 6624 7848 6642 7866
rect 6624 7866 6642 7884
rect 6624 7884 6642 7902
rect 6624 7902 6642 7920
rect 6624 7920 6642 7938
rect 6624 7938 6642 7956
rect 6624 7956 6642 7974
rect 6624 7974 6642 7992
rect 6624 7992 6642 8010
rect 6624 8010 6642 8028
rect 6624 8028 6642 8046
rect 6624 8046 6642 8064
rect 6624 8064 6642 8082
rect 6624 8082 6642 8100
rect 6624 8100 6642 8118
rect 6624 8118 6642 8136
rect 6624 8136 6642 8154
rect 6624 8154 6642 8172
rect 6624 8172 6642 8190
rect 6624 8190 6642 8208
rect 6624 8208 6642 8226
rect 6624 8226 6642 8244
rect 6624 8244 6642 8262
rect 6624 8262 6642 8280
rect 6624 8280 6642 8298
rect 6624 8298 6642 8316
rect 6624 8316 6642 8334
rect 6624 8334 6642 8352
rect 6624 8352 6642 8370
rect 6624 8370 6642 8388
rect 6624 8388 6642 8406
rect 6624 8406 6642 8424
rect 6624 8424 6642 8442
rect 6624 8442 6642 8460
rect 6624 8460 6642 8478
rect 6624 8478 6642 8496
rect 6624 8496 6642 8514
rect 6624 8514 6642 8532
rect 6624 8532 6642 8550
rect 6624 8550 6642 8568
rect 6624 8568 6642 8586
rect 6624 8586 6642 8604
rect 6624 8604 6642 8622
rect 6624 8622 6642 8640
rect 6624 8640 6642 8658
rect 6624 8658 6642 8676
rect 6624 8676 6642 8694
rect 6624 8694 6642 8712
rect 6624 8712 6642 8730
rect 6624 8730 6642 8748
rect 6624 8748 6642 8766
rect 6624 8766 6642 8784
rect 6624 8784 6642 8802
rect 6624 8802 6642 8820
rect 6624 8820 6642 8838
rect 6624 8838 6642 8856
rect 6624 8856 6642 8874
rect 6624 8874 6642 8892
rect 6624 8892 6642 8910
rect 6624 8910 6642 8928
rect 6624 8928 6642 8946
rect 6624 8946 6642 8964
rect 6624 8964 6642 8982
rect 6624 8982 6642 9000
rect 6624 9000 6642 9018
rect 6624 9018 6642 9036
rect 6624 9036 6642 9054
rect 6624 9054 6642 9072
rect 6624 9072 6642 9090
rect 6624 9090 6642 9108
rect 6624 9108 6642 9126
rect 6624 9126 6642 9144
rect 6624 9144 6642 9162
rect 6624 9162 6642 9180
rect 6624 9180 6642 9198
rect 6624 9198 6642 9216
rect 6624 9216 6642 9234
rect 6624 9234 6642 9252
rect 6624 9252 6642 9270
rect 6624 9270 6642 9288
rect 6624 9288 6642 9306
rect 6624 9306 6642 9324
rect 6624 9324 6642 9342
rect 6624 9342 6642 9360
rect 6624 9360 6642 9378
rect 6624 9378 6642 9396
rect 6624 9396 6642 9414
rect 6624 9414 6642 9432
rect 6624 9432 6642 9450
rect 6624 9450 6642 9468
rect 6624 9468 6642 9486
rect 6624 9486 6642 9504
rect 6624 9504 6642 9522
rect 6624 9522 6642 9540
rect 6624 9540 6642 9558
rect 6624 9558 6642 9576
rect 6624 9576 6642 9594
rect 6624 9594 6642 9612
rect 6624 9612 6642 9630
rect 6624 9630 6642 9648
rect 6624 9648 6642 9666
rect 6624 9666 6642 9684
rect 6624 9684 6642 9702
rect 6624 9702 6642 9720
rect 6624 9720 6642 9738
rect 6624 9738 6642 9756
rect 6624 9756 6642 9774
rect 6624 9774 6642 9792
rect 6624 9792 6642 9810
rect 6624 9810 6642 9828
rect 6624 9828 6642 9846
rect 6624 9846 6642 9864
rect 6624 9864 6642 9882
rect 6624 9882 6642 9900
rect 6624 9900 6642 9918
rect 6624 9918 6642 9936
rect 6624 9936 6642 9954
rect 6624 9954 6642 9972
rect 6624 9972 6642 9990
rect 6624 9990 6642 10008
rect 6624 10008 6642 10026
rect 6642 1566 6660 1584
rect 6642 1584 6660 1602
rect 6642 1602 6660 1620
rect 6642 1620 6660 1638
rect 6642 1638 6660 1656
rect 6642 1656 6660 1674
rect 6642 1674 6660 1692
rect 6642 1692 6660 1710
rect 6642 1710 6660 1728
rect 6642 1728 6660 1746
rect 6642 1746 6660 1764
rect 6642 1764 6660 1782
rect 6642 1782 6660 1800
rect 6642 1800 6660 1818
rect 6642 1818 6660 1836
rect 6642 1836 6660 1854
rect 6642 1854 6660 1872
rect 6642 1872 6660 1890
rect 6642 1890 6660 1908
rect 6642 1908 6660 1926
rect 6642 1926 6660 1944
rect 6642 1944 6660 1962
rect 6642 1962 6660 1980
rect 6642 1980 6660 1998
rect 6642 1998 6660 2016
rect 6642 2016 6660 2034
rect 6642 2034 6660 2052
rect 6642 2052 6660 2070
rect 6642 2070 6660 2088
rect 6642 2088 6660 2106
rect 6642 2106 6660 2124
rect 6642 2124 6660 2142
rect 6642 2142 6660 2160
rect 6642 2160 6660 2178
rect 6642 2178 6660 2196
rect 6642 2196 6660 2214
rect 6642 2214 6660 2232
rect 6642 2232 6660 2250
rect 6642 2250 6660 2268
rect 6642 2268 6660 2286
rect 6642 2286 6660 2304
rect 6642 2304 6660 2322
rect 6642 2322 6660 2340
rect 6642 2340 6660 2358
rect 6642 2358 6660 2376
rect 6642 2376 6660 2394
rect 6642 2394 6660 2412
rect 6642 2412 6660 2430
rect 6642 2430 6660 2448
rect 6642 2448 6660 2466
rect 6642 2466 6660 2484
rect 6642 2484 6660 2502
rect 6642 2502 6660 2520
rect 6642 2520 6660 2538
rect 6642 2538 6660 2556
rect 6642 2556 6660 2574
rect 6642 2574 6660 2592
rect 6642 2592 6660 2610
rect 6642 2610 6660 2628
rect 6642 2628 6660 2646
rect 6642 2646 6660 2664
rect 6642 2664 6660 2682
rect 6642 2682 6660 2700
rect 6642 2700 6660 2718
rect 6642 2718 6660 2736
rect 6642 2736 6660 2754
rect 6642 2754 6660 2772
rect 6642 2772 6660 2790
rect 6642 2790 6660 2808
rect 6642 2808 6660 2826
rect 6642 2826 6660 2844
rect 6642 2844 6660 2862
rect 6642 2862 6660 2880
rect 6642 2880 6660 2898
rect 6642 2898 6660 2916
rect 6642 2916 6660 2934
rect 6642 2934 6660 2952
rect 6642 2952 6660 2970
rect 6642 2970 6660 2988
rect 6642 3150 6660 3168
rect 6642 3168 6660 3186
rect 6642 3186 6660 3204
rect 6642 3204 6660 3222
rect 6642 3222 6660 3240
rect 6642 3240 6660 3258
rect 6642 3258 6660 3276
rect 6642 3276 6660 3294
rect 6642 3294 6660 3312
rect 6642 3312 6660 3330
rect 6642 3330 6660 3348
rect 6642 3348 6660 3366
rect 6642 3366 6660 3384
rect 6642 3384 6660 3402
rect 6642 3582 6660 3600
rect 6642 3600 6660 3618
rect 6642 3618 6660 3636
rect 6642 3636 6660 3654
rect 6642 3654 6660 3672
rect 6642 3672 6660 3690
rect 6642 3690 6660 3708
rect 6642 3708 6660 3726
rect 6642 3726 6660 3744
rect 6642 3744 6660 3762
rect 6642 3762 6660 3780
rect 6642 3780 6660 3798
rect 6642 3798 6660 3816
rect 6642 3816 6660 3834
rect 6642 3834 6660 3852
rect 6642 3852 6660 3870
rect 6642 3870 6660 3888
rect 6642 3888 6660 3906
rect 6642 3906 6660 3924
rect 6642 3924 6660 3942
rect 6642 3942 6660 3960
rect 6642 3960 6660 3978
rect 6642 3978 6660 3996
rect 6642 3996 6660 4014
rect 6642 4014 6660 4032
rect 6642 4032 6660 4050
rect 6642 4050 6660 4068
rect 6642 4068 6660 4086
rect 6642 4086 6660 4104
rect 6642 4104 6660 4122
rect 6642 4122 6660 4140
rect 6642 4140 6660 4158
rect 6642 4158 6660 4176
rect 6642 4176 6660 4194
rect 6642 4194 6660 4212
rect 6642 4212 6660 4230
rect 6642 4230 6660 4248
rect 6642 4248 6660 4266
rect 6642 4266 6660 4284
rect 6642 4284 6660 4302
rect 6642 4302 6660 4320
rect 6642 4320 6660 4338
rect 6642 4338 6660 4356
rect 6642 4356 6660 4374
rect 6642 4374 6660 4392
rect 6642 4392 6660 4410
rect 6642 4410 6660 4428
rect 6642 4428 6660 4446
rect 6642 4446 6660 4464
rect 6642 4464 6660 4482
rect 6642 4482 6660 4500
rect 6642 4500 6660 4518
rect 6642 4518 6660 4536
rect 6642 4536 6660 4554
rect 6642 4554 6660 4572
rect 6642 4572 6660 4590
rect 6642 4590 6660 4608
rect 6642 4608 6660 4626
rect 6642 4626 6660 4644
rect 6642 4644 6660 4662
rect 6642 4662 6660 4680
rect 6642 4680 6660 4698
rect 6642 4698 6660 4716
rect 6642 4716 6660 4734
rect 6642 4734 6660 4752
rect 6642 4752 6660 4770
rect 6642 4770 6660 4788
rect 6642 4788 6660 4806
rect 6642 4806 6660 4824
rect 6642 4824 6660 4842
rect 6642 4842 6660 4860
rect 6642 4860 6660 4878
rect 6642 4878 6660 4896
rect 6642 4896 6660 4914
rect 6642 4914 6660 4932
rect 6642 4932 6660 4950
rect 6642 4950 6660 4968
rect 6642 4968 6660 4986
rect 6642 4986 6660 5004
rect 6642 5004 6660 5022
rect 6642 5022 6660 5040
rect 6642 5040 6660 5058
rect 6642 5058 6660 5076
rect 6642 5076 6660 5094
rect 6642 5094 6660 5112
rect 6642 5112 6660 5130
rect 6642 5130 6660 5148
rect 6642 5148 6660 5166
rect 6642 5166 6660 5184
rect 6642 5184 6660 5202
rect 6642 5202 6660 5220
rect 6642 5220 6660 5238
rect 6642 5238 6660 5256
rect 6642 5256 6660 5274
rect 6642 5274 6660 5292
rect 6642 5292 6660 5310
rect 6642 5310 6660 5328
rect 6642 5328 6660 5346
rect 6642 5346 6660 5364
rect 6642 5364 6660 5382
rect 6642 5382 6660 5400
rect 6642 5400 6660 5418
rect 6642 5418 6660 5436
rect 6642 5436 6660 5454
rect 6642 5454 6660 5472
rect 6642 5472 6660 5490
rect 6642 5490 6660 5508
rect 6642 5508 6660 5526
rect 6642 5526 6660 5544
rect 6642 5544 6660 5562
rect 6642 5562 6660 5580
rect 6642 5580 6660 5598
rect 6642 5598 6660 5616
rect 6642 5616 6660 5634
rect 6642 5634 6660 5652
rect 6642 5652 6660 5670
rect 6642 5670 6660 5688
rect 6642 5688 6660 5706
rect 6642 5706 6660 5724
rect 6642 5724 6660 5742
rect 6642 5742 6660 5760
rect 6642 5760 6660 5778
rect 6642 5778 6660 5796
rect 6642 5796 6660 5814
rect 6642 5814 6660 5832
rect 6642 5832 6660 5850
rect 6642 5850 6660 5868
rect 6642 5868 6660 5886
rect 6642 5886 6660 5904
rect 6642 5904 6660 5922
rect 6642 5922 6660 5940
rect 6642 5940 6660 5958
rect 6642 6930 6660 6948
rect 6642 6948 6660 6966
rect 6642 6966 6660 6984
rect 6642 6984 6660 7002
rect 6642 7002 6660 7020
rect 6642 7020 6660 7038
rect 6642 7038 6660 7056
rect 6642 7056 6660 7074
rect 6642 7074 6660 7092
rect 6642 7092 6660 7110
rect 6642 7110 6660 7128
rect 6642 7128 6660 7146
rect 6642 7146 6660 7164
rect 6642 7164 6660 7182
rect 6642 7182 6660 7200
rect 6642 7200 6660 7218
rect 6642 7218 6660 7236
rect 6642 7236 6660 7254
rect 6642 7254 6660 7272
rect 6642 7272 6660 7290
rect 6642 7290 6660 7308
rect 6642 7308 6660 7326
rect 6642 7326 6660 7344
rect 6642 7344 6660 7362
rect 6642 7362 6660 7380
rect 6642 7380 6660 7398
rect 6642 7398 6660 7416
rect 6642 7416 6660 7434
rect 6642 7434 6660 7452
rect 6642 7452 6660 7470
rect 6642 7470 6660 7488
rect 6642 7488 6660 7506
rect 6642 7506 6660 7524
rect 6642 7524 6660 7542
rect 6642 7542 6660 7560
rect 6642 7560 6660 7578
rect 6642 7578 6660 7596
rect 6642 7596 6660 7614
rect 6642 7614 6660 7632
rect 6642 7632 6660 7650
rect 6642 7650 6660 7668
rect 6642 7668 6660 7686
rect 6642 7686 6660 7704
rect 6642 7704 6660 7722
rect 6642 7722 6660 7740
rect 6642 7740 6660 7758
rect 6642 7758 6660 7776
rect 6642 7776 6660 7794
rect 6642 7794 6660 7812
rect 6642 7812 6660 7830
rect 6642 7830 6660 7848
rect 6642 7848 6660 7866
rect 6642 7866 6660 7884
rect 6642 7884 6660 7902
rect 6642 7902 6660 7920
rect 6642 7920 6660 7938
rect 6642 7938 6660 7956
rect 6642 7956 6660 7974
rect 6642 7974 6660 7992
rect 6642 7992 6660 8010
rect 6642 8010 6660 8028
rect 6642 8028 6660 8046
rect 6642 8046 6660 8064
rect 6642 8064 6660 8082
rect 6642 8082 6660 8100
rect 6642 8100 6660 8118
rect 6642 8118 6660 8136
rect 6642 8136 6660 8154
rect 6642 8154 6660 8172
rect 6642 8172 6660 8190
rect 6642 8190 6660 8208
rect 6642 8208 6660 8226
rect 6642 8226 6660 8244
rect 6642 8244 6660 8262
rect 6642 8262 6660 8280
rect 6642 8280 6660 8298
rect 6642 8298 6660 8316
rect 6642 8316 6660 8334
rect 6642 8334 6660 8352
rect 6642 8352 6660 8370
rect 6642 8370 6660 8388
rect 6642 8388 6660 8406
rect 6642 8406 6660 8424
rect 6642 8424 6660 8442
rect 6642 8442 6660 8460
rect 6642 8460 6660 8478
rect 6642 8478 6660 8496
rect 6642 8496 6660 8514
rect 6642 8514 6660 8532
rect 6642 8532 6660 8550
rect 6642 8550 6660 8568
rect 6642 8568 6660 8586
rect 6642 8586 6660 8604
rect 6642 8604 6660 8622
rect 6642 8622 6660 8640
rect 6642 8640 6660 8658
rect 6642 8658 6660 8676
rect 6642 8676 6660 8694
rect 6642 8694 6660 8712
rect 6642 8712 6660 8730
rect 6642 8730 6660 8748
rect 6642 8748 6660 8766
rect 6642 8766 6660 8784
rect 6642 8784 6660 8802
rect 6642 8802 6660 8820
rect 6642 8820 6660 8838
rect 6642 8838 6660 8856
rect 6642 8856 6660 8874
rect 6642 8874 6660 8892
rect 6642 8892 6660 8910
rect 6642 8910 6660 8928
rect 6642 8928 6660 8946
rect 6642 8946 6660 8964
rect 6642 8964 6660 8982
rect 6642 8982 6660 9000
rect 6642 9000 6660 9018
rect 6642 9018 6660 9036
rect 6642 9036 6660 9054
rect 6642 9054 6660 9072
rect 6642 9072 6660 9090
rect 6642 9090 6660 9108
rect 6642 9108 6660 9126
rect 6642 9126 6660 9144
rect 6642 9144 6660 9162
rect 6642 9162 6660 9180
rect 6642 9180 6660 9198
rect 6642 9198 6660 9216
rect 6642 9216 6660 9234
rect 6642 9234 6660 9252
rect 6642 9252 6660 9270
rect 6642 9270 6660 9288
rect 6642 9288 6660 9306
rect 6642 9306 6660 9324
rect 6642 9324 6660 9342
rect 6642 9342 6660 9360
rect 6642 9360 6660 9378
rect 6642 9378 6660 9396
rect 6642 9396 6660 9414
rect 6642 9414 6660 9432
rect 6642 9432 6660 9450
rect 6642 9450 6660 9468
rect 6642 9468 6660 9486
rect 6642 9486 6660 9504
rect 6642 9504 6660 9522
rect 6642 9522 6660 9540
rect 6642 9540 6660 9558
rect 6642 9558 6660 9576
rect 6642 9576 6660 9594
rect 6642 9594 6660 9612
rect 6642 9612 6660 9630
rect 6642 9630 6660 9648
rect 6642 9648 6660 9666
rect 6642 9666 6660 9684
rect 6642 9684 6660 9702
rect 6642 9702 6660 9720
rect 6642 9720 6660 9738
rect 6642 9738 6660 9756
rect 6642 9756 6660 9774
rect 6642 9774 6660 9792
rect 6642 9792 6660 9810
rect 6642 9810 6660 9828
rect 6642 9828 6660 9846
rect 6642 9846 6660 9864
rect 6642 9864 6660 9882
rect 6642 9882 6660 9900
rect 6642 9900 6660 9918
rect 6642 9918 6660 9936
rect 6642 9936 6660 9954
rect 6642 9954 6660 9972
rect 6642 9972 6660 9990
rect 6642 9990 6660 10008
rect 6642 10008 6660 10026
rect 6642 10026 6660 10044
rect 6660 1584 6678 1602
rect 6660 1602 6678 1620
rect 6660 1620 6678 1638
rect 6660 1638 6678 1656
rect 6660 1656 6678 1674
rect 6660 1674 6678 1692
rect 6660 1692 6678 1710
rect 6660 1710 6678 1728
rect 6660 1728 6678 1746
rect 6660 1746 6678 1764
rect 6660 1764 6678 1782
rect 6660 1782 6678 1800
rect 6660 1800 6678 1818
rect 6660 1818 6678 1836
rect 6660 1836 6678 1854
rect 6660 1854 6678 1872
rect 6660 1872 6678 1890
rect 6660 1890 6678 1908
rect 6660 1908 6678 1926
rect 6660 1926 6678 1944
rect 6660 1944 6678 1962
rect 6660 1962 6678 1980
rect 6660 1980 6678 1998
rect 6660 1998 6678 2016
rect 6660 2016 6678 2034
rect 6660 2034 6678 2052
rect 6660 2052 6678 2070
rect 6660 2070 6678 2088
rect 6660 2088 6678 2106
rect 6660 2106 6678 2124
rect 6660 2124 6678 2142
rect 6660 2142 6678 2160
rect 6660 2160 6678 2178
rect 6660 2178 6678 2196
rect 6660 2196 6678 2214
rect 6660 2214 6678 2232
rect 6660 2232 6678 2250
rect 6660 2250 6678 2268
rect 6660 2268 6678 2286
rect 6660 2286 6678 2304
rect 6660 2304 6678 2322
rect 6660 2322 6678 2340
rect 6660 2340 6678 2358
rect 6660 2358 6678 2376
rect 6660 2376 6678 2394
rect 6660 2394 6678 2412
rect 6660 2412 6678 2430
rect 6660 2430 6678 2448
rect 6660 2448 6678 2466
rect 6660 2466 6678 2484
rect 6660 2484 6678 2502
rect 6660 2502 6678 2520
rect 6660 2520 6678 2538
rect 6660 2538 6678 2556
rect 6660 2556 6678 2574
rect 6660 2574 6678 2592
rect 6660 2592 6678 2610
rect 6660 2610 6678 2628
rect 6660 2628 6678 2646
rect 6660 2646 6678 2664
rect 6660 2664 6678 2682
rect 6660 2682 6678 2700
rect 6660 2700 6678 2718
rect 6660 2718 6678 2736
rect 6660 2736 6678 2754
rect 6660 2754 6678 2772
rect 6660 2772 6678 2790
rect 6660 2790 6678 2808
rect 6660 2808 6678 2826
rect 6660 2826 6678 2844
rect 6660 2844 6678 2862
rect 6660 2862 6678 2880
rect 6660 2880 6678 2898
rect 6660 2898 6678 2916
rect 6660 2916 6678 2934
rect 6660 2934 6678 2952
rect 6660 2952 6678 2970
rect 6660 2970 6678 2988
rect 6660 3150 6678 3168
rect 6660 3168 6678 3186
rect 6660 3186 6678 3204
rect 6660 3204 6678 3222
rect 6660 3222 6678 3240
rect 6660 3240 6678 3258
rect 6660 3258 6678 3276
rect 6660 3276 6678 3294
rect 6660 3294 6678 3312
rect 6660 3312 6678 3330
rect 6660 3330 6678 3348
rect 6660 3348 6678 3366
rect 6660 3366 6678 3384
rect 6660 3384 6678 3402
rect 6660 3402 6678 3420
rect 6660 3618 6678 3636
rect 6660 3636 6678 3654
rect 6660 3654 6678 3672
rect 6660 3672 6678 3690
rect 6660 3690 6678 3708
rect 6660 3708 6678 3726
rect 6660 3726 6678 3744
rect 6660 3744 6678 3762
rect 6660 3762 6678 3780
rect 6660 3780 6678 3798
rect 6660 3798 6678 3816
rect 6660 3816 6678 3834
rect 6660 3834 6678 3852
rect 6660 3852 6678 3870
rect 6660 3870 6678 3888
rect 6660 3888 6678 3906
rect 6660 3906 6678 3924
rect 6660 3924 6678 3942
rect 6660 3942 6678 3960
rect 6660 3960 6678 3978
rect 6660 3978 6678 3996
rect 6660 3996 6678 4014
rect 6660 4014 6678 4032
rect 6660 4032 6678 4050
rect 6660 4050 6678 4068
rect 6660 4068 6678 4086
rect 6660 4086 6678 4104
rect 6660 4104 6678 4122
rect 6660 4122 6678 4140
rect 6660 4140 6678 4158
rect 6660 4158 6678 4176
rect 6660 4176 6678 4194
rect 6660 4194 6678 4212
rect 6660 4212 6678 4230
rect 6660 4230 6678 4248
rect 6660 4248 6678 4266
rect 6660 4266 6678 4284
rect 6660 4284 6678 4302
rect 6660 4302 6678 4320
rect 6660 4320 6678 4338
rect 6660 4338 6678 4356
rect 6660 4356 6678 4374
rect 6660 4374 6678 4392
rect 6660 4392 6678 4410
rect 6660 4410 6678 4428
rect 6660 4428 6678 4446
rect 6660 4446 6678 4464
rect 6660 4464 6678 4482
rect 6660 4482 6678 4500
rect 6660 4500 6678 4518
rect 6660 4518 6678 4536
rect 6660 4536 6678 4554
rect 6660 4554 6678 4572
rect 6660 4572 6678 4590
rect 6660 4590 6678 4608
rect 6660 4608 6678 4626
rect 6660 4626 6678 4644
rect 6660 4644 6678 4662
rect 6660 4662 6678 4680
rect 6660 4680 6678 4698
rect 6660 4698 6678 4716
rect 6660 4716 6678 4734
rect 6660 4734 6678 4752
rect 6660 4752 6678 4770
rect 6660 4770 6678 4788
rect 6660 4788 6678 4806
rect 6660 4806 6678 4824
rect 6660 4824 6678 4842
rect 6660 4842 6678 4860
rect 6660 4860 6678 4878
rect 6660 4878 6678 4896
rect 6660 4896 6678 4914
rect 6660 4914 6678 4932
rect 6660 4932 6678 4950
rect 6660 4950 6678 4968
rect 6660 4968 6678 4986
rect 6660 4986 6678 5004
rect 6660 5004 6678 5022
rect 6660 5022 6678 5040
rect 6660 5040 6678 5058
rect 6660 5058 6678 5076
rect 6660 5076 6678 5094
rect 6660 5094 6678 5112
rect 6660 5112 6678 5130
rect 6660 5130 6678 5148
rect 6660 5148 6678 5166
rect 6660 5166 6678 5184
rect 6660 5184 6678 5202
rect 6660 5202 6678 5220
rect 6660 5220 6678 5238
rect 6660 5238 6678 5256
rect 6660 5256 6678 5274
rect 6660 5274 6678 5292
rect 6660 5292 6678 5310
rect 6660 5310 6678 5328
rect 6660 5328 6678 5346
rect 6660 5346 6678 5364
rect 6660 5364 6678 5382
rect 6660 5382 6678 5400
rect 6660 5400 6678 5418
rect 6660 5418 6678 5436
rect 6660 5436 6678 5454
rect 6660 5454 6678 5472
rect 6660 5472 6678 5490
rect 6660 5490 6678 5508
rect 6660 5508 6678 5526
rect 6660 5526 6678 5544
rect 6660 5544 6678 5562
rect 6660 5562 6678 5580
rect 6660 5580 6678 5598
rect 6660 5598 6678 5616
rect 6660 5616 6678 5634
rect 6660 5634 6678 5652
rect 6660 5652 6678 5670
rect 6660 5670 6678 5688
rect 6660 5688 6678 5706
rect 6660 5706 6678 5724
rect 6660 5724 6678 5742
rect 6660 5742 6678 5760
rect 6660 5760 6678 5778
rect 6660 5778 6678 5796
rect 6660 5796 6678 5814
rect 6660 5814 6678 5832
rect 6660 5832 6678 5850
rect 6660 5850 6678 5868
rect 6660 5868 6678 5886
rect 6660 5886 6678 5904
rect 6660 5904 6678 5922
rect 6660 5922 6678 5940
rect 6660 5940 6678 5958
rect 6660 5958 6678 5976
rect 6660 6984 6678 7002
rect 6660 7002 6678 7020
rect 6660 7020 6678 7038
rect 6660 7038 6678 7056
rect 6660 7056 6678 7074
rect 6660 7074 6678 7092
rect 6660 7092 6678 7110
rect 6660 7110 6678 7128
rect 6660 7128 6678 7146
rect 6660 7146 6678 7164
rect 6660 7164 6678 7182
rect 6660 7182 6678 7200
rect 6660 7200 6678 7218
rect 6660 7218 6678 7236
rect 6660 7236 6678 7254
rect 6660 7254 6678 7272
rect 6660 7272 6678 7290
rect 6660 7290 6678 7308
rect 6660 7308 6678 7326
rect 6660 7326 6678 7344
rect 6660 7344 6678 7362
rect 6660 7362 6678 7380
rect 6660 7380 6678 7398
rect 6660 7398 6678 7416
rect 6660 7416 6678 7434
rect 6660 7434 6678 7452
rect 6660 7452 6678 7470
rect 6660 7470 6678 7488
rect 6660 7488 6678 7506
rect 6660 7506 6678 7524
rect 6660 7524 6678 7542
rect 6660 7542 6678 7560
rect 6660 7560 6678 7578
rect 6660 7578 6678 7596
rect 6660 7596 6678 7614
rect 6660 7614 6678 7632
rect 6660 7632 6678 7650
rect 6660 7650 6678 7668
rect 6660 7668 6678 7686
rect 6660 7686 6678 7704
rect 6660 7704 6678 7722
rect 6660 7722 6678 7740
rect 6660 7740 6678 7758
rect 6660 7758 6678 7776
rect 6660 7776 6678 7794
rect 6660 7794 6678 7812
rect 6660 7812 6678 7830
rect 6660 7830 6678 7848
rect 6660 7848 6678 7866
rect 6660 7866 6678 7884
rect 6660 7884 6678 7902
rect 6660 7902 6678 7920
rect 6660 7920 6678 7938
rect 6660 7938 6678 7956
rect 6660 7956 6678 7974
rect 6660 7974 6678 7992
rect 6660 7992 6678 8010
rect 6660 8010 6678 8028
rect 6660 8028 6678 8046
rect 6660 8046 6678 8064
rect 6660 8064 6678 8082
rect 6660 8082 6678 8100
rect 6660 8100 6678 8118
rect 6660 8118 6678 8136
rect 6660 8136 6678 8154
rect 6660 8154 6678 8172
rect 6660 8172 6678 8190
rect 6660 8190 6678 8208
rect 6660 8208 6678 8226
rect 6660 8226 6678 8244
rect 6660 8244 6678 8262
rect 6660 8262 6678 8280
rect 6660 8280 6678 8298
rect 6660 8298 6678 8316
rect 6660 8316 6678 8334
rect 6660 8334 6678 8352
rect 6660 8352 6678 8370
rect 6660 8370 6678 8388
rect 6660 8388 6678 8406
rect 6660 8406 6678 8424
rect 6660 8424 6678 8442
rect 6660 8442 6678 8460
rect 6660 8460 6678 8478
rect 6660 8478 6678 8496
rect 6660 8496 6678 8514
rect 6660 8514 6678 8532
rect 6660 8532 6678 8550
rect 6660 8550 6678 8568
rect 6660 8568 6678 8586
rect 6660 8586 6678 8604
rect 6660 8604 6678 8622
rect 6660 8622 6678 8640
rect 6660 8640 6678 8658
rect 6660 8658 6678 8676
rect 6660 8676 6678 8694
rect 6660 8694 6678 8712
rect 6660 8712 6678 8730
rect 6660 8730 6678 8748
rect 6660 8748 6678 8766
rect 6660 8766 6678 8784
rect 6660 8784 6678 8802
rect 6660 8802 6678 8820
rect 6660 8820 6678 8838
rect 6660 8838 6678 8856
rect 6660 8856 6678 8874
rect 6660 8874 6678 8892
rect 6660 8892 6678 8910
rect 6660 8910 6678 8928
rect 6660 8928 6678 8946
rect 6660 8946 6678 8964
rect 6660 8964 6678 8982
rect 6660 8982 6678 9000
rect 6660 9000 6678 9018
rect 6660 9018 6678 9036
rect 6660 9036 6678 9054
rect 6660 9054 6678 9072
rect 6660 9072 6678 9090
rect 6660 9090 6678 9108
rect 6660 9108 6678 9126
rect 6660 9126 6678 9144
rect 6660 9144 6678 9162
rect 6660 9162 6678 9180
rect 6660 9180 6678 9198
rect 6660 9198 6678 9216
rect 6660 9216 6678 9234
rect 6660 9234 6678 9252
rect 6660 9252 6678 9270
rect 6660 9270 6678 9288
rect 6660 9288 6678 9306
rect 6660 9306 6678 9324
rect 6660 9324 6678 9342
rect 6660 9342 6678 9360
rect 6660 9360 6678 9378
rect 6660 9378 6678 9396
rect 6660 9396 6678 9414
rect 6660 9414 6678 9432
rect 6660 9432 6678 9450
rect 6660 9450 6678 9468
rect 6660 9468 6678 9486
rect 6660 9486 6678 9504
rect 6660 9504 6678 9522
rect 6660 9522 6678 9540
rect 6660 9540 6678 9558
rect 6660 9558 6678 9576
rect 6660 9576 6678 9594
rect 6660 9594 6678 9612
rect 6660 9612 6678 9630
rect 6660 9630 6678 9648
rect 6660 9648 6678 9666
rect 6660 9666 6678 9684
rect 6660 9684 6678 9702
rect 6660 9702 6678 9720
rect 6660 9720 6678 9738
rect 6660 9738 6678 9756
rect 6660 9756 6678 9774
rect 6660 9774 6678 9792
rect 6660 9792 6678 9810
rect 6660 9810 6678 9828
rect 6660 9828 6678 9846
rect 6660 9846 6678 9864
rect 6660 9864 6678 9882
rect 6660 9882 6678 9900
rect 6660 9900 6678 9918
rect 6660 9918 6678 9936
rect 6660 9936 6678 9954
rect 6660 9954 6678 9972
rect 6660 9972 6678 9990
rect 6660 9990 6678 10008
rect 6660 10008 6678 10026
rect 6660 10026 6678 10044
rect 6660 10044 6678 10062
rect 6678 1602 6696 1620
rect 6678 1620 6696 1638
rect 6678 1638 6696 1656
rect 6678 1656 6696 1674
rect 6678 1674 6696 1692
rect 6678 1692 6696 1710
rect 6678 1710 6696 1728
rect 6678 1728 6696 1746
rect 6678 1746 6696 1764
rect 6678 1764 6696 1782
rect 6678 1782 6696 1800
rect 6678 1800 6696 1818
rect 6678 1818 6696 1836
rect 6678 1836 6696 1854
rect 6678 1854 6696 1872
rect 6678 1872 6696 1890
rect 6678 1890 6696 1908
rect 6678 1908 6696 1926
rect 6678 1926 6696 1944
rect 6678 1944 6696 1962
rect 6678 1962 6696 1980
rect 6678 1980 6696 1998
rect 6678 1998 6696 2016
rect 6678 2016 6696 2034
rect 6678 2034 6696 2052
rect 6678 2052 6696 2070
rect 6678 2070 6696 2088
rect 6678 2088 6696 2106
rect 6678 2106 6696 2124
rect 6678 2124 6696 2142
rect 6678 2142 6696 2160
rect 6678 2160 6696 2178
rect 6678 2178 6696 2196
rect 6678 2196 6696 2214
rect 6678 2214 6696 2232
rect 6678 2232 6696 2250
rect 6678 2250 6696 2268
rect 6678 2268 6696 2286
rect 6678 2286 6696 2304
rect 6678 2304 6696 2322
rect 6678 2322 6696 2340
rect 6678 2340 6696 2358
rect 6678 2358 6696 2376
rect 6678 2376 6696 2394
rect 6678 2394 6696 2412
rect 6678 2412 6696 2430
rect 6678 2430 6696 2448
rect 6678 2448 6696 2466
rect 6678 2466 6696 2484
rect 6678 2484 6696 2502
rect 6678 2502 6696 2520
rect 6678 2520 6696 2538
rect 6678 2538 6696 2556
rect 6678 2556 6696 2574
rect 6678 2574 6696 2592
rect 6678 2592 6696 2610
rect 6678 2610 6696 2628
rect 6678 2628 6696 2646
rect 6678 2646 6696 2664
rect 6678 2664 6696 2682
rect 6678 2682 6696 2700
rect 6678 2700 6696 2718
rect 6678 2718 6696 2736
rect 6678 2736 6696 2754
rect 6678 2754 6696 2772
rect 6678 2772 6696 2790
rect 6678 2790 6696 2808
rect 6678 2808 6696 2826
rect 6678 2826 6696 2844
rect 6678 2844 6696 2862
rect 6678 2862 6696 2880
rect 6678 2880 6696 2898
rect 6678 2898 6696 2916
rect 6678 2916 6696 2934
rect 6678 2934 6696 2952
rect 6678 2952 6696 2970
rect 6678 2970 6696 2988
rect 6678 3150 6696 3168
rect 6678 3168 6696 3186
rect 6678 3186 6696 3204
rect 6678 3204 6696 3222
rect 6678 3222 6696 3240
rect 6678 3240 6696 3258
rect 6678 3258 6696 3276
rect 6678 3276 6696 3294
rect 6678 3294 6696 3312
rect 6678 3312 6696 3330
rect 6678 3330 6696 3348
rect 6678 3348 6696 3366
rect 6678 3366 6696 3384
rect 6678 3384 6696 3402
rect 6678 3402 6696 3420
rect 6678 3420 6696 3438
rect 6678 3438 6696 3456
rect 6678 3636 6696 3654
rect 6678 3654 6696 3672
rect 6678 3672 6696 3690
rect 6678 3690 6696 3708
rect 6678 3708 6696 3726
rect 6678 3726 6696 3744
rect 6678 3744 6696 3762
rect 6678 3762 6696 3780
rect 6678 3780 6696 3798
rect 6678 3798 6696 3816
rect 6678 3816 6696 3834
rect 6678 3834 6696 3852
rect 6678 3852 6696 3870
rect 6678 3870 6696 3888
rect 6678 3888 6696 3906
rect 6678 3906 6696 3924
rect 6678 3924 6696 3942
rect 6678 3942 6696 3960
rect 6678 3960 6696 3978
rect 6678 3978 6696 3996
rect 6678 3996 6696 4014
rect 6678 4014 6696 4032
rect 6678 4032 6696 4050
rect 6678 4050 6696 4068
rect 6678 4068 6696 4086
rect 6678 4086 6696 4104
rect 6678 4104 6696 4122
rect 6678 4122 6696 4140
rect 6678 4140 6696 4158
rect 6678 4158 6696 4176
rect 6678 4176 6696 4194
rect 6678 4194 6696 4212
rect 6678 4212 6696 4230
rect 6678 4230 6696 4248
rect 6678 4248 6696 4266
rect 6678 4266 6696 4284
rect 6678 4284 6696 4302
rect 6678 4302 6696 4320
rect 6678 4320 6696 4338
rect 6678 4338 6696 4356
rect 6678 4356 6696 4374
rect 6678 4374 6696 4392
rect 6678 4392 6696 4410
rect 6678 4410 6696 4428
rect 6678 4428 6696 4446
rect 6678 4446 6696 4464
rect 6678 4464 6696 4482
rect 6678 4482 6696 4500
rect 6678 4500 6696 4518
rect 6678 4518 6696 4536
rect 6678 4536 6696 4554
rect 6678 4554 6696 4572
rect 6678 4572 6696 4590
rect 6678 4590 6696 4608
rect 6678 4608 6696 4626
rect 6678 4626 6696 4644
rect 6678 4644 6696 4662
rect 6678 4662 6696 4680
rect 6678 4680 6696 4698
rect 6678 4698 6696 4716
rect 6678 4716 6696 4734
rect 6678 4734 6696 4752
rect 6678 4752 6696 4770
rect 6678 4770 6696 4788
rect 6678 4788 6696 4806
rect 6678 4806 6696 4824
rect 6678 4824 6696 4842
rect 6678 4842 6696 4860
rect 6678 4860 6696 4878
rect 6678 4878 6696 4896
rect 6678 4896 6696 4914
rect 6678 4914 6696 4932
rect 6678 4932 6696 4950
rect 6678 4950 6696 4968
rect 6678 4968 6696 4986
rect 6678 4986 6696 5004
rect 6678 5004 6696 5022
rect 6678 5022 6696 5040
rect 6678 5040 6696 5058
rect 6678 5058 6696 5076
rect 6678 5076 6696 5094
rect 6678 5094 6696 5112
rect 6678 5112 6696 5130
rect 6678 5130 6696 5148
rect 6678 5148 6696 5166
rect 6678 5166 6696 5184
rect 6678 5184 6696 5202
rect 6678 5202 6696 5220
rect 6678 5220 6696 5238
rect 6678 5238 6696 5256
rect 6678 5256 6696 5274
rect 6678 5274 6696 5292
rect 6678 5292 6696 5310
rect 6678 5310 6696 5328
rect 6678 5328 6696 5346
rect 6678 5346 6696 5364
rect 6678 5364 6696 5382
rect 6678 5382 6696 5400
rect 6678 5400 6696 5418
rect 6678 5418 6696 5436
rect 6678 5436 6696 5454
rect 6678 5454 6696 5472
rect 6678 5472 6696 5490
rect 6678 5490 6696 5508
rect 6678 5508 6696 5526
rect 6678 5526 6696 5544
rect 6678 5544 6696 5562
rect 6678 5562 6696 5580
rect 6678 5580 6696 5598
rect 6678 5598 6696 5616
rect 6678 5616 6696 5634
rect 6678 5634 6696 5652
rect 6678 5652 6696 5670
rect 6678 5670 6696 5688
rect 6678 5688 6696 5706
rect 6678 5706 6696 5724
rect 6678 5724 6696 5742
rect 6678 5742 6696 5760
rect 6678 5760 6696 5778
rect 6678 5778 6696 5796
rect 6678 5796 6696 5814
rect 6678 5814 6696 5832
rect 6678 5832 6696 5850
rect 6678 5850 6696 5868
rect 6678 5868 6696 5886
rect 6678 5886 6696 5904
rect 6678 5904 6696 5922
rect 6678 5922 6696 5940
rect 6678 5940 6696 5958
rect 6678 5958 6696 5976
rect 6678 5976 6696 5994
rect 6678 7020 6696 7038
rect 6678 7038 6696 7056
rect 6678 7056 6696 7074
rect 6678 7074 6696 7092
rect 6678 7092 6696 7110
rect 6678 7110 6696 7128
rect 6678 7128 6696 7146
rect 6678 7146 6696 7164
rect 6678 7164 6696 7182
rect 6678 7182 6696 7200
rect 6678 7200 6696 7218
rect 6678 7218 6696 7236
rect 6678 7236 6696 7254
rect 6678 7254 6696 7272
rect 6678 7272 6696 7290
rect 6678 7290 6696 7308
rect 6678 7308 6696 7326
rect 6678 7326 6696 7344
rect 6678 7344 6696 7362
rect 6678 7362 6696 7380
rect 6678 7380 6696 7398
rect 6678 7398 6696 7416
rect 6678 7416 6696 7434
rect 6678 7434 6696 7452
rect 6678 7452 6696 7470
rect 6678 7470 6696 7488
rect 6678 7488 6696 7506
rect 6678 7506 6696 7524
rect 6678 7524 6696 7542
rect 6678 7542 6696 7560
rect 6678 7560 6696 7578
rect 6678 7578 6696 7596
rect 6678 7596 6696 7614
rect 6678 7614 6696 7632
rect 6678 7632 6696 7650
rect 6678 7650 6696 7668
rect 6678 7668 6696 7686
rect 6678 7686 6696 7704
rect 6678 7704 6696 7722
rect 6678 7722 6696 7740
rect 6678 7740 6696 7758
rect 6678 7758 6696 7776
rect 6678 7776 6696 7794
rect 6678 7794 6696 7812
rect 6678 7812 6696 7830
rect 6678 7830 6696 7848
rect 6678 7848 6696 7866
rect 6678 7866 6696 7884
rect 6678 7884 6696 7902
rect 6678 7902 6696 7920
rect 6678 7920 6696 7938
rect 6678 7938 6696 7956
rect 6678 7956 6696 7974
rect 6678 7974 6696 7992
rect 6678 7992 6696 8010
rect 6678 8010 6696 8028
rect 6678 8028 6696 8046
rect 6678 8046 6696 8064
rect 6678 8064 6696 8082
rect 6678 8082 6696 8100
rect 6678 8100 6696 8118
rect 6678 8118 6696 8136
rect 6678 8136 6696 8154
rect 6678 8154 6696 8172
rect 6678 8172 6696 8190
rect 6678 8190 6696 8208
rect 6678 8208 6696 8226
rect 6678 8226 6696 8244
rect 6678 8244 6696 8262
rect 6678 8262 6696 8280
rect 6678 8280 6696 8298
rect 6678 8298 6696 8316
rect 6678 8316 6696 8334
rect 6678 8334 6696 8352
rect 6678 8352 6696 8370
rect 6678 8370 6696 8388
rect 6678 8388 6696 8406
rect 6678 8406 6696 8424
rect 6678 8424 6696 8442
rect 6678 8442 6696 8460
rect 6678 8460 6696 8478
rect 6678 8478 6696 8496
rect 6678 8496 6696 8514
rect 6678 8514 6696 8532
rect 6678 8532 6696 8550
rect 6678 8550 6696 8568
rect 6678 8568 6696 8586
rect 6678 8586 6696 8604
rect 6678 8604 6696 8622
rect 6678 8622 6696 8640
rect 6678 8640 6696 8658
rect 6678 8658 6696 8676
rect 6678 8676 6696 8694
rect 6678 8694 6696 8712
rect 6678 8712 6696 8730
rect 6678 8730 6696 8748
rect 6678 8748 6696 8766
rect 6678 8766 6696 8784
rect 6678 8784 6696 8802
rect 6678 8802 6696 8820
rect 6678 8820 6696 8838
rect 6678 8838 6696 8856
rect 6678 8856 6696 8874
rect 6678 8874 6696 8892
rect 6678 8892 6696 8910
rect 6678 8910 6696 8928
rect 6678 8928 6696 8946
rect 6678 8946 6696 8964
rect 6678 8964 6696 8982
rect 6678 8982 6696 9000
rect 6678 9000 6696 9018
rect 6678 9018 6696 9036
rect 6678 9036 6696 9054
rect 6678 9054 6696 9072
rect 6678 9072 6696 9090
rect 6678 9090 6696 9108
rect 6678 9108 6696 9126
rect 6678 9126 6696 9144
rect 6678 9144 6696 9162
rect 6678 9162 6696 9180
rect 6678 9180 6696 9198
rect 6678 9198 6696 9216
rect 6678 9216 6696 9234
rect 6678 9234 6696 9252
rect 6678 9252 6696 9270
rect 6678 9270 6696 9288
rect 6678 9288 6696 9306
rect 6678 9306 6696 9324
rect 6678 9324 6696 9342
rect 6678 9342 6696 9360
rect 6678 9360 6696 9378
rect 6678 9378 6696 9396
rect 6678 9396 6696 9414
rect 6678 9414 6696 9432
rect 6678 9432 6696 9450
rect 6678 9450 6696 9468
rect 6678 9468 6696 9486
rect 6678 9486 6696 9504
rect 6678 9504 6696 9522
rect 6678 9522 6696 9540
rect 6678 9540 6696 9558
rect 6678 9558 6696 9576
rect 6678 9576 6696 9594
rect 6678 9594 6696 9612
rect 6678 9612 6696 9630
rect 6678 9630 6696 9648
rect 6678 9648 6696 9666
rect 6678 9666 6696 9684
rect 6678 9684 6696 9702
rect 6678 9702 6696 9720
rect 6678 9720 6696 9738
rect 6678 9738 6696 9756
rect 6678 9756 6696 9774
rect 6678 9774 6696 9792
rect 6678 9792 6696 9810
rect 6678 9810 6696 9828
rect 6678 9828 6696 9846
rect 6678 9846 6696 9864
rect 6678 9864 6696 9882
rect 6678 9882 6696 9900
rect 6678 9900 6696 9918
rect 6678 9918 6696 9936
rect 6678 9936 6696 9954
rect 6678 9954 6696 9972
rect 6678 9972 6696 9990
rect 6678 9990 6696 10008
rect 6678 10008 6696 10026
rect 6678 10026 6696 10044
rect 6678 10044 6696 10062
rect 6678 10062 6696 10080
rect 6696 1602 6714 1620
rect 6696 1620 6714 1638
rect 6696 1638 6714 1656
rect 6696 1656 6714 1674
rect 6696 1674 6714 1692
rect 6696 1692 6714 1710
rect 6696 1710 6714 1728
rect 6696 1728 6714 1746
rect 6696 1746 6714 1764
rect 6696 1764 6714 1782
rect 6696 1782 6714 1800
rect 6696 1800 6714 1818
rect 6696 1818 6714 1836
rect 6696 1836 6714 1854
rect 6696 1854 6714 1872
rect 6696 1872 6714 1890
rect 6696 1890 6714 1908
rect 6696 1908 6714 1926
rect 6696 1926 6714 1944
rect 6696 1944 6714 1962
rect 6696 1962 6714 1980
rect 6696 1980 6714 1998
rect 6696 1998 6714 2016
rect 6696 2016 6714 2034
rect 6696 2034 6714 2052
rect 6696 2052 6714 2070
rect 6696 2070 6714 2088
rect 6696 2088 6714 2106
rect 6696 2106 6714 2124
rect 6696 2124 6714 2142
rect 6696 2142 6714 2160
rect 6696 2160 6714 2178
rect 6696 2178 6714 2196
rect 6696 2196 6714 2214
rect 6696 2214 6714 2232
rect 6696 2232 6714 2250
rect 6696 2250 6714 2268
rect 6696 2268 6714 2286
rect 6696 2286 6714 2304
rect 6696 2304 6714 2322
rect 6696 2322 6714 2340
rect 6696 2340 6714 2358
rect 6696 2358 6714 2376
rect 6696 2376 6714 2394
rect 6696 2394 6714 2412
rect 6696 2412 6714 2430
rect 6696 2430 6714 2448
rect 6696 2448 6714 2466
rect 6696 2466 6714 2484
rect 6696 2484 6714 2502
rect 6696 2502 6714 2520
rect 6696 2520 6714 2538
rect 6696 2538 6714 2556
rect 6696 2556 6714 2574
rect 6696 2574 6714 2592
rect 6696 2592 6714 2610
rect 6696 2610 6714 2628
rect 6696 2628 6714 2646
rect 6696 2646 6714 2664
rect 6696 2664 6714 2682
rect 6696 2682 6714 2700
rect 6696 2700 6714 2718
rect 6696 2718 6714 2736
rect 6696 2736 6714 2754
rect 6696 2754 6714 2772
rect 6696 2772 6714 2790
rect 6696 2790 6714 2808
rect 6696 2808 6714 2826
rect 6696 2826 6714 2844
rect 6696 2844 6714 2862
rect 6696 2862 6714 2880
rect 6696 2880 6714 2898
rect 6696 2898 6714 2916
rect 6696 2916 6714 2934
rect 6696 2934 6714 2952
rect 6696 2952 6714 2970
rect 6696 2970 6714 2988
rect 6696 2988 6714 3006
rect 6696 3168 6714 3186
rect 6696 3186 6714 3204
rect 6696 3204 6714 3222
rect 6696 3222 6714 3240
rect 6696 3240 6714 3258
rect 6696 3258 6714 3276
rect 6696 3276 6714 3294
rect 6696 3294 6714 3312
rect 6696 3312 6714 3330
rect 6696 3330 6714 3348
rect 6696 3348 6714 3366
rect 6696 3366 6714 3384
rect 6696 3384 6714 3402
rect 6696 3402 6714 3420
rect 6696 3420 6714 3438
rect 6696 3438 6714 3456
rect 6696 3456 6714 3474
rect 6696 3654 6714 3672
rect 6696 3672 6714 3690
rect 6696 3690 6714 3708
rect 6696 3708 6714 3726
rect 6696 3726 6714 3744
rect 6696 3744 6714 3762
rect 6696 3762 6714 3780
rect 6696 3780 6714 3798
rect 6696 3798 6714 3816
rect 6696 3816 6714 3834
rect 6696 3834 6714 3852
rect 6696 3852 6714 3870
rect 6696 3870 6714 3888
rect 6696 3888 6714 3906
rect 6696 3906 6714 3924
rect 6696 3924 6714 3942
rect 6696 3942 6714 3960
rect 6696 3960 6714 3978
rect 6696 3978 6714 3996
rect 6696 3996 6714 4014
rect 6696 4014 6714 4032
rect 6696 4032 6714 4050
rect 6696 4050 6714 4068
rect 6696 4068 6714 4086
rect 6696 4086 6714 4104
rect 6696 4104 6714 4122
rect 6696 4122 6714 4140
rect 6696 4140 6714 4158
rect 6696 4158 6714 4176
rect 6696 4176 6714 4194
rect 6696 4194 6714 4212
rect 6696 4212 6714 4230
rect 6696 4230 6714 4248
rect 6696 4248 6714 4266
rect 6696 4266 6714 4284
rect 6696 4284 6714 4302
rect 6696 4302 6714 4320
rect 6696 4320 6714 4338
rect 6696 4338 6714 4356
rect 6696 4356 6714 4374
rect 6696 4374 6714 4392
rect 6696 4392 6714 4410
rect 6696 4410 6714 4428
rect 6696 4428 6714 4446
rect 6696 4446 6714 4464
rect 6696 4464 6714 4482
rect 6696 4482 6714 4500
rect 6696 4500 6714 4518
rect 6696 4518 6714 4536
rect 6696 4536 6714 4554
rect 6696 4554 6714 4572
rect 6696 4572 6714 4590
rect 6696 4590 6714 4608
rect 6696 4608 6714 4626
rect 6696 4626 6714 4644
rect 6696 4644 6714 4662
rect 6696 4662 6714 4680
rect 6696 4680 6714 4698
rect 6696 4698 6714 4716
rect 6696 4716 6714 4734
rect 6696 4734 6714 4752
rect 6696 4752 6714 4770
rect 6696 4770 6714 4788
rect 6696 4788 6714 4806
rect 6696 4806 6714 4824
rect 6696 4824 6714 4842
rect 6696 4842 6714 4860
rect 6696 4860 6714 4878
rect 6696 4878 6714 4896
rect 6696 4896 6714 4914
rect 6696 4914 6714 4932
rect 6696 4932 6714 4950
rect 6696 4950 6714 4968
rect 6696 4968 6714 4986
rect 6696 4986 6714 5004
rect 6696 5004 6714 5022
rect 6696 5022 6714 5040
rect 6696 5040 6714 5058
rect 6696 5058 6714 5076
rect 6696 5076 6714 5094
rect 6696 5094 6714 5112
rect 6696 5112 6714 5130
rect 6696 5130 6714 5148
rect 6696 5148 6714 5166
rect 6696 5166 6714 5184
rect 6696 5184 6714 5202
rect 6696 5202 6714 5220
rect 6696 5220 6714 5238
rect 6696 5238 6714 5256
rect 6696 5256 6714 5274
rect 6696 5274 6714 5292
rect 6696 5292 6714 5310
rect 6696 5310 6714 5328
rect 6696 5328 6714 5346
rect 6696 5346 6714 5364
rect 6696 5364 6714 5382
rect 6696 5382 6714 5400
rect 6696 5400 6714 5418
rect 6696 5418 6714 5436
rect 6696 5436 6714 5454
rect 6696 5454 6714 5472
rect 6696 5472 6714 5490
rect 6696 5490 6714 5508
rect 6696 5508 6714 5526
rect 6696 5526 6714 5544
rect 6696 5544 6714 5562
rect 6696 5562 6714 5580
rect 6696 5580 6714 5598
rect 6696 5598 6714 5616
rect 6696 5616 6714 5634
rect 6696 5634 6714 5652
rect 6696 5652 6714 5670
rect 6696 5670 6714 5688
rect 6696 5688 6714 5706
rect 6696 5706 6714 5724
rect 6696 5724 6714 5742
rect 6696 5742 6714 5760
rect 6696 5760 6714 5778
rect 6696 5778 6714 5796
rect 6696 5796 6714 5814
rect 6696 5814 6714 5832
rect 6696 5832 6714 5850
rect 6696 5850 6714 5868
rect 6696 5868 6714 5886
rect 6696 5886 6714 5904
rect 6696 5904 6714 5922
rect 6696 5922 6714 5940
rect 6696 5940 6714 5958
rect 6696 5958 6714 5976
rect 6696 5976 6714 5994
rect 6696 5994 6714 6012
rect 6696 7074 6714 7092
rect 6696 7092 6714 7110
rect 6696 7110 6714 7128
rect 6696 7128 6714 7146
rect 6696 7146 6714 7164
rect 6696 7164 6714 7182
rect 6696 7182 6714 7200
rect 6696 7200 6714 7218
rect 6696 7218 6714 7236
rect 6696 7236 6714 7254
rect 6696 7254 6714 7272
rect 6696 7272 6714 7290
rect 6696 7290 6714 7308
rect 6696 7308 6714 7326
rect 6696 7326 6714 7344
rect 6696 7344 6714 7362
rect 6696 7362 6714 7380
rect 6696 7380 6714 7398
rect 6696 7398 6714 7416
rect 6696 7416 6714 7434
rect 6696 7434 6714 7452
rect 6696 7452 6714 7470
rect 6696 7470 6714 7488
rect 6696 7488 6714 7506
rect 6696 7506 6714 7524
rect 6696 7524 6714 7542
rect 6696 7542 6714 7560
rect 6696 7560 6714 7578
rect 6696 7578 6714 7596
rect 6696 7596 6714 7614
rect 6696 7614 6714 7632
rect 6696 7632 6714 7650
rect 6696 7650 6714 7668
rect 6696 7668 6714 7686
rect 6696 7686 6714 7704
rect 6696 7704 6714 7722
rect 6696 7722 6714 7740
rect 6696 7740 6714 7758
rect 6696 7758 6714 7776
rect 6696 7776 6714 7794
rect 6696 7794 6714 7812
rect 6696 7812 6714 7830
rect 6696 7830 6714 7848
rect 6696 7848 6714 7866
rect 6696 7866 6714 7884
rect 6696 7884 6714 7902
rect 6696 7902 6714 7920
rect 6696 7920 6714 7938
rect 6696 7938 6714 7956
rect 6696 7956 6714 7974
rect 6696 7974 6714 7992
rect 6696 7992 6714 8010
rect 6696 8010 6714 8028
rect 6696 8028 6714 8046
rect 6696 8046 6714 8064
rect 6696 8064 6714 8082
rect 6696 8082 6714 8100
rect 6696 8100 6714 8118
rect 6696 8118 6714 8136
rect 6696 8136 6714 8154
rect 6696 8154 6714 8172
rect 6696 8172 6714 8190
rect 6696 8190 6714 8208
rect 6696 8208 6714 8226
rect 6696 8226 6714 8244
rect 6696 8244 6714 8262
rect 6696 8262 6714 8280
rect 6696 8280 6714 8298
rect 6696 8298 6714 8316
rect 6696 8316 6714 8334
rect 6696 8334 6714 8352
rect 6696 8352 6714 8370
rect 6696 8370 6714 8388
rect 6696 8388 6714 8406
rect 6696 8406 6714 8424
rect 6696 8424 6714 8442
rect 6696 8442 6714 8460
rect 6696 8460 6714 8478
rect 6696 8478 6714 8496
rect 6696 8496 6714 8514
rect 6696 8514 6714 8532
rect 6696 8532 6714 8550
rect 6696 8550 6714 8568
rect 6696 8568 6714 8586
rect 6696 8586 6714 8604
rect 6696 8604 6714 8622
rect 6696 8622 6714 8640
rect 6696 8640 6714 8658
rect 6696 8658 6714 8676
rect 6696 8676 6714 8694
rect 6696 8694 6714 8712
rect 6696 8712 6714 8730
rect 6696 8730 6714 8748
rect 6696 8748 6714 8766
rect 6696 8766 6714 8784
rect 6696 8784 6714 8802
rect 6696 8802 6714 8820
rect 6696 8820 6714 8838
rect 6696 8838 6714 8856
rect 6696 8856 6714 8874
rect 6696 8874 6714 8892
rect 6696 8892 6714 8910
rect 6696 8910 6714 8928
rect 6696 8928 6714 8946
rect 6696 8946 6714 8964
rect 6696 8964 6714 8982
rect 6696 8982 6714 9000
rect 6696 9000 6714 9018
rect 6696 9018 6714 9036
rect 6696 9036 6714 9054
rect 6696 9054 6714 9072
rect 6696 9072 6714 9090
rect 6696 9090 6714 9108
rect 6696 9108 6714 9126
rect 6696 9126 6714 9144
rect 6696 9144 6714 9162
rect 6696 9162 6714 9180
rect 6696 9180 6714 9198
rect 6696 9198 6714 9216
rect 6696 9216 6714 9234
rect 6696 9234 6714 9252
rect 6696 9252 6714 9270
rect 6696 9270 6714 9288
rect 6696 9288 6714 9306
rect 6696 9306 6714 9324
rect 6696 9324 6714 9342
rect 6696 9342 6714 9360
rect 6696 9360 6714 9378
rect 6696 9378 6714 9396
rect 6696 9396 6714 9414
rect 6696 9414 6714 9432
rect 6696 9432 6714 9450
rect 6696 9450 6714 9468
rect 6696 9468 6714 9486
rect 6696 9486 6714 9504
rect 6696 9504 6714 9522
rect 6696 9522 6714 9540
rect 6696 9540 6714 9558
rect 6696 9558 6714 9576
rect 6696 9576 6714 9594
rect 6696 9594 6714 9612
rect 6696 9612 6714 9630
rect 6696 9630 6714 9648
rect 6696 9648 6714 9666
rect 6696 9666 6714 9684
rect 6696 9684 6714 9702
rect 6696 9702 6714 9720
rect 6696 9720 6714 9738
rect 6696 9738 6714 9756
rect 6696 9756 6714 9774
rect 6696 9774 6714 9792
rect 6696 9792 6714 9810
rect 6696 9810 6714 9828
rect 6696 9828 6714 9846
rect 6696 9846 6714 9864
rect 6696 9864 6714 9882
rect 6696 9882 6714 9900
rect 6696 9900 6714 9918
rect 6696 9918 6714 9936
rect 6696 9936 6714 9954
rect 6696 9954 6714 9972
rect 6696 9972 6714 9990
rect 6696 9990 6714 10008
rect 6696 10008 6714 10026
rect 6696 10026 6714 10044
rect 6696 10044 6714 10062
rect 6696 10062 6714 10080
rect 6696 10080 6714 10098
rect 6696 10098 6714 10116
rect 6714 1620 6732 1638
rect 6714 1638 6732 1656
rect 6714 1656 6732 1674
rect 6714 1674 6732 1692
rect 6714 1692 6732 1710
rect 6714 1710 6732 1728
rect 6714 1728 6732 1746
rect 6714 1746 6732 1764
rect 6714 1764 6732 1782
rect 6714 1782 6732 1800
rect 6714 1800 6732 1818
rect 6714 1818 6732 1836
rect 6714 1836 6732 1854
rect 6714 1854 6732 1872
rect 6714 1872 6732 1890
rect 6714 1890 6732 1908
rect 6714 1908 6732 1926
rect 6714 1926 6732 1944
rect 6714 1944 6732 1962
rect 6714 1962 6732 1980
rect 6714 1980 6732 1998
rect 6714 1998 6732 2016
rect 6714 2016 6732 2034
rect 6714 2034 6732 2052
rect 6714 2052 6732 2070
rect 6714 2070 6732 2088
rect 6714 2088 6732 2106
rect 6714 2106 6732 2124
rect 6714 2124 6732 2142
rect 6714 2142 6732 2160
rect 6714 2160 6732 2178
rect 6714 2178 6732 2196
rect 6714 2196 6732 2214
rect 6714 2214 6732 2232
rect 6714 2232 6732 2250
rect 6714 2250 6732 2268
rect 6714 2268 6732 2286
rect 6714 2286 6732 2304
rect 6714 2304 6732 2322
rect 6714 2322 6732 2340
rect 6714 2340 6732 2358
rect 6714 2358 6732 2376
rect 6714 2376 6732 2394
rect 6714 2394 6732 2412
rect 6714 2412 6732 2430
rect 6714 2430 6732 2448
rect 6714 2448 6732 2466
rect 6714 2466 6732 2484
rect 6714 2484 6732 2502
rect 6714 2502 6732 2520
rect 6714 2520 6732 2538
rect 6714 2538 6732 2556
rect 6714 2556 6732 2574
rect 6714 2574 6732 2592
rect 6714 2592 6732 2610
rect 6714 2610 6732 2628
rect 6714 2628 6732 2646
rect 6714 2646 6732 2664
rect 6714 2664 6732 2682
rect 6714 2682 6732 2700
rect 6714 2700 6732 2718
rect 6714 2718 6732 2736
rect 6714 2736 6732 2754
rect 6714 2754 6732 2772
rect 6714 2772 6732 2790
rect 6714 2790 6732 2808
rect 6714 2808 6732 2826
rect 6714 2826 6732 2844
rect 6714 2844 6732 2862
rect 6714 2862 6732 2880
rect 6714 2880 6732 2898
rect 6714 2898 6732 2916
rect 6714 2916 6732 2934
rect 6714 2934 6732 2952
rect 6714 2952 6732 2970
rect 6714 2970 6732 2988
rect 6714 2988 6732 3006
rect 6714 3168 6732 3186
rect 6714 3186 6732 3204
rect 6714 3204 6732 3222
rect 6714 3222 6732 3240
rect 6714 3240 6732 3258
rect 6714 3258 6732 3276
rect 6714 3276 6732 3294
rect 6714 3294 6732 3312
rect 6714 3312 6732 3330
rect 6714 3330 6732 3348
rect 6714 3348 6732 3366
rect 6714 3366 6732 3384
rect 6714 3384 6732 3402
rect 6714 3402 6732 3420
rect 6714 3420 6732 3438
rect 6714 3438 6732 3456
rect 6714 3456 6732 3474
rect 6714 3474 6732 3492
rect 6714 3672 6732 3690
rect 6714 3690 6732 3708
rect 6714 3708 6732 3726
rect 6714 3726 6732 3744
rect 6714 3744 6732 3762
rect 6714 3762 6732 3780
rect 6714 3780 6732 3798
rect 6714 3798 6732 3816
rect 6714 3816 6732 3834
rect 6714 3834 6732 3852
rect 6714 3852 6732 3870
rect 6714 3870 6732 3888
rect 6714 3888 6732 3906
rect 6714 3906 6732 3924
rect 6714 3924 6732 3942
rect 6714 3942 6732 3960
rect 6714 3960 6732 3978
rect 6714 3978 6732 3996
rect 6714 3996 6732 4014
rect 6714 4014 6732 4032
rect 6714 4032 6732 4050
rect 6714 4050 6732 4068
rect 6714 4068 6732 4086
rect 6714 4086 6732 4104
rect 6714 4104 6732 4122
rect 6714 4122 6732 4140
rect 6714 4140 6732 4158
rect 6714 4158 6732 4176
rect 6714 4176 6732 4194
rect 6714 4194 6732 4212
rect 6714 4212 6732 4230
rect 6714 4230 6732 4248
rect 6714 4248 6732 4266
rect 6714 4266 6732 4284
rect 6714 4284 6732 4302
rect 6714 4302 6732 4320
rect 6714 4320 6732 4338
rect 6714 4338 6732 4356
rect 6714 4356 6732 4374
rect 6714 4374 6732 4392
rect 6714 4392 6732 4410
rect 6714 4410 6732 4428
rect 6714 4428 6732 4446
rect 6714 4446 6732 4464
rect 6714 4464 6732 4482
rect 6714 4482 6732 4500
rect 6714 4500 6732 4518
rect 6714 4518 6732 4536
rect 6714 4536 6732 4554
rect 6714 4554 6732 4572
rect 6714 4572 6732 4590
rect 6714 4590 6732 4608
rect 6714 4608 6732 4626
rect 6714 4626 6732 4644
rect 6714 4644 6732 4662
rect 6714 4662 6732 4680
rect 6714 4680 6732 4698
rect 6714 4698 6732 4716
rect 6714 4716 6732 4734
rect 6714 4734 6732 4752
rect 6714 4752 6732 4770
rect 6714 4770 6732 4788
rect 6714 4788 6732 4806
rect 6714 4806 6732 4824
rect 6714 4824 6732 4842
rect 6714 4842 6732 4860
rect 6714 4860 6732 4878
rect 6714 4878 6732 4896
rect 6714 4896 6732 4914
rect 6714 4914 6732 4932
rect 6714 4932 6732 4950
rect 6714 4950 6732 4968
rect 6714 4968 6732 4986
rect 6714 4986 6732 5004
rect 6714 5004 6732 5022
rect 6714 5022 6732 5040
rect 6714 5040 6732 5058
rect 6714 5058 6732 5076
rect 6714 5076 6732 5094
rect 6714 5094 6732 5112
rect 6714 5112 6732 5130
rect 6714 5130 6732 5148
rect 6714 5148 6732 5166
rect 6714 5166 6732 5184
rect 6714 5184 6732 5202
rect 6714 5202 6732 5220
rect 6714 5220 6732 5238
rect 6714 5238 6732 5256
rect 6714 5256 6732 5274
rect 6714 5274 6732 5292
rect 6714 5292 6732 5310
rect 6714 5310 6732 5328
rect 6714 5328 6732 5346
rect 6714 5346 6732 5364
rect 6714 5364 6732 5382
rect 6714 5382 6732 5400
rect 6714 5400 6732 5418
rect 6714 5418 6732 5436
rect 6714 5436 6732 5454
rect 6714 5454 6732 5472
rect 6714 5472 6732 5490
rect 6714 5490 6732 5508
rect 6714 5508 6732 5526
rect 6714 5526 6732 5544
rect 6714 5544 6732 5562
rect 6714 5562 6732 5580
rect 6714 5580 6732 5598
rect 6714 5598 6732 5616
rect 6714 5616 6732 5634
rect 6714 5634 6732 5652
rect 6714 5652 6732 5670
rect 6714 5670 6732 5688
rect 6714 5688 6732 5706
rect 6714 5706 6732 5724
rect 6714 5724 6732 5742
rect 6714 5742 6732 5760
rect 6714 5760 6732 5778
rect 6714 5778 6732 5796
rect 6714 5796 6732 5814
rect 6714 5814 6732 5832
rect 6714 5832 6732 5850
rect 6714 5850 6732 5868
rect 6714 5868 6732 5886
rect 6714 5886 6732 5904
rect 6714 5904 6732 5922
rect 6714 5922 6732 5940
rect 6714 5940 6732 5958
rect 6714 5958 6732 5976
rect 6714 5976 6732 5994
rect 6714 5994 6732 6012
rect 6714 6012 6732 6030
rect 6714 7110 6732 7128
rect 6714 7128 6732 7146
rect 6714 7146 6732 7164
rect 6714 7164 6732 7182
rect 6714 7182 6732 7200
rect 6714 7200 6732 7218
rect 6714 7218 6732 7236
rect 6714 7236 6732 7254
rect 6714 7254 6732 7272
rect 6714 7272 6732 7290
rect 6714 7290 6732 7308
rect 6714 7308 6732 7326
rect 6714 7326 6732 7344
rect 6714 7344 6732 7362
rect 6714 7362 6732 7380
rect 6714 7380 6732 7398
rect 6714 7398 6732 7416
rect 6714 7416 6732 7434
rect 6714 7434 6732 7452
rect 6714 7452 6732 7470
rect 6714 7470 6732 7488
rect 6714 7488 6732 7506
rect 6714 7506 6732 7524
rect 6714 7524 6732 7542
rect 6714 7542 6732 7560
rect 6714 7560 6732 7578
rect 6714 7578 6732 7596
rect 6714 7596 6732 7614
rect 6714 7614 6732 7632
rect 6714 7632 6732 7650
rect 6714 7650 6732 7668
rect 6714 7668 6732 7686
rect 6714 7686 6732 7704
rect 6714 7704 6732 7722
rect 6714 7722 6732 7740
rect 6714 7740 6732 7758
rect 6714 7758 6732 7776
rect 6714 7776 6732 7794
rect 6714 7794 6732 7812
rect 6714 7812 6732 7830
rect 6714 7830 6732 7848
rect 6714 7848 6732 7866
rect 6714 7866 6732 7884
rect 6714 7884 6732 7902
rect 6714 7902 6732 7920
rect 6714 7920 6732 7938
rect 6714 7938 6732 7956
rect 6714 7956 6732 7974
rect 6714 7974 6732 7992
rect 6714 7992 6732 8010
rect 6714 8010 6732 8028
rect 6714 8028 6732 8046
rect 6714 8046 6732 8064
rect 6714 8064 6732 8082
rect 6714 8082 6732 8100
rect 6714 8100 6732 8118
rect 6714 8118 6732 8136
rect 6714 8136 6732 8154
rect 6714 8154 6732 8172
rect 6714 8172 6732 8190
rect 6714 8190 6732 8208
rect 6714 8208 6732 8226
rect 6714 8226 6732 8244
rect 6714 8244 6732 8262
rect 6714 8262 6732 8280
rect 6714 8280 6732 8298
rect 6714 8298 6732 8316
rect 6714 8316 6732 8334
rect 6714 8334 6732 8352
rect 6714 8352 6732 8370
rect 6714 8370 6732 8388
rect 6714 8388 6732 8406
rect 6714 8406 6732 8424
rect 6714 8424 6732 8442
rect 6714 8442 6732 8460
rect 6714 8460 6732 8478
rect 6714 8478 6732 8496
rect 6714 8496 6732 8514
rect 6714 8514 6732 8532
rect 6714 8532 6732 8550
rect 6714 8550 6732 8568
rect 6714 8568 6732 8586
rect 6714 8586 6732 8604
rect 6714 8604 6732 8622
rect 6714 8622 6732 8640
rect 6714 8640 6732 8658
rect 6714 8658 6732 8676
rect 6714 8676 6732 8694
rect 6714 8694 6732 8712
rect 6714 8712 6732 8730
rect 6714 8730 6732 8748
rect 6714 8748 6732 8766
rect 6714 8766 6732 8784
rect 6714 8784 6732 8802
rect 6714 8802 6732 8820
rect 6714 8820 6732 8838
rect 6714 8838 6732 8856
rect 6714 8856 6732 8874
rect 6714 8874 6732 8892
rect 6714 8892 6732 8910
rect 6714 8910 6732 8928
rect 6714 8928 6732 8946
rect 6714 8946 6732 8964
rect 6714 8964 6732 8982
rect 6714 8982 6732 9000
rect 6714 9000 6732 9018
rect 6714 9018 6732 9036
rect 6714 9036 6732 9054
rect 6714 9054 6732 9072
rect 6714 9072 6732 9090
rect 6714 9090 6732 9108
rect 6714 9108 6732 9126
rect 6714 9126 6732 9144
rect 6714 9144 6732 9162
rect 6714 9162 6732 9180
rect 6714 9180 6732 9198
rect 6714 9198 6732 9216
rect 6714 9216 6732 9234
rect 6714 9234 6732 9252
rect 6714 9252 6732 9270
rect 6714 9270 6732 9288
rect 6714 9288 6732 9306
rect 6714 9306 6732 9324
rect 6714 9324 6732 9342
rect 6714 9342 6732 9360
rect 6714 9360 6732 9378
rect 6714 9378 6732 9396
rect 6714 9396 6732 9414
rect 6714 9414 6732 9432
rect 6714 9432 6732 9450
rect 6714 9450 6732 9468
rect 6714 9468 6732 9486
rect 6714 9486 6732 9504
rect 6714 9504 6732 9522
rect 6714 9522 6732 9540
rect 6714 9540 6732 9558
rect 6714 9558 6732 9576
rect 6714 9576 6732 9594
rect 6714 9594 6732 9612
rect 6714 9612 6732 9630
rect 6714 9630 6732 9648
rect 6714 9648 6732 9666
rect 6714 9666 6732 9684
rect 6714 9684 6732 9702
rect 6714 9702 6732 9720
rect 6714 9720 6732 9738
rect 6714 9738 6732 9756
rect 6714 9756 6732 9774
rect 6714 9774 6732 9792
rect 6714 9792 6732 9810
rect 6714 9810 6732 9828
rect 6714 9828 6732 9846
rect 6714 9846 6732 9864
rect 6714 9864 6732 9882
rect 6714 9882 6732 9900
rect 6714 9900 6732 9918
rect 6714 9918 6732 9936
rect 6714 9936 6732 9954
rect 6714 9954 6732 9972
rect 6714 9972 6732 9990
rect 6714 9990 6732 10008
rect 6714 10008 6732 10026
rect 6714 10026 6732 10044
rect 6714 10044 6732 10062
rect 6714 10062 6732 10080
rect 6714 10080 6732 10098
rect 6714 10098 6732 10116
rect 6714 10116 6732 10134
rect 6732 1620 6750 1638
rect 6732 1638 6750 1656
rect 6732 1656 6750 1674
rect 6732 1674 6750 1692
rect 6732 1692 6750 1710
rect 6732 1710 6750 1728
rect 6732 1728 6750 1746
rect 6732 1746 6750 1764
rect 6732 1764 6750 1782
rect 6732 1782 6750 1800
rect 6732 1800 6750 1818
rect 6732 1818 6750 1836
rect 6732 1836 6750 1854
rect 6732 1854 6750 1872
rect 6732 1872 6750 1890
rect 6732 1890 6750 1908
rect 6732 1908 6750 1926
rect 6732 1926 6750 1944
rect 6732 1944 6750 1962
rect 6732 1962 6750 1980
rect 6732 1980 6750 1998
rect 6732 1998 6750 2016
rect 6732 2016 6750 2034
rect 6732 2034 6750 2052
rect 6732 2052 6750 2070
rect 6732 2070 6750 2088
rect 6732 2088 6750 2106
rect 6732 2106 6750 2124
rect 6732 2124 6750 2142
rect 6732 2142 6750 2160
rect 6732 2160 6750 2178
rect 6732 2178 6750 2196
rect 6732 2196 6750 2214
rect 6732 2214 6750 2232
rect 6732 2232 6750 2250
rect 6732 2250 6750 2268
rect 6732 2268 6750 2286
rect 6732 2286 6750 2304
rect 6732 2304 6750 2322
rect 6732 2322 6750 2340
rect 6732 2340 6750 2358
rect 6732 2358 6750 2376
rect 6732 2376 6750 2394
rect 6732 2394 6750 2412
rect 6732 2412 6750 2430
rect 6732 2430 6750 2448
rect 6732 2448 6750 2466
rect 6732 2466 6750 2484
rect 6732 2484 6750 2502
rect 6732 2502 6750 2520
rect 6732 2520 6750 2538
rect 6732 2538 6750 2556
rect 6732 2556 6750 2574
rect 6732 2574 6750 2592
rect 6732 2592 6750 2610
rect 6732 2610 6750 2628
rect 6732 2628 6750 2646
rect 6732 2646 6750 2664
rect 6732 2664 6750 2682
rect 6732 2682 6750 2700
rect 6732 2700 6750 2718
rect 6732 2718 6750 2736
rect 6732 2736 6750 2754
rect 6732 2754 6750 2772
rect 6732 2772 6750 2790
rect 6732 2790 6750 2808
rect 6732 2808 6750 2826
rect 6732 2826 6750 2844
rect 6732 2844 6750 2862
rect 6732 2862 6750 2880
rect 6732 2880 6750 2898
rect 6732 2898 6750 2916
rect 6732 2916 6750 2934
rect 6732 2934 6750 2952
rect 6732 2952 6750 2970
rect 6732 2970 6750 2988
rect 6732 2988 6750 3006
rect 6732 3168 6750 3186
rect 6732 3186 6750 3204
rect 6732 3204 6750 3222
rect 6732 3222 6750 3240
rect 6732 3240 6750 3258
rect 6732 3258 6750 3276
rect 6732 3276 6750 3294
rect 6732 3294 6750 3312
rect 6732 3312 6750 3330
rect 6732 3330 6750 3348
rect 6732 3348 6750 3366
rect 6732 3366 6750 3384
rect 6732 3384 6750 3402
rect 6732 3402 6750 3420
rect 6732 3420 6750 3438
rect 6732 3438 6750 3456
rect 6732 3456 6750 3474
rect 6732 3474 6750 3492
rect 6732 3492 6750 3510
rect 6732 3690 6750 3708
rect 6732 3708 6750 3726
rect 6732 3726 6750 3744
rect 6732 3744 6750 3762
rect 6732 3762 6750 3780
rect 6732 3780 6750 3798
rect 6732 3798 6750 3816
rect 6732 3816 6750 3834
rect 6732 3834 6750 3852
rect 6732 3852 6750 3870
rect 6732 3870 6750 3888
rect 6732 3888 6750 3906
rect 6732 3906 6750 3924
rect 6732 3924 6750 3942
rect 6732 3942 6750 3960
rect 6732 3960 6750 3978
rect 6732 3978 6750 3996
rect 6732 3996 6750 4014
rect 6732 4014 6750 4032
rect 6732 4032 6750 4050
rect 6732 4050 6750 4068
rect 6732 4068 6750 4086
rect 6732 4086 6750 4104
rect 6732 4104 6750 4122
rect 6732 4122 6750 4140
rect 6732 4140 6750 4158
rect 6732 4158 6750 4176
rect 6732 4176 6750 4194
rect 6732 4194 6750 4212
rect 6732 4212 6750 4230
rect 6732 4230 6750 4248
rect 6732 4248 6750 4266
rect 6732 4266 6750 4284
rect 6732 4284 6750 4302
rect 6732 4302 6750 4320
rect 6732 4320 6750 4338
rect 6732 4338 6750 4356
rect 6732 4356 6750 4374
rect 6732 4374 6750 4392
rect 6732 4392 6750 4410
rect 6732 4410 6750 4428
rect 6732 4428 6750 4446
rect 6732 4446 6750 4464
rect 6732 4464 6750 4482
rect 6732 4482 6750 4500
rect 6732 4500 6750 4518
rect 6732 4518 6750 4536
rect 6732 4536 6750 4554
rect 6732 4554 6750 4572
rect 6732 4572 6750 4590
rect 6732 4590 6750 4608
rect 6732 4608 6750 4626
rect 6732 4626 6750 4644
rect 6732 4644 6750 4662
rect 6732 4662 6750 4680
rect 6732 4680 6750 4698
rect 6732 4698 6750 4716
rect 6732 4716 6750 4734
rect 6732 4734 6750 4752
rect 6732 4752 6750 4770
rect 6732 4770 6750 4788
rect 6732 4788 6750 4806
rect 6732 4806 6750 4824
rect 6732 4824 6750 4842
rect 6732 4842 6750 4860
rect 6732 4860 6750 4878
rect 6732 4878 6750 4896
rect 6732 4896 6750 4914
rect 6732 4914 6750 4932
rect 6732 4932 6750 4950
rect 6732 4950 6750 4968
rect 6732 4968 6750 4986
rect 6732 4986 6750 5004
rect 6732 5004 6750 5022
rect 6732 5022 6750 5040
rect 6732 5040 6750 5058
rect 6732 5058 6750 5076
rect 6732 5076 6750 5094
rect 6732 5094 6750 5112
rect 6732 5112 6750 5130
rect 6732 5130 6750 5148
rect 6732 5148 6750 5166
rect 6732 5166 6750 5184
rect 6732 5184 6750 5202
rect 6732 5202 6750 5220
rect 6732 5220 6750 5238
rect 6732 5238 6750 5256
rect 6732 5256 6750 5274
rect 6732 5274 6750 5292
rect 6732 5292 6750 5310
rect 6732 5310 6750 5328
rect 6732 5328 6750 5346
rect 6732 5346 6750 5364
rect 6732 5364 6750 5382
rect 6732 5382 6750 5400
rect 6732 5400 6750 5418
rect 6732 5418 6750 5436
rect 6732 5436 6750 5454
rect 6732 5454 6750 5472
rect 6732 5472 6750 5490
rect 6732 5490 6750 5508
rect 6732 5508 6750 5526
rect 6732 5526 6750 5544
rect 6732 5544 6750 5562
rect 6732 5562 6750 5580
rect 6732 5580 6750 5598
rect 6732 5598 6750 5616
rect 6732 5616 6750 5634
rect 6732 5634 6750 5652
rect 6732 5652 6750 5670
rect 6732 5670 6750 5688
rect 6732 5688 6750 5706
rect 6732 5706 6750 5724
rect 6732 5724 6750 5742
rect 6732 5742 6750 5760
rect 6732 5760 6750 5778
rect 6732 5778 6750 5796
rect 6732 5796 6750 5814
rect 6732 5814 6750 5832
rect 6732 5832 6750 5850
rect 6732 5850 6750 5868
rect 6732 5868 6750 5886
rect 6732 5886 6750 5904
rect 6732 5904 6750 5922
rect 6732 5922 6750 5940
rect 6732 5940 6750 5958
rect 6732 5958 6750 5976
rect 6732 5976 6750 5994
rect 6732 5994 6750 6012
rect 6732 6012 6750 6030
rect 6732 7164 6750 7182
rect 6732 7182 6750 7200
rect 6732 7200 6750 7218
rect 6732 7218 6750 7236
rect 6732 7236 6750 7254
rect 6732 7254 6750 7272
rect 6732 7272 6750 7290
rect 6732 7290 6750 7308
rect 6732 7308 6750 7326
rect 6732 7326 6750 7344
rect 6732 7344 6750 7362
rect 6732 7362 6750 7380
rect 6732 7380 6750 7398
rect 6732 7398 6750 7416
rect 6732 7416 6750 7434
rect 6732 7434 6750 7452
rect 6732 7452 6750 7470
rect 6732 7470 6750 7488
rect 6732 7488 6750 7506
rect 6732 7506 6750 7524
rect 6732 7524 6750 7542
rect 6732 7542 6750 7560
rect 6732 7560 6750 7578
rect 6732 7578 6750 7596
rect 6732 7596 6750 7614
rect 6732 7614 6750 7632
rect 6732 7632 6750 7650
rect 6732 7650 6750 7668
rect 6732 7668 6750 7686
rect 6732 7686 6750 7704
rect 6732 7704 6750 7722
rect 6732 7722 6750 7740
rect 6732 7740 6750 7758
rect 6732 7758 6750 7776
rect 6732 7776 6750 7794
rect 6732 7794 6750 7812
rect 6732 7812 6750 7830
rect 6732 7830 6750 7848
rect 6732 7848 6750 7866
rect 6732 7866 6750 7884
rect 6732 7884 6750 7902
rect 6732 7902 6750 7920
rect 6732 7920 6750 7938
rect 6732 7938 6750 7956
rect 6732 7956 6750 7974
rect 6732 7974 6750 7992
rect 6732 7992 6750 8010
rect 6732 8010 6750 8028
rect 6732 8028 6750 8046
rect 6732 8046 6750 8064
rect 6732 8064 6750 8082
rect 6732 8082 6750 8100
rect 6732 8100 6750 8118
rect 6732 8118 6750 8136
rect 6732 8136 6750 8154
rect 6732 8154 6750 8172
rect 6732 8172 6750 8190
rect 6732 8190 6750 8208
rect 6732 8208 6750 8226
rect 6732 8226 6750 8244
rect 6732 8244 6750 8262
rect 6732 8262 6750 8280
rect 6732 8280 6750 8298
rect 6732 8298 6750 8316
rect 6732 8316 6750 8334
rect 6732 8334 6750 8352
rect 6732 8352 6750 8370
rect 6732 8370 6750 8388
rect 6732 8388 6750 8406
rect 6732 8406 6750 8424
rect 6732 8424 6750 8442
rect 6732 8442 6750 8460
rect 6732 8460 6750 8478
rect 6732 8478 6750 8496
rect 6732 8496 6750 8514
rect 6732 8514 6750 8532
rect 6732 8532 6750 8550
rect 6732 8550 6750 8568
rect 6732 8568 6750 8586
rect 6732 8586 6750 8604
rect 6732 8604 6750 8622
rect 6732 8622 6750 8640
rect 6732 8640 6750 8658
rect 6732 8658 6750 8676
rect 6732 8676 6750 8694
rect 6732 8694 6750 8712
rect 6732 8712 6750 8730
rect 6732 8730 6750 8748
rect 6732 8748 6750 8766
rect 6732 8766 6750 8784
rect 6732 8784 6750 8802
rect 6732 8802 6750 8820
rect 6732 8820 6750 8838
rect 6732 8838 6750 8856
rect 6732 8856 6750 8874
rect 6732 8874 6750 8892
rect 6732 8892 6750 8910
rect 6732 8910 6750 8928
rect 6732 8928 6750 8946
rect 6732 8946 6750 8964
rect 6732 8964 6750 8982
rect 6732 8982 6750 9000
rect 6732 9000 6750 9018
rect 6732 9018 6750 9036
rect 6732 9036 6750 9054
rect 6732 9054 6750 9072
rect 6732 9072 6750 9090
rect 6732 9090 6750 9108
rect 6732 9108 6750 9126
rect 6732 9126 6750 9144
rect 6732 9144 6750 9162
rect 6732 9162 6750 9180
rect 6732 9180 6750 9198
rect 6732 9198 6750 9216
rect 6732 9216 6750 9234
rect 6732 9234 6750 9252
rect 6732 9252 6750 9270
rect 6732 9270 6750 9288
rect 6732 9288 6750 9306
rect 6732 9306 6750 9324
rect 6732 9324 6750 9342
rect 6732 9342 6750 9360
rect 6732 9360 6750 9378
rect 6732 9378 6750 9396
rect 6732 9396 6750 9414
rect 6732 9414 6750 9432
rect 6732 9432 6750 9450
rect 6732 9450 6750 9468
rect 6732 9468 6750 9486
rect 6732 9486 6750 9504
rect 6732 9504 6750 9522
rect 6732 9522 6750 9540
rect 6732 9540 6750 9558
rect 6732 9558 6750 9576
rect 6732 9576 6750 9594
rect 6732 9594 6750 9612
rect 6732 9612 6750 9630
rect 6732 9630 6750 9648
rect 6732 9648 6750 9666
rect 6732 9666 6750 9684
rect 6732 9684 6750 9702
rect 6732 9702 6750 9720
rect 6732 9720 6750 9738
rect 6732 9738 6750 9756
rect 6732 9756 6750 9774
rect 6732 9774 6750 9792
rect 6732 9792 6750 9810
rect 6732 9810 6750 9828
rect 6732 9828 6750 9846
rect 6732 9846 6750 9864
rect 6732 9864 6750 9882
rect 6732 9882 6750 9900
rect 6732 9900 6750 9918
rect 6732 9918 6750 9936
rect 6732 9936 6750 9954
rect 6732 9954 6750 9972
rect 6732 9972 6750 9990
rect 6732 9990 6750 10008
rect 6732 10008 6750 10026
rect 6732 10026 6750 10044
rect 6732 10044 6750 10062
rect 6732 10062 6750 10080
rect 6732 10080 6750 10098
rect 6732 10098 6750 10116
rect 6732 10116 6750 10134
rect 6732 10134 6750 10152
rect 6750 1638 6768 1656
rect 6750 1656 6768 1674
rect 6750 1674 6768 1692
rect 6750 1692 6768 1710
rect 6750 1710 6768 1728
rect 6750 1728 6768 1746
rect 6750 1746 6768 1764
rect 6750 1764 6768 1782
rect 6750 1782 6768 1800
rect 6750 1800 6768 1818
rect 6750 1818 6768 1836
rect 6750 1836 6768 1854
rect 6750 1854 6768 1872
rect 6750 1872 6768 1890
rect 6750 1890 6768 1908
rect 6750 1908 6768 1926
rect 6750 1926 6768 1944
rect 6750 1944 6768 1962
rect 6750 1962 6768 1980
rect 6750 1980 6768 1998
rect 6750 1998 6768 2016
rect 6750 2016 6768 2034
rect 6750 2034 6768 2052
rect 6750 2052 6768 2070
rect 6750 2070 6768 2088
rect 6750 2088 6768 2106
rect 6750 2106 6768 2124
rect 6750 2124 6768 2142
rect 6750 2142 6768 2160
rect 6750 2160 6768 2178
rect 6750 2178 6768 2196
rect 6750 2196 6768 2214
rect 6750 2214 6768 2232
rect 6750 2232 6768 2250
rect 6750 2250 6768 2268
rect 6750 2268 6768 2286
rect 6750 2286 6768 2304
rect 6750 2304 6768 2322
rect 6750 2322 6768 2340
rect 6750 2340 6768 2358
rect 6750 2358 6768 2376
rect 6750 2376 6768 2394
rect 6750 2394 6768 2412
rect 6750 2412 6768 2430
rect 6750 2430 6768 2448
rect 6750 2448 6768 2466
rect 6750 2466 6768 2484
rect 6750 2484 6768 2502
rect 6750 2502 6768 2520
rect 6750 2520 6768 2538
rect 6750 2538 6768 2556
rect 6750 2556 6768 2574
rect 6750 2574 6768 2592
rect 6750 2592 6768 2610
rect 6750 2610 6768 2628
rect 6750 2628 6768 2646
rect 6750 2646 6768 2664
rect 6750 2664 6768 2682
rect 6750 2682 6768 2700
rect 6750 2700 6768 2718
rect 6750 2718 6768 2736
rect 6750 2736 6768 2754
rect 6750 2754 6768 2772
rect 6750 2772 6768 2790
rect 6750 2790 6768 2808
rect 6750 2808 6768 2826
rect 6750 2826 6768 2844
rect 6750 2844 6768 2862
rect 6750 2862 6768 2880
rect 6750 2880 6768 2898
rect 6750 2898 6768 2916
rect 6750 2916 6768 2934
rect 6750 2934 6768 2952
rect 6750 2952 6768 2970
rect 6750 2970 6768 2988
rect 6750 2988 6768 3006
rect 6750 3006 6768 3024
rect 6750 3186 6768 3204
rect 6750 3204 6768 3222
rect 6750 3222 6768 3240
rect 6750 3240 6768 3258
rect 6750 3258 6768 3276
rect 6750 3276 6768 3294
rect 6750 3294 6768 3312
rect 6750 3312 6768 3330
rect 6750 3330 6768 3348
rect 6750 3348 6768 3366
rect 6750 3366 6768 3384
rect 6750 3384 6768 3402
rect 6750 3402 6768 3420
rect 6750 3420 6768 3438
rect 6750 3438 6768 3456
rect 6750 3456 6768 3474
rect 6750 3474 6768 3492
rect 6750 3492 6768 3510
rect 6750 3510 6768 3528
rect 6750 3726 6768 3744
rect 6750 3744 6768 3762
rect 6750 3762 6768 3780
rect 6750 3780 6768 3798
rect 6750 3798 6768 3816
rect 6750 3816 6768 3834
rect 6750 3834 6768 3852
rect 6750 3852 6768 3870
rect 6750 3870 6768 3888
rect 6750 3888 6768 3906
rect 6750 3906 6768 3924
rect 6750 3924 6768 3942
rect 6750 3942 6768 3960
rect 6750 3960 6768 3978
rect 6750 3978 6768 3996
rect 6750 3996 6768 4014
rect 6750 4014 6768 4032
rect 6750 4032 6768 4050
rect 6750 4050 6768 4068
rect 6750 4068 6768 4086
rect 6750 4086 6768 4104
rect 6750 4104 6768 4122
rect 6750 4122 6768 4140
rect 6750 4140 6768 4158
rect 6750 4158 6768 4176
rect 6750 4176 6768 4194
rect 6750 4194 6768 4212
rect 6750 4212 6768 4230
rect 6750 4230 6768 4248
rect 6750 4248 6768 4266
rect 6750 4266 6768 4284
rect 6750 4284 6768 4302
rect 6750 4302 6768 4320
rect 6750 4320 6768 4338
rect 6750 4338 6768 4356
rect 6750 4356 6768 4374
rect 6750 4374 6768 4392
rect 6750 4392 6768 4410
rect 6750 4410 6768 4428
rect 6750 4428 6768 4446
rect 6750 4446 6768 4464
rect 6750 4464 6768 4482
rect 6750 4482 6768 4500
rect 6750 4500 6768 4518
rect 6750 4518 6768 4536
rect 6750 4536 6768 4554
rect 6750 4554 6768 4572
rect 6750 4572 6768 4590
rect 6750 4590 6768 4608
rect 6750 4608 6768 4626
rect 6750 4626 6768 4644
rect 6750 4644 6768 4662
rect 6750 4662 6768 4680
rect 6750 4680 6768 4698
rect 6750 4698 6768 4716
rect 6750 4716 6768 4734
rect 6750 4734 6768 4752
rect 6750 4752 6768 4770
rect 6750 4770 6768 4788
rect 6750 4788 6768 4806
rect 6750 4806 6768 4824
rect 6750 4824 6768 4842
rect 6750 4842 6768 4860
rect 6750 4860 6768 4878
rect 6750 4878 6768 4896
rect 6750 4896 6768 4914
rect 6750 4914 6768 4932
rect 6750 4932 6768 4950
rect 6750 4950 6768 4968
rect 6750 4968 6768 4986
rect 6750 4986 6768 5004
rect 6750 5004 6768 5022
rect 6750 5022 6768 5040
rect 6750 5040 6768 5058
rect 6750 5058 6768 5076
rect 6750 5076 6768 5094
rect 6750 5094 6768 5112
rect 6750 5112 6768 5130
rect 6750 5130 6768 5148
rect 6750 5148 6768 5166
rect 6750 5166 6768 5184
rect 6750 5184 6768 5202
rect 6750 5202 6768 5220
rect 6750 5220 6768 5238
rect 6750 5238 6768 5256
rect 6750 5256 6768 5274
rect 6750 5274 6768 5292
rect 6750 5292 6768 5310
rect 6750 5310 6768 5328
rect 6750 5328 6768 5346
rect 6750 5346 6768 5364
rect 6750 5364 6768 5382
rect 6750 5382 6768 5400
rect 6750 5400 6768 5418
rect 6750 5418 6768 5436
rect 6750 5436 6768 5454
rect 6750 5454 6768 5472
rect 6750 5472 6768 5490
rect 6750 5490 6768 5508
rect 6750 5508 6768 5526
rect 6750 5526 6768 5544
rect 6750 5544 6768 5562
rect 6750 5562 6768 5580
rect 6750 5580 6768 5598
rect 6750 5598 6768 5616
rect 6750 5616 6768 5634
rect 6750 5634 6768 5652
rect 6750 5652 6768 5670
rect 6750 5670 6768 5688
rect 6750 5688 6768 5706
rect 6750 5706 6768 5724
rect 6750 5724 6768 5742
rect 6750 5742 6768 5760
rect 6750 5760 6768 5778
rect 6750 5778 6768 5796
rect 6750 5796 6768 5814
rect 6750 5814 6768 5832
rect 6750 5832 6768 5850
rect 6750 5850 6768 5868
rect 6750 5868 6768 5886
rect 6750 5886 6768 5904
rect 6750 5904 6768 5922
rect 6750 5922 6768 5940
rect 6750 5940 6768 5958
rect 6750 5958 6768 5976
rect 6750 5976 6768 5994
rect 6750 5994 6768 6012
rect 6750 6012 6768 6030
rect 6750 6030 6768 6048
rect 6750 7200 6768 7218
rect 6750 7218 6768 7236
rect 6750 7236 6768 7254
rect 6750 7254 6768 7272
rect 6750 7272 6768 7290
rect 6750 7290 6768 7308
rect 6750 7308 6768 7326
rect 6750 7326 6768 7344
rect 6750 7344 6768 7362
rect 6750 7362 6768 7380
rect 6750 7380 6768 7398
rect 6750 7398 6768 7416
rect 6750 7416 6768 7434
rect 6750 7434 6768 7452
rect 6750 7452 6768 7470
rect 6750 7470 6768 7488
rect 6750 7488 6768 7506
rect 6750 7506 6768 7524
rect 6750 7524 6768 7542
rect 6750 7542 6768 7560
rect 6750 7560 6768 7578
rect 6750 7578 6768 7596
rect 6750 7596 6768 7614
rect 6750 7614 6768 7632
rect 6750 7632 6768 7650
rect 6750 7650 6768 7668
rect 6750 7668 6768 7686
rect 6750 7686 6768 7704
rect 6750 7704 6768 7722
rect 6750 7722 6768 7740
rect 6750 7740 6768 7758
rect 6750 7758 6768 7776
rect 6750 7776 6768 7794
rect 6750 7794 6768 7812
rect 6750 7812 6768 7830
rect 6750 7830 6768 7848
rect 6750 7848 6768 7866
rect 6750 7866 6768 7884
rect 6750 7884 6768 7902
rect 6750 7902 6768 7920
rect 6750 7920 6768 7938
rect 6750 7938 6768 7956
rect 6750 7956 6768 7974
rect 6750 7974 6768 7992
rect 6750 7992 6768 8010
rect 6750 8010 6768 8028
rect 6750 8028 6768 8046
rect 6750 8046 6768 8064
rect 6750 8064 6768 8082
rect 6750 8082 6768 8100
rect 6750 8100 6768 8118
rect 6750 8118 6768 8136
rect 6750 8136 6768 8154
rect 6750 8154 6768 8172
rect 6750 8172 6768 8190
rect 6750 8190 6768 8208
rect 6750 8208 6768 8226
rect 6750 8226 6768 8244
rect 6750 8244 6768 8262
rect 6750 8262 6768 8280
rect 6750 8280 6768 8298
rect 6750 8298 6768 8316
rect 6750 8316 6768 8334
rect 6750 8334 6768 8352
rect 6750 8352 6768 8370
rect 6750 8370 6768 8388
rect 6750 8388 6768 8406
rect 6750 8406 6768 8424
rect 6750 8424 6768 8442
rect 6750 8442 6768 8460
rect 6750 8460 6768 8478
rect 6750 8478 6768 8496
rect 6750 8496 6768 8514
rect 6750 8514 6768 8532
rect 6750 8532 6768 8550
rect 6750 8550 6768 8568
rect 6750 8568 6768 8586
rect 6750 8586 6768 8604
rect 6750 8604 6768 8622
rect 6750 8622 6768 8640
rect 6750 8640 6768 8658
rect 6750 8658 6768 8676
rect 6750 8676 6768 8694
rect 6750 8694 6768 8712
rect 6750 8712 6768 8730
rect 6750 8730 6768 8748
rect 6750 8748 6768 8766
rect 6750 8766 6768 8784
rect 6750 8784 6768 8802
rect 6750 8802 6768 8820
rect 6750 8820 6768 8838
rect 6750 8838 6768 8856
rect 6750 8856 6768 8874
rect 6750 8874 6768 8892
rect 6750 8892 6768 8910
rect 6750 8910 6768 8928
rect 6750 8928 6768 8946
rect 6750 8946 6768 8964
rect 6750 8964 6768 8982
rect 6750 8982 6768 9000
rect 6750 9000 6768 9018
rect 6750 9018 6768 9036
rect 6750 9036 6768 9054
rect 6750 9054 6768 9072
rect 6750 9072 6768 9090
rect 6750 9090 6768 9108
rect 6750 9108 6768 9126
rect 6750 9126 6768 9144
rect 6750 9144 6768 9162
rect 6750 9162 6768 9180
rect 6750 9180 6768 9198
rect 6750 9198 6768 9216
rect 6750 9216 6768 9234
rect 6750 9234 6768 9252
rect 6750 9252 6768 9270
rect 6750 9270 6768 9288
rect 6750 9288 6768 9306
rect 6750 9306 6768 9324
rect 6750 9324 6768 9342
rect 6750 9342 6768 9360
rect 6750 9360 6768 9378
rect 6750 9378 6768 9396
rect 6750 9396 6768 9414
rect 6750 9414 6768 9432
rect 6750 9432 6768 9450
rect 6750 9450 6768 9468
rect 6750 9468 6768 9486
rect 6750 9486 6768 9504
rect 6750 9504 6768 9522
rect 6750 9522 6768 9540
rect 6750 9540 6768 9558
rect 6750 9558 6768 9576
rect 6750 9576 6768 9594
rect 6750 9594 6768 9612
rect 6750 9612 6768 9630
rect 6750 9630 6768 9648
rect 6750 9648 6768 9666
rect 6750 9666 6768 9684
rect 6750 9684 6768 9702
rect 6750 9702 6768 9720
rect 6750 9720 6768 9738
rect 6750 9738 6768 9756
rect 6750 9756 6768 9774
rect 6750 9774 6768 9792
rect 6750 9792 6768 9810
rect 6750 9810 6768 9828
rect 6750 9828 6768 9846
rect 6750 9846 6768 9864
rect 6750 9864 6768 9882
rect 6750 9882 6768 9900
rect 6750 9900 6768 9918
rect 6750 9918 6768 9936
rect 6750 9936 6768 9954
rect 6750 9954 6768 9972
rect 6750 9972 6768 9990
rect 6750 9990 6768 10008
rect 6750 10008 6768 10026
rect 6750 10026 6768 10044
rect 6750 10044 6768 10062
rect 6750 10062 6768 10080
rect 6750 10080 6768 10098
rect 6750 10098 6768 10116
rect 6750 10116 6768 10134
rect 6750 10134 6768 10152
rect 6750 10152 6768 10170
rect 6768 1656 6786 1674
rect 6768 1674 6786 1692
rect 6768 1692 6786 1710
rect 6768 1710 6786 1728
rect 6768 1728 6786 1746
rect 6768 1746 6786 1764
rect 6768 1764 6786 1782
rect 6768 1782 6786 1800
rect 6768 1800 6786 1818
rect 6768 1818 6786 1836
rect 6768 1836 6786 1854
rect 6768 1854 6786 1872
rect 6768 1872 6786 1890
rect 6768 1890 6786 1908
rect 6768 1908 6786 1926
rect 6768 1926 6786 1944
rect 6768 1944 6786 1962
rect 6768 1962 6786 1980
rect 6768 1980 6786 1998
rect 6768 1998 6786 2016
rect 6768 2016 6786 2034
rect 6768 2034 6786 2052
rect 6768 2052 6786 2070
rect 6768 2070 6786 2088
rect 6768 2088 6786 2106
rect 6768 2106 6786 2124
rect 6768 2124 6786 2142
rect 6768 2142 6786 2160
rect 6768 2160 6786 2178
rect 6768 2178 6786 2196
rect 6768 2196 6786 2214
rect 6768 2214 6786 2232
rect 6768 2232 6786 2250
rect 6768 2250 6786 2268
rect 6768 2268 6786 2286
rect 6768 2286 6786 2304
rect 6768 2304 6786 2322
rect 6768 2322 6786 2340
rect 6768 2340 6786 2358
rect 6768 2358 6786 2376
rect 6768 2376 6786 2394
rect 6768 2394 6786 2412
rect 6768 2412 6786 2430
rect 6768 2430 6786 2448
rect 6768 2448 6786 2466
rect 6768 2466 6786 2484
rect 6768 2484 6786 2502
rect 6768 2502 6786 2520
rect 6768 2520 6786 2538
rect 6768 2538 6786 2556
rect 6768 2556 6786 2574
rect 6768 2574 6786 2592
rect 6768 2592 6786 2610
rect 6768 2610 6786 2628
rect 6768 2628 6786 2646
rect 6768 2646 6786 2664
rect 6768 2664 6786 2682
rect 6768 2682 6786 2700
rect 6768 2700 6786 2718
rect 6768 2718 6786 2736
rect 6768 2736 6786 2754
rect 6768 2754 6786 2772
rect 6768 2772 6786 2790
rect 6768 2790 6786 2808
rect 6768 2808 6786 2826
rect 6768 2826 6786 2844
rect 6768 2844 6786 2862
rect 6768 2862 6786 2880
rect 6768 2880 6786 2898
rect 6768 2898 6786 2916
rect 6768 2916 6786 2934
rect 6768 2934 6786 2952
rect 6768 2952 6786 2970
rect 6768 2970 6786 2988
rect 6768 2988 6786 3006
rect 6768 3006 6786 3024
rect 6768 3186 6786 3204
rect 6768 3204 6786 3222
rect 6768 3222 6786 3240
rect 6768 3240 6786 3258
rect 6768 3258 6786 3276
rect 6768 3276 6786 3294
rect 6768 3294 6786 3312
rect 6768 3312 6786 3330
rect 6768 3330 6786 3348
rect 6768 3348 6786 3366
rect 6768 3366 6786 3384
rect 6768 3384 6786 3402
rect 6768 3402 6786 3420
rect 6768 3420 6786 3438
rect 6768 3438 6786 3456
rect 6768 3456 6786 3474
rect 6768 3474 6786 3492
rect 6768 3492 6786 3510
rect 6768 3510 6786 3528
rect 6768 3528 6786 3546
rect 6768 3744 6786 3762
rect 6768 3762 6786 3780
rect 6768 3780 6786 3798
rect 6768 3798 6786 3816
rect 6768 3816 6786 3834
rect 6768 3834 6786 3852
rect 6768 3852 6786 3870
rect 6768 3870 6786 3888
rect 6768 3888 6786 3906
rect 6768 3906 6786 3924
rect 6768 3924 6786 3942
rect 6768 3942 6786 3960
rect 6768 3960 6786 3978
rect 6768 3978 6786 3996
rect 6768 3996 6786 4014
rect 6768 4014 6786 4032
rect 6768 4032 6786 4050
rect 6768 4050 6786 4068
rect 6768 4068 6786 4086
rect 6768 4086 6786 4104
rect 6768 4104 6786 4122
rect 6768 4122 6786 4140
rect 6768 4140 6786 4158
rect 6768 4158 6786 4176
rect 6768 4176 6786 4194
rect 6768 4194 6786 4212
rect 6768 4212 6786 4230
rect 6768 4230 6786 4248
rect 6768 4248 6786 4266
rect 6768 4266 6786 4284
rect 6768 4284 6786 4302
rect 6768 4302 6786 4320
rect 6768 4320 6786 4338
rect 6768 4338 6786 4356
rect 6768 4356 6786 4374
rect 6768 4374 6786 4392
rect 6768 4392 6786 4410
rect 6768 4410 6786 4428
rect 6768 4428 6786 4446
rect 6768 4446 6786 4464
rect 6768 4464 6786 4482
rect 6768 4482 6786 4500
rect 6768 4500 6786 4518
rect 6768 4518 6786 4536
rect 6768 4536 6786 4554
rect 6768 4554 6786 4572
rect 6768 4572 6786 4590
rect 6768 4590 6786 4608
rect 6768 4608 6786 4626
rect 6768 4626 6786 4644
rect 6768 4644 6786 4662
rect 6768 4662 6786 4680
rect 6768 4680 6786 4698
rect 6768 4698 6786 4716
rect 6768 4716 6786 4734
rect 6768 4734 6786 4752
rect 6768 4752 6786 4770
rect 6768 4770 6786 4788
rect 6768 4788 6786 4806
rect 6768 4806 6786 4824
rect 6768 4824 6786 4842
rect 6768 4842 6786 4860
rect 6768 4860 6786 4878
rect 6768 4878 6786 4896
rect 6768 4896 6786 4914
rect 6768 4914 6786 4932
rect 6768 4932 6786 4950
rect 6768 4950 6786 4968
rect 6768 4968 6786 4986
rect 6768 4986 6786 5004
rect 6768 5004 6786 5022
rect 6768 5022 6786 5040
rect 6768 5040 6786 5058
rect 6768 5058 6786 5076
rect 6768 5076 6786 5094
rect 6768 5094 6786 5112
rect 6768 5112 6786 5130
rect 6768 5130 6786 5148
rect 6768 5148 6786 5166
rect 6768 5166 6786 5184
rect 6768 5184 6786 5202
rect 6768 5202 6786 5220
rect 6768 5220 6786 5238
rect 6768 5238 6786 5256
rect 6768 5256 6786 5274
rect 6768 5274 6786 5292
rect 6768 5292 6786 5310
rect 6768 5310 6786 5328
rect 6768 5328 6786 5346
rect 6768 5346 6786 5364
rect 6768 5364 6786 5382
rect 6768 5382 6786 5400
rect 6768 5400 6786 5418
rect 6768 5418 6786 5436
rect 6768 5436 6786 5454
rect 6768 5454 6786 5472
rect 6768 5472 6786 5490
rect 6768 5490 6786 5508
rect 6768 5508 6786 5526
rect 6768 5526 6786 5544
rect 6768 5544 6786 5562
rect 6768 5562 6786 5580
rect 6768 5580 6786 5598
rect 6768 5598 6786 5616
rect 6768 5616 6786 5634
rect 6768 5634 6786 5652
rect 6768 5652 6786 5670
rect 6768 5670 6786 5688
rect 6768 5688 6786 5706
rect 6768 5706 6786 5724
rect 6768 5724 6786 5742
rect 6768 5742 6786 5760
rect 6768 5760 6786 5778
rect 6768 5778 6786 5796
rect 6768 5796 6786 5814
rect 6768 5814 6786 5832
rect 6768 5832 6786 5850
rect 6768 5850 6786 5868
rect 6768 5868 6786 5886
rect 6768 5886 6786 5904
rect 6768 5904 6786 5922
rect 6768 5922 6786 5940
rect 6768 5940 6786 5958
rect 6768 5958 6786 5976
rect 6768 5976 6786 5994
rect 6768 5994 6786 6012
rect 6768 6012 6786 6030
rect 6768 6030 6786 6048
rect 6768 6048 6786 6066
rect 6768 7254 6786 7272
rect 6768 7272 6786 7290
rect 6768 7290 6786 7308
rect 6768 7308 6786 7326
rect 6768 7326 6786 7344
rect 6768 7344 6786 7362
rect 6768 7362 6786 7380
rect 6768 7380 6786 7398
rect 6768 7398 6786 7416
rect 6768 7416 6786 7434
rect 6768 7434 6786 7452
rect 6768 7452 6786 7470
rect 6768 7470 6786 7488
rect 6768 7488 6786 7506
rect 6768 7506 6786 7524
rect 6768 7524 6786 7542
rect 6768 7542 6786 7560
rect 6768 7560 6786 7578
rect 6768 7578 6786 7596
rect 6768 7596 6786 7614
rect 6768 7614 6786 7632
rect 6768 7632 6786 7650
rect 6768 7650 6786 7668
rect 6768 7668 6786 7686
rect 6768 7686 6786 7704
rect 6768 7704 6786 7722
rect 6768 7722 6786 7740
rect 6768 7740 6786 7758
rect 6768 7758 6786 7776
rect 6768 7776 6786 7794
rect 6768 7794 6786 7812
rect 6768 7812 6786 7830
rect 6768 7830 6786 7848
rect 6768 7848 6786 7866
rect 6768 7866 6786 7884
rect 6768 7884 6786 7902
rect 6768 7902 6786 7920
rect 6768 7920 6786 7938
rect 6768 7938 6786 7956
rect 6768 7956 6786 7974
rect 6768 7974 6786 7992
rect 6768 7992 6786 8010
rect 6768 8010 6786 8028
rect 6768 8028 6786 8046
rect 6768 8046 6786 8064
rect 6768 8064 6786 8082
rect 6768 8082 6786 8100
rect 6768 8100 6786 8118
rect 6768 8118 6786 8136
rect 6768 8136 6786 8154
rect 6768 8154 6786 8172
rect 6768 8172 6786 8190
rect 6768 8190 6786 8208
rect 6768 8208 6786 8226
rect 6768 8226 6786 8244
rect 6768 8244 6786 8262
rect 6768 8262 6786 8280
rect 6768 8280 6786 8298
rect 6768 8298 6786 8316
rect 6768 8316 6786 8334
rect 6768 8334 6786 8352
rect 6768 8352 6786 8370
rect 6768 8370 6786 8388
rect 6768 8388 6786 8406
rect 6768 8406 6786 8424
rect 6768 8424 6786 8442
rect 6768 8442 6786 8460
rect 6768 8460 6786 8478
rect 6768 8478 6786 8496
rect 6768 8496 6786 8514
rect 6768 8514 6786 8532
rect 6768 8532 6786 8550
rect 6768 8550 6786 8568
rect 6768 8568 6786 8586
rect 6768 8586 6786 8604
rect 6768 8604 6786 8622
rect 6768 8622 6786 8640
rect 6768 8640 6786 8658
rect 6768 8658 6786 8676
rect 6768 8676 6786 8694
rect 6768 8694 6786 8712
rect 6768 8712 6786 8730
rect 6768 8730 6786 8748
rect 6768 8748 6786 8766
rect 6768 8766 6786 8784
rect 6768 8784 6786 8802
rect 6768 8802 6786 8820
rect 6768 8820 6786 8838
rect 6768 8838 6786 8856
rect 6768 8856 6786 8874
rect 6768 8874 6786 8892
rect 6768 8892 6786 8910
rect 6768 8910 6786 8928
rect 6768 8928 6786 8946
rect 6768 8946 6786 8964
rect 6768 8964 6786 8982
rect 6768 8982 6786 9000
rect 6768 9000 6786 9018
rect 6768 9018 6786 9036
rect 6768 9036 6786 9054
rect 6768 9054 6786 9072
rect 6768 9072 6786 9090
rect 6768 9090 6786 9108
rect 6768 9108 6786 9126
rect 6768 9126 6786 9144
rect 6768 9144 6786 9162
rect 6768 9162 6786 9180
rect 6768 9180 6786 9198
rect 6768 9198 6786 9216
rect 6768 9216 6786 9234
rect 6768 9234 6786 9252
rect 6768 9252 6786 9270
rect 6768 9270 6786 9288
rect 6768 9288 6786 9306
rect 6768 9306 6786 9324
rect 6768 9324 6786 9342
rect 6768 9342 6786 9360
rect 6768 9360 6786 9378
rect 6768 9378 6786 9396
rect 6768 9396 6786 9414
rect 6768 9414 6786 9432
rect 6768 9432 6786 9450
rect 6768 9450 6786 9468
rect 6768 9468 6786 9486
rect 6768 9486 6786 9504
rect 6768 9504 6786 9522
rect 6768 9522 6786 9540
rect 6768 9540 6786 9558
rect 6768 9558 6786 9576
rect 6768 9576 6786 9594
rect 6768 9594 6786 9612
rect 6768 9612 6786 9630
rect 6768 9630 6786 9648
rect 6768 9648 6786 9666
rect 6768 9666 6786 9684
rect 6768 9684 6786 9702
rect 6768 9702 6786 9720
rect 6768 9720 6786 9738
rect 6768 9738 6786 9756
rect 6768 9756 6786 9774
rect 6768 9774 6786 9792
rect 6768 9792 6786 9810
rect 6768 9810 6786 9828
rect 6768 9828 6786 9846
rect 6768 9846 6786 9864
rect 6768 9864 6786 9882
rect 6768 9882 6786 9900
rect 6768 9900 6786 9918
rect 6768 9918 6786 9936
rect 6768 9936 6786 9954
rect 6768 9954 6786 9972
rect 6768 9972 6786 9990
rect 6768 9990 6786 10008
rect 6768 10008 6786 10026
rect 6768 10026 6786 10044
rect 6768 10044 6786 10062
rect 6768 10062 6786 10080
rect 6768 10080 6786 10098
rect 6768 10098 6786 10116
rect 6768 10116 6786 10134
rect 6768 10134 6786 10152
rect 6768 10152 6786 10170
rect 6768 10170 6786 10188
rect 6768 10188 6786 10206
rect 6786 1656 6804 1674
rect 6786 1674 6804 1692
rect 6786 1692 6804 1710
rect 6786 1710 6804 1728
rect 6786 1728 6804 1746
rect 6786 1746 6804 1764
rect 6786 1764 6804 1782
rect 6786 1782 6804 1800
rect 6786 1800 6804 1818
rect 6786 1818 6804 1836
rect 6786 1836 6804 1854
rect 6786 1854 6804 1872
rect 6786 1872 6804 1890
rect 6786 1890 6804 1908
rect 6786 1908 6804 1926
rect 6786 1926 6804 1944
rect 6786 1944 6804 1962
rect 6786 1962 6804 1980
rect 6786 1980 6804 1998
rect 6786 1998 6804 2016
rect 6786 2016 6804 2034
rect 6786 2034 6804 2052
rect 6786 2052 6804 2070
rect 6786 2070 6804 2088
rect 6786 2088 6804 2106
rect 6786 2106 6804 2124
rect 6786 2124 6804 2142
rect 6786 2142 6804 2160
rect 6786 2160 6804 2178
rect 6786 2178 6804 2196
rect 6786 2196 6804 2214
rect 6786 2214 6804 2232
rect 6786 2232 6804 2250
rect 6786 2250 6804 2268
rect 6786 2268 6804 2286
rect 6786 2286 6804 2304
rect 6786 2304 6804 2322
rect 6786 2322 6804 2340
rect 6786 2340 6804 2358
rect 6786 2358 6804 2376
rect 6786 2376 6804 2394
rect 6786 2394 6804 2412
rect 6786 2412 6804 2430
rect 6786 2430 6804 2448
rect 6786 2448 6804 2466
rect 6786 2466 6804 2484
rect 6786 2484 6804 2502
rect 6786 2502 6804 2520
rect 6786 2520 6804 2538
rect 6786 2538 6804 2556
rect 6786 2556 6804 2574
rect 6786 2574 6804 2592
rect 6786 2592 6804 2610
rect 6786 2610 6804 2628
rect 6786 2628 6804 2646
rect 6786 2646 6804 2664
rect 6786 2664 6804 2682
rect 6786 2682 6804 2700
rect 6786 2700 6804 2718
rect 6786 2718 6804 2736
rect 6786 2736 6804 2754
rect 6786 2754 6804 2772
rect 6786 2772 6804 2790
rect 6786 2790 6804 2808
rect 6786 2808 6804 2826
rect 6786 2826 6804 2844
rect 6786 2844 6804 2862
rect 6786 2862 6804 2880
rect 6786 2880 6804 2898
rect 6786 2898 6804 2916
rect 6786 2916 6804 2934
rect 6786 2934 6804 2952
rect 6786 2952 6804 2970
rect 6786 2970 6804 2988
rect 6786 2988 6804 3006
rect 6786 3006 6804 3024
rect 6786 3186 6804 3204
rect 6786 3204 6804 3222
rect 6786 3222 6804 3240
rect 6786 3240 6804 3258
rect 6786 3258 6804 3276
rect 6786 3276 6804 3294
rect 6786 3294 6804 3312
rect 6786 3312 6804 3330
rect 6786 3330 6804 3348
rect 6786 3348 6804 3366
rect 6786 3366 6804 3384
rect 6786 3384 6804 3402
rect 6786 3402 6804 3420
rect 6786 3420 6804 3438
rect 6786 3438 6804 3456
rect 6786 3456 6804 3474
rect 6786 3474 6804 3492
rect 6786 3492 6804 3510
rect 6786 3510 6804 3528
rect 6786 3528 6804 3546
rect 6786 3546 6804 3564
rect 6786 3564 6804 3582
rect 6786 3762 6804 3780
rect 6786 3780 6804 3798
rect 6786 3798 6804 3816
rect 6786 3816 6804 3834
rect 6786 3834 6804 3852
rect 6786 3852 6804 3870
rect 6786 3870 6804 3888
rect 6786 3888 6804 3906
rect 6786 3906 6804 3924
rect 6786 3924 6804 3942
rect 6786 3942 6804 3960
rect 6786 3960 6804 3978
rect 6786 3978 6804 3996
rect 6786 3996 6804 4014
rect 6786 4014 6804 4032
rect 6786 4032 6804 4050
rect 6786 4050 6804 4068
rect 6786 4068 6804 4086
rect 6786 4086 6804 4104
rect 6786 4104 6804 4122
rect 6786 4122 6804 4140
rect 6786 4140 6804 4158
rect 6786 4158 6804 4176
rect 6786 4176 6804 4194
rect 6786 4194 6804 4212
rect 6786 4212 6804 4230
rect 6786 4230 6804 4248
rect 6786 4248 6804 4266
rect 6786 4266 6804 4284
rect 6786 4284 6804 4302
rect 6786 4302 6804 4320
rect 6786 4320 6804 4338
rect 6786 4338 6804 4356
rect 6786 4356 6804 4374
rect 6786 4374 6804 4392
rect 6786 4392 6804 4410
rect 6786 4410 6804 4428
rect 6786 4428 6804 4446
rect 6786 4446 6804 4464
rect 6786 4464 6804 4482
rect 6786 4482 6804 4500
rect 6786 4500 6804 4518
rect 6786 4518 6804 4536
rect 6786 4536 6804 4554
rect 6786 4554 6804 4572
rect 6786 4572 6804 4590
rect 6786 4590 6804 4608
rect 6786 4608 6804 4626
rect 6786 4626 6804 4644
rect 6786 4644 6804 4662
rect 6786 4662 6804 4680
rect 6786 4680 6804 4698
rect 6786 4698 6804 4716
rect 6786 4716 6804 4734
rect 6786 4734 6804 4752
rect 6786 4752 6804 4770
rect 6786 4770 6804 4788
rect 6786 4788 6804 4806
rect 6786 4806 6804 4824
rect 6786 4824 6804 4842
rect 6786 4842 6804 4860
rect 6786 4860 6804 4878
rect 6786 4878 6804 4896
rect 6786 4896 6804 4914
rect 6786 4914 6804 4932
rect 6786 4932 6804 4950
rect 6786 4950 6804 4968
rect 6786 4968 6804 4986
rect 6786 4986 6804 5004
rect 6786 5004 6804 5022
rect 6786 5022 6804 5040
rect 6786 5040 6804 5058
rect 6786 5058 6804 5076
rect 6786 5076 6804 5094
rect 6786 5094 6804 5112
rect 6786 5112 6804 5130
rect 6786 5130 6804 5148
rect 6786 5148 6804 5166
rect 6786 5166 6804 5184
rect 6786 5184 6804 5202
rect 6786 5202 6804 5220
rect 6786 5220 6804 5238
rect 6786 5238 6804 5256
rect 6786 5256 6804 5274
rect 6786 5274 6804 5292
rect 6786 5292 6804 5310
rect 6786 5310 6804 5328
rect 6786 5328 6804 5346
rect 6786 5346 6804 5364
rect 6786 5364 6804 5382
rect 6786 5382 6804 5400
rect 6786 5400 6804 5418
rect 6786 5418 6804 5436
rect 6786 5436 6804 5454
rect 6786 5454 6804 5472
rect 6786 5472 6804 5490
rect 6786 5490 6804 5508
rect 6786 5508 6804 5526
rect 6786 5526 6804 5544
rect 6786 5544 6804 5562
rect 6786 5562 6804 5580
rect 6786 5580 6804 5598
rect 6786 5598 6804 5616
rect 6786 5616 6804 5634
rect 6786 5634 6804 5652
rect 6786 5652 6804 5670
rect 6786 5670 6804 5688
rect 6786 5688 6804 5706
rect 6786 5706 6804 5724
rect 6786 5724 6804 5742
rect 6786 5742 6804 5760
rect 6786 5760 6804 5778
rect 6786 5778 6804 5796
rect 6786 5796 6804 5814
rect 6786 5814 6804 5832
rect 6786 5832 6804 5850
rect 6786 5850 6804 5868
rect 6786 5868 6804 5886
rect 6786 5886 6804 5904
rect 6786 5904 6804 5922
rect 6786 5922 6804 5940
rect 6786 5940 6804 5958
rect 6786 5958 6804 5976
rect 6786 5976 6804 5994
rect 6786 5994 6804 6012
rect 6786 6012 6804 6030
rect 6786 6030 6804 6048
rect 6786 6048 6804 6066
rect 6786 6066 6804 6084
rect 6786 7290 6804 7308
rect 6786 7308 6804 7326
rect 6786 7326 6804 7344
rect 6786 7344 6804 7362
rect 6786 7362 6804 7380
rect 6786 7380 6804 7398
rect 6786 7398 6804 7416
rect 6786 7416 6804 7434
rect 6786 7434 6804 7452
rect 6786 7452 6804 7470
rect 6786 7470 6804 7488
rect 6786 7488 6804 7506
rect 6786 7506 6804 7524
rect 6786 7524 6804 7542
rect 6786 7542 6804 7560
rect 6786 7560 6804 7578
rect 6786 7578 6804 7596
rect 6786 7596 6804 7614
rect 6786 7614 6804 7632
rect 6786 7632 6804 7650
rect 6786 7650 6804 7668
rect 6786 7668 6804 7686
rect 6786 7686 6804 7704
rect 6786 7704 6804 7722
rect 6786 7722 6804 7740
rect 6786 7740 6804 7758
rect 6786 7758 6804 7776
rect 6786 7776 6804 7794
rect 6786 7794 6804 7812
rect 6786 7812 6804 7830
rect 6786 7830 6804 7848
rect 6786 7848 6804 7866
rect 6786 7866 6804 7884
rect 6786 7884 6804 7902
rect 6786 7902 6804 7920
rect 6786 7920 6804 7938
rect 6786 7938 6804 7956
rect 6786 7956 6804 7974
rect 6786 7974 6804 7992
rect 6786 7992 6804 8010
rect 6786 8010 6804 8028
rect 6786 8028 6804 8046
rect 6786 8046 6804 8064
rect 6786 8064 6804 8082
rect 6786 8082 6804 8100
rect 6786 8100 6804 8118
rect 6786 8118 6804 8136
rect 6786 8136 6804 8154
rect 6786 8154 6804 8172
rect 6786 8172 6804 8190
rect 6786 8190 6804 8208
rect 6786 8208 6804 8226
rect 6786 8226 6804 8244
rect 6786 8244 6804 8262
rect 6786 8262 6804 8280
rect 6786 8280 6804 8298
rect 6786 8298 6804 8316
rect 6786 8316 6804 8334
rect 6786 8334 6804 8352
rect 6786 8352 6804 8370
rect 6786 8370 6804 8388
rect 6786 8388 6804 8406
rect 6786 8406 6804 8424
rect 6786 8424 6804 8442
rect 6786 8442 6804 8460
rect 6786 8460 6804 8478
rect 6786 8478 6804 8496
rect 6786 8496 6804 8514
rect 6786 8514 6804 8532
rect 6786 8532 6804 8550
rect 6786 8550 6804 8568
rect 6786 8568 6804 8586
rect 6786 8586 6804 8604
rect 6786 8604 6804 8622
rect 6786 8622 6804 8640
rect 6786 8640 6804 8658
rect 6786 8658 6804 8676
rect 6786 8676 6804 8694
rect 6786 8694 6804 8712
rect 6786 8712 6804 8730
rect 6786 8730 6804 8748
rect 6786 8748 6804 8766
rect 6786 8766 6804 8784
rect 6786 8784 6804 8802
rect 6786 8802 6804 8820
rect 6786 8820 6804 8838
rect 6786 8838 6804 8856
rect 6786 8856 6804 8874
rect 6786 8874 6804 8892
rect 6786 8892 6804 8910
rect 6786 8910 6804 8928
rect 6786 8928 6804 8946
rect 6786 8946 6804 8964
rect 6786 8964 6804 8982
rect 6786 8982 6804 9000
rect 6786 9000 6804 9018
rect 6786 9018 6804 9036
rect 6786 9036 6804 9054
rect 6786 9054 6804 9072
rect 6786 9072 6804 9090
rect 6786 9090 6804 9108
rect 6786 9108 6804 9126
rect 6786 9126 6804 9144
rect 6786 9144 6804 9162
rect 6786 9162 6804 9180
rect 6786 9180 6804 9198
rect 6786 9198 6804 9216
rect 6786 9216 6804 9234
rect 6786 9234 6804 9252
rect 6786 9252 6804 9270
rect 6786 9270 6804 9288
rect 6786 9288 6804 9306
rect 6786 9306 6804 9324
rect 6786 9324 6804 9342
rect 6786 9342 6804 9360
rect 6786 9360 6804 9378
rect 6786 9378 6804 9396
rect 6786 9396 6804 9414
rect 6786 9414 6804 9432
rect 6786 9432 6804 9450
rect 6786 9450 6804 9468
rect 6786 9468 6804 9486
rect 6786 9486 6804 9504
rect 6786 9504 6804 9522
rect 6786 9522 6804 9540
rect 6786 9540 6804 9558
rect 6786 9558 6804 9576
rect 6786 9576 6804 9594
rect 6786 9594 6804 9612
rect 6786 9612 6804 9630
rect 6786 9630 6804 9648
rect 6786 9648 6804 9666
rect 6786 9666 6804 9684
rect 6786 9684 6804 9702
rect 6786 9702 6804 9720
rect 6786 9720 6804 9738
rect 6786 9738 6804 9756
rect 6786 9756 6804 9774
rect 6786 9774 6804 9792
rect 6786 9792 6804 9810
rect 6786 9810 6804 9828
rect 6786 9828 6804 9846
rect 6786 9846 6804 9864
rect 6786 9864 6804 9882
rect 6786 9882 6804 9900
rect 6786 9900 6804 9918
rect 6786 9918 6804 9936
rect 6786 9936 6804 9954
rect 6786 9954 6804 9972
rect 6786 9972 6804 9990
rect 6786 9990 6804 10008
rect 6786 10008 6804 10026
rect 6786 10026 6804 10044
rect 6786 10044 6804 10062
rect 6786 10062 6804 10080
rect 6786 10080 6804 10098
rect 6786 10098 6804 10116
rect 6786 10116 6804 10134
rect 6786 10134 6804 10152
rect 6786 10152 6804 10170
rect 6786 10170 6804 10188
rect 6786 10188 6804 10206
rect 6786 10206 6804 10224
rect 6804 1674 6822 1692
rect 6804 1692 6822 1710
rect 6804 1710 6822 1728
rect 6804 1728 6822 1746
rect 6804 1746 6822 1764
rect 6804 1764 6822 1782
rect 6804 1782 6822 1800
rect 6804 1800 6822 1818
rect 6804 1818 6822 1836
rect 6804 1836 6822 1854
rect 6804 1854 6822 1872
rect 6804 1872 6822 1890
rect 6804 1890 6822 1908
rect 6804 1908 6822 1926
rect 6804 1926 6822 1944
rect 6804 1944 6822 1962
rect 6804 1962 6822 1980
rect 6804 1980 6822 1998
rect 6804 1998 6822 2016
rect 6804 2016 6822 2034
rect 6804 2034 6822 2052
rect 6804 2052 6822 2070
rect 6804 2070 6822 2088
rect 6804 2088 6822 2106
rect 6804 2106 6822 2124
rect 6804 2124 6822 2142
rect 6804 2142 6822 2160
rect 6804 2160 6822 2178
rect 6804 2178 6822 2196
rect 6804 2196 6822 2214
rect 6804 2214 6822 2232
rect 6804 2232 6822 2250
rect 6804 2250 6822 2268
rect 6804 2268 6822 2286
rect 6804 2286 6822 2304
rect 6804 2304 6822 2322
rect 6804 2322 6822 2340
rect 6804 2340 6822 2358
rect 6804 2358 6822 2376
rect 6804 2376 6822 2394
rect 6804 2394 6822 2412
rect 6804 2412 6822 2430
rect 6804 2430 6822 2448
rect 6804 2448 6822 2466
rect 6804 2466 6822 2484
rect 6804 2484 6822 2502
rect 6804 2502 6822 2520
rect 6804 2520 6822 2538
rect 6804 2538 6822 2556
rect 6804 2556 6822 2574
rect 6804 2574 6822 2592
rect 6804 2592 6822 2610
rect 6804 2610 6822 2628
rect 6804 2628 6822 2646
rect 6804 2646 6822 2664
rect 6804 2664 6822 2682
rect 6804 2682 6822 2700
rect 6804 2700 6822 2718
rect 6804 2718 6822 2736
rect 6804 2736 6822 2754
rect 6804 2754 6822 2772
rect 6804 2772 6822 2790
rect 6804 2790 6822 2808
rect 6804 2808 6822 2826
rect 6804 2826 6822 2844
rect 6804 2844 6822 2862
rect 6804 2862 6822 2880
rect 6804 2880 6822 2898
rect 6804 2898 6822 2916
rect 6804 2916 6822 2934
rect 6804 2934 6822 2952
rect 6804 2952 6822 2970
rect 6804 2970 6822 2988
rect 6804 2988 6822 3006
rect 6804 3006 6822 3024
rect 6804 3024 6822 3042
rect 6804 3204 6822 3222
rect 6804 3222 6822 3240
rect 6804 3240 6822 3258
rect 6804 3258 6822 3276
rect 6804 3276 6822 3294
rect 6804 3294 6822 3312
rect 6804 3312 6822 3330
rect 6804 3330 6822 3348
rect 6804 3348 6822 3366
rect 6804 3366 6822 3384
rect 6804 3384 6822 3402
rect 6804 3402 6822 3420
rect 6804 3420 6822 3438
rect 6804 3438 6822 3456
rect 6804 3456 6822 3474
rect 6804 3474 6822 3492
rect 6804 3492 6822 3510
rect 6804 3510 6822 3528
rect 6804 3528 6822 3546
rect 6804 3546 6822 3564
rect 6804 3564 6822 3582
rect 6804 3582 6822 3600
rect 6804 3780 6822 3798
rect 6804 3798 6822 3816
rect 6804 3816 6822 3834
rect 6804 3834 6822 3852
rect 6804 3852 6822 3870
rect 6804 3870 6822 3888
rect 6804 3888 6822 3906
rect 6804 3906 6822 3924
rect 6804 3924 6822 3942
rect 6804 3942 6822 3960
rect 6804 3960 6822 3978
rect 6804 3978 6822 3996
rect 6804 3996 6822 4014
rect 6804 4014 6822 4032
rect 6804 4032 6822 4050
rect 6804 4050 6822 4068
rect 6804 4068 6822 4086
rect 6804 4086 6822 4104
rect 6804 4104 6822 4122
rect 6804 4122 6822 4140
rect 6804 4140 6822 4158
rect 6804 4158 6822 4176
rect 6804 4176 6822 4194
rect 6804 4194 6822 4212
rect 6804 4212 6822 4230
rect 6804 4230 6822 4248
rect 6804 4248 6822 4266
rect 6804 4266 6822 4284
rect 6804 4284 6822 4302
rect 6804 4302 6822 4320
rect 6804 4320 6822 4338
rect 6804 4338 6822 4356
rect 6804 4356 6822 4374
rect 6804 4374 6822 4392
rect 6804 4392 6822 4410
rect 6804 4410 6822 4428
rect 6804 4428 6822 4446
rect 6804 4446 6822 4464
rect 6804 4464 6822 4482
rect 6804 4482 6822 4500
rect 6804 4500 6822 4518
rect 6804 4518 6822 4536
rect 6804 4536 6822 4554
rect 6804 4554 6822 4572
rect 6804 4572 6822 4590
rect 6804 4590 6822 4608
rect 6804 4608 6822 4626
rect 6804 4626 6822 4644
rect 6804 4644 6822 4662
rect 6804 4662 6822 4680
rect 6804 4680 6822 4698
rect 6804 4698 6822 4716
rect 6804 4716 6822 4734
rect 6804 4734 6822 4752
rect 6804 4752 6822 4770
rect 6804 4770 6822 4788
rect 6804 4788 6822 4806
rect 6804 4806 6822 4824
rect 6804 4824 6822 4842
rect 6804 4842 6822 4860
rect 6804 4860 6822 4878
rect 6804 4878 6822 4896
rect 6804 4896 6822 4914
rect 6804 4914 6822 4932
rect 6804 4932 6822 4950
rect 6804 4950 6822 4968
rect 6804 4968 6822 4986
rect 6804 4986 6822 5004
rect 6804 5004 6822 5022
rect 6804 5022 6822 5040
rect 6804 5040 6822 5058
rect 6804 5058 6822 5076
rect 6804 5076 6822 5094
rect 6804 5094 6822 5112
rect 6804 5112 6822 5130
rect 6804 5130 6822 5148
rect 6804 5148 6822 5166
rect 6804 5166 6822 5184
rect 6804 5184 6822 5202
rect 6804 5202 6822 5220
rect 6804 5220 6822 5238
rect 6804 5238 6822 5256
rect 6804 5256 6822 5274
rect 6804 5274 6822 5292
rect 6804 5292 6822 5310
rect 6804 5310 6822 5328
rect 6804 5328 6822 5346
rect 6804 5346 6822 5364
rect 6804 5364 6822 5382
rect 6804 5382 6822 5400
rect 6804 5400 6822 5418
rect 6804 5418 6822 5436
rect 6804 5436 6822 5454
rect 6804 5454 6822 5472
rect 6804 5472 6822 5490
rect 6804 5490 6822 5508
rect 6804 5508 6822 5526
rect 6804 5526 6822 5544
rect 6804 5544 6822 5562
rect 6804 5562 6822 5580
rect 6804 5580 6822 5598
rect 6804 5598 6822 5616
rect 6804 5616 6822 5634
rect 6804 5634 6822 5652
rect 6804 5652 6822 5670
rect 6804 5670 6822 5688
rect 6804 5688 6822 5706
rect 6804 5706 6822 5724
rect 6804 5724 6822 5742
rect 6804 5742 6822 5760
rect 6804 5760 6822 5778
rect 6804 5778 6822 5796
rect 6804 5796 6822 5814
rect 6804 5814 6822 5832
rect 6804 5832 6822 5850
rect 6804 5850 6822 5868
rect 6804 5868 6822 5886
rect 6804 5886 6822 5904
rect 6804 5904 6822 5922
rect 6804 5922 6822 5940
rect 6804 5940 6822 5958
rect 6804 5958 6822 5976
rect 6804 5976 6822 5994
rect 6804 5994 6822 6012
rect 6804 6012 6822 6030
rect 6804 6030 6822 6048
rect 6804 6048 6822 6066
rect 6804 6066 6822 6084
rect 6804 6084 6822 6102
rect 6804 7344 6822 7362
rect 6804 7362 6822 7380
rect 6804 7380 6822 7398
rect 6804 7398 6822 7416
rect 6804 7416 6822 7434
rect 6804 7434 6822 7452
rect 6804 7452 6822 7470
rect 6804 7470 6822 7488
rect 6804 7488 6822 7506
rect 6804 7506 6822 7524
rect 6804 7524 6822 7542
rect 6804 7542 6822 7560
rect 6804 7560 6822 7578
rect 6804 7578 6822 7596
rect 6804 7596 6822 7614
rect 6804 7614 6822 7632
rect 6804 7632 6822 7650
rect 6804 7650 6822 7668
rect 6804 7668 6822 7686
rect 6804 7686 6822 7704
rect 6804 7704 6822 7722
rect 6804 7722 6822 7740
rect 6804 7740 6822 7758
rect 6804 7758 6822 7776
rect 6804 7776 6822 7794
rect 6804 7794 6822 7812
rect 6804 7812 6822 7830
rect 6804 7830 6822 7848
rect 6804 7848 6822 7866
rect 6804 7866 6822 7884
rect 6804 7884 6822 7902
rect 6804 7902 6822 7920
rect 6804 7920 6822 7938
rect 6804 7938 6822 7956
rect 6804 7956 6822 7974
rect 6804 7974 6822 7992
rect 6804 7992 6822 8010
rect 6804 8010 6822 8028
rect 6804 8028 6822 8046
rect 6804 8046 6822 8064
rect 6804 8064 6822 8082
rect 6804 8082 6822 8100
rect 6804 8100 6822 8118
rect 6804 8118 6822 8136
rect 6804 8136 6822 8154
rect 6804 8154 6822 8172
rect 6804 8172 6822 8190
rect 6804 8190 6822 8208
rect 6804 8208 6822 8226
rect 6804 8226 6822 8244
rect 6804 8244 6822 8262
rect 6804 8262 6822 8280
rect 6804 8280 6822 8298
rect 6804 8298 6822 8316
rect 6804 8316 6822 8334
rect 6804 8334 6822 8352
rect 6804 8352 6822 8370
rect 6804 8370 6822 8388
rect 6804 8388 6822 8406
rect 6804 8406 6822 8424
rect 6804 8424 6822 8442
rect 6804 8442 6822 8460
rect 6804 8460 6822 8478
rect 6804 8478 6822 8496
rect 6804 8496 6822 8514
rect 6804 8514 6822 8532
rect 6804 8532 6822 8550
rect 6804 8550 6822 8568
rect 6804 8568 6822 8586
rect 6804 8586 6822 8604
rect 6804 8604 6822 8622
rect 6804 8622 6822 8640
rect 6804 8640 6822 8658
rect 6804 8658 6822 8676
rect 6804 8676 6822 8694
rect 6804 8694 6822 8712
rect 6804 8712 6822 8730
rect 6804 8730 6822 8748
rect 6804 8748 6822 8766
rect 6804 8766 6822 8784
rect 6804 8784 6822 8802
rect 6804 8802 6822 8820
rect 6804 8820 6822 8838
rect 6804 8838 6822 8856
rect 6804 8856 6822 8874
rect 6804 8874 6822 8892
rect 6804 8892 6822 8910
rect 6804 8910 6822 8928
rect 6804 8928 6822 8946
rect 6804 8946 6822 8964
rect 6804 8964 6822 8982
rect 6804 8982 6822 9000
rect 6804 9000 6822 9018
rect 6804 9018 6822 9036
rect 6804 9036 6822 9054
rect 6804 9054 6822 9072
rect 6804 9072 6822 9090
rect 6804 9090 6822 9108
rect 6804 9108 6822 9126
rect 6804 9126 6822 9144
rect 6804 9144 6822 9162
rect 6804 9162 6822 9180
rect 6804 9180 6822 9198
rect 6804 9198 6822 9216
rect 6804 9216 6822 9234
rect 6804 9234 6822 9252
rect 6804 9252 6822 9270
rect 6804 9270 6822 9288
rect 6804 9288 6822 9306
rect 6804 9306 6822 9324
rect 6804 9324 6822 9342
rect 6804 9342 6822 9360
rect 6804 9360 6822 9378
rect 6804 9378 6822 9396
rect 6804 9396 6822 9414
rect 6804 9414 6822 9432
rect 6804 9432 6822 9450
rect 6804 9450 6822 9468
rect 6804 9468 6822 9486
rect 6804 9486 6822 9504
rect 6804 9504 6822 9522
rect 6804 9522 6822 9540
rect 6804 9540 6822 9558
rect 6804 9558 6822 9576
rect 6804 9576 6822 9594
rect 6804 9594 6822 9612
rect 6804 9612 6822 9630
rect 6804 9630 6822 9648
rect 6804 9648 6822 9666
rect 6804 9666 6822 9684
rect 6804 9684 6822 9702
rect 6804 9702 6822 9720
rect 6804 9720 6822 9738
rect 6804 9738 6822 9756
rect 6804 9756 6822 9774
rect 6804 9774 6822 9792
rect 6804 9792 6822 9810
rect 6804 9810 6822 9828
rect 6804 9828 6822 9846
rect 6804 9846 6822 9864
rect 6804 9864 6822 9882
rect 6804 9882 6822 9900
rect 6804 9900 6822 9918
rect 6804 9918 6822 9936
rect 6804 9936 6822 9954
rect 6804 9954 6822 9972
rect 6804 9972 6822 9990
rect 6804 9990 6822 10008
rect 6804 10008 6822 10026
rect 6804 10026 6822 10044
rect 6804 10044 6822 10062
rect 6804 10062 6822 10080
rect 6804 10080 6822 10098
rect 6804 10098 6822 10116
rect 6804 10116 6822 10134
rect 6804 10134 6822 10152
rect 6804 10152 6822 10170
rect 6804 10170 6822 10188
rect 6804 10188 6822 10206
rect 6804 10206 6822 10224
rect 6804 10224 6822 10242
rect 6822 1674 6840 1692
rect 6822 1692 6840 1710
rect 6822 1710 6840 1728
rect 6822 1728 6840 1746
rect 6822 1746 6840 1764
rect 6822 1764 6840 1782
rect 6822 1782 6840 1800
rect 6822 1800 6840 1818
rect 6822 1818 6840 1836
rect 6822 1836 6840 1854
rect 6822 1854 6840 1872
rect 6822 1872 6840 1890
rect 6822 1890 6840 1908
rect 6822 1908 6840 1926
rect 6822 1926 6840 1944
rect 6822 1944 6840 1962
rect 6822 1962 6840 1980
rect 6822 1980 6840 1998
rect 6822 1998 6840 2016
rect 6822 2016 6840 2034
rect 6822 2034 6840 2052
rect 6822 2052 6840 2070
rect 6822 2070 6840 2088
rect 6822 2088 6840 2106
rect 6822 2106 6840 2124
rect 6822 2124 6840 2142
rect 6822 2142 6840 2160
rect 6822 2160 6840 2178
rect 6822 2178 6840 2196
rect 6822 2196 6840 2214
rect 6822 2214 6840 2232
rect 6822 2232 6840 2250
rect 6822 2250 6840 2268
rect 6822 2268 6840 2286
rect 6822 2286 6840 2304
rect 6822 2304 6840 2322
rect 6822 2322 6840 2340
rect 6822 2340 6840 2358
rect 6822 2358 6840 2376
rect 6822 2376 6840 2394
rect 6822 2394 6840 2412
rect 6822 2412 6840 2430
rect 6822 2430 6840 2448
rect 6822 2448 6840 2466
rect 6822 2466 6840 2484
rect 6822 2484 6840 2502
rect 6822 2502 6840 2520
rect 6822 2520 6840 2538
rect 6822 2538 6840 2556
rect 6822 2556 6840 2574
rect 6822 2574 6840 2592
rect 6822 2592 6840 2610
rect 6822 2610 6840 2628
rect 6822 2628 6840 2646
rect 6822 2646 6840 2664
rect 6822 2664 6840 2682
rect 6822 2682 6840 2700
rect 6822 2700 6840 2718
rect 6822 2718 6840 2736
rect 6822 2736 6840 2754
rect 6822 2754 6840 2772
rect 6822 2772 6840 2790
rect 6822 2790 6840 2808
rect 6822 2808 6840 2826
rect 6822 2826 6840 2844
rect 6822 2844 6840 2862
rect 6822 2862 6840 2880
rect 6822 2880 6840 2898
rect 6822 2898 6840 2916
rect 6822 2916 6840 2934
rect 6822 2934 6840 2952
rect 6822 2952 6840 2970
rect 6822 2970 6840 2988
rect 6822 2988 6840 3006
rect 6822 3006 6840 3024
rect 6822 3024 6840 3042
rect 6822 3204 6840 3222
rect 6822 3222 6840 3240
rect 6822 3240 6840 3258
rect 6822 3258 6840 3276
rect 6822 3276 6840 3294
rect 6822 3294 6840 3312
rect 6822 3312 6840 3330
rect 6822 3330 6840 3348
rect 6822 3348 6840 3366
rect 6822 3366 6840 3384
rect 6822 3384 6840 3402
rect 6822 3402 6840 3420
rect 6822 3420 6840 3438
rect 6822 3438 6840 3456
rect 6822 3456 6840 3474
rect 6822 3474 6840 3492
rect 6822 3492 6840 3510
rect 6822 3510 6840 3528
rect 6822 3528 6840 3546
rect 6822 3546 6840 3564
rect 6822 3564 6840 3582
rect 6822 3582 6840 3600
rect 6822 3600 6840 3618
rect 6822 3816 6840 3834
rect 6822 3834 6840 3852
rect 6822 3852 6840 3870
rect 6822 3870 6840 3888
rect 6822 3888 6840 3906
rect 6822 3906 6840 3924
rect 6822 3924 6840 3942
rect 6822 3942 6840 3960
rect 6822 3960 6840 3978
rect 6822 3978 6840 3996
rect 6822 3996 6840 4014
rect 6822 4014 6840 4032
rect 6822 4032 6840 4050
rect 6822 4050 6840 4068
rect 6822 4068 6840 4086
rect 6822 4086 6840 4104
rect 6822 4104 6840 4122
rect 6822 4122 6840 4140
rect 6822 4140 6840 4158
rect 6822 4158 6840 4176
rect 6822 4176 6840 4194
rect 6822 4194 6840 4212
rect 6822 4212 6840 4230
rect 6822 4230 6840 4248
rect 6822 4248 6840 4266
rect 6822 4266 6840 4284
rect 6822 4284 6840 4302
rect 6822 4302 6840 4320
rect 6822 4320 6840 4338
rect 6822 4338 6840 4356
rect 6822 4356 6840 4374
rect 6822 4374 6840 4392
rect 6822 4392 6840 4410
rect 6822 4410 6840 4428
rect 6822 4428 6840 4446
rect 6822 4446 6840 4464
rect 6822 4464 6840 4482
rect 6822 4482 6840 4500
rect 6822 4500 6840 4518
rect 6822 4518 6840 4536
rect 6822 4536 6840 4554
rect 6822 4554 6840 4572
rect 6822 4572 6840 4590
rect 6822 4590 6840 4608
rect 6822 4608 6840 4626
rect 6822 4626 6840 4644
rect 6822 4644 6840 4662
rect 6822 4662 6840 4680
rect 6822 4680 6840 4698
rect 6822 4698 6840 4716
rect 6822 4716 6840 4734
rect 6822 4734 6840 4752
rect 6822 4752 6840 4770
rect 6822 4770 6840 4788
rect 6822 4788 6840 4806
rect 6822 4806 6840 4824
rect 6822 4824 6840 4842
rect 6822 4842 6840 4860
rect 6822 4860 6840 4878
rect 6822 4878 6840 4896
rect 6822 4896 6840 4914
rect 6822 4914 6840 4932
rect 6822 4932 6840 4950
rect 6822 4950 6840 4968
rect 6822 4968 6840 4986
rect 6822 4986 6840 5004
rect 6822 5004 6840 5022
rect 6822 5022 6840 5040
rect 6822 5040 6840 5058
rect 6822 5058 6840 5076
rect 6822 5076 6840 5094
rect 6822 5094 6840 5112
rect 6822 5112 6840 5130
rect 6822 5130 6840 5148
rect 6822 5148 6840 5166
rect 6822 5166 6840 5184
rect 6822 5184 6840 5202
rect 6822 5202 6840 5220
rect 6822 5220 6840 5238
rect 6822 5238 6840 5256
rect 6822 5256 6840 5274
rect 6822 5274 6840 5292
rect 6822 5292 6840 5310
rect 6822 5310 6840 5328
rect 6822 5328 6840 5346
rect 6822 5346 6840 5364
rect 6822 5364 6840 5382
rect 6822 5382 6840 5400
rect 6822 5400 6840 5418
rect 6822 5418 6840 5436
rect 6822 5436 6840 5454
rect 6822 5454 6840 5472
rect 6822 5472 6840 5490
rect 6822 5490 6840 5508
rect 6822 5508 6840 5526
rect 6822 5526 6840 5544
rect 6822 5544 6840 5562
rect 6822 5562 6840 5580
rect 6822 5580 6840 5598
rect 6822 5598 6840 5616
rect 6822 5616 6840 5634
rect 6822 5634 6840 5652
rect 6822 5652 6840 5670
rect 6822 5670 6840 5688
rect 6822 5688 6840 5706
rect 6822 5706 6840 5724
rect 6822 5724 6840 5742
rect 6822 5742 6840 5760
rect 6822 5760 6840 5778
rect 6822 5778 6840 5796
rect 6822 5796 6840 5814
rect 6822 5814 6840 5832
rect 6822 5832 6840 5850
rect 6822 5850 6840 5868
rect 6822 5868 6840 5886
rect 6822 5886 6840 5904
rect 6822 5904 6840 5922
rect 6822 5922 6840 5940
rect 6822 5940 6840 5958
rect 6822 5958 6840 5976
rect 6822 5976 6840 5994
rect 6822 5994 6840 6012
rect 6822 6012 6840 6030
rect 6822 6030 6840 6048
rect 6822 6048 6840 6066
rect 6822 6066 6840 6084
rect 6822 6084 6840 6102
rect 6822 6102 6840 6120
rect 6822 7380 6840 7398
rect 6822 7398 6840 7416
rect 6822 7416 6840 7434
rect 6822 7434 6840 7452
rect 6822 7452 6840 7470
rect 6822 7470 6840 7488
rect 6822 7488 6840 7506
rect 6822 7506 6840 7524
rect 6822 7524 6840 7542
rect 6822 7542 6840 7560
rect 6822 7560 6840 7578
rect 6822 7578 6840 7596
rect 6822 7596 6840 7614
rect 6822 7614 6840 7632
rect 6822 7632 6840 7650
rect 6822 7650 6840 7668
rect 6822 7668 6840 7686
rect 6822 7686 6840 7704
rect 6822 7704 6840 7722
rect 6822 7722 6840 7740
rect 6822 7740 6840 7758
rect 6822 7758 6840 7776
rect 6822 7776 6840 7794
rect 6822 7794 6840 7812
rect 6822 7812 6840 7830
rect 6822 7830 6840 7848
rect 6822 7848 6840 7866
rect 6822 7866 6840 7884
rect 6822 7884 6840 7902
rect 6822 7902 6840 7920
rect 6822 7920 6840 7938
rect 6822 7938 6840 7956
rect 6822 7956 6840 7974
rect 6822 7974 6840 7992
rect 6822 7992 6840 8010
rect 6822 8010 6840 8028
rect 6822 8028 6840 8046
rect 6822 8046 6840 8064
rect 6822 8064 6840 8082
rect 6822 8082 6840 8100
rect 6822 8100 6840 8118
rect 6822 8118 6840 8136
rect 6822 8136 6840 8154
rect 6822 8154 6840 8172
rect 6822 8172 6840 8190
rect 6822 8190 6840 8208
rect 6822 8208 6840 8226
rect 6822 8226 6840 8244
rect 6822 8244 6840 8262
rect 6822 8262 6840 8280
rect 6822 8280 6840 8298
rect 6822 8298 6840 8316
rect 6822 8316 6840 8334
rect 6822 8334 6840 8352
rect 6822 8352 6840 8370
rect 6822 8370 6840 8388
rect 6822 8388 6840 8406
rect 6822 8406 6840 8424
rect 6822 8424 6840 8442
rect 6822 8442 6840 8460
rect 6822 8460 6840 8478
rect 6822 8478 6840 8496
rect 6822 8496 6840 8514
rect 6822 8514 6840 8532
rect 6822 8532 6840 8550
rect 6822 8550 6840 8568
rect 6822 8568 6840 8586
rect 6822 8586 6840 8604
rect 6822 8604 6840 8622
rect 6822 8622 6840 8640
rect 6822 8640 6840 8658
rect 6822 8658 6840 8676
rect 6822 8676 6840 8694
rect 6822 8694 6840 8712
rect 6822 8712 6840 8730
rect 6822 8730 6840 8748
rect 6822 8748 6840 8766
rect 6822 8766 6840 8784
rect 6822 8784 6840 8802
rect 6822 8802 6840 8820
rect 6822 8820 6840 8838
rect 6822 8838 6840 8856
rect 6822 8856 6840 8874
rect 6822 8874 6840 8892
rect 6822 8892 6840 8910
rect 6822 8910 6840 8928
rect 6822 8928 6840 8946
rect 6822 8946 6840 8964
rect 6822 8964 6840 8982
rect 6822 8982 6840 9000
rect 6822 9000 6840 9018
rect 6822 9018 6840 9036
rect 6822 9036 6840 9054
rect 6822 9054 6840 9072
rect 6822 9072 6840 9090
rect 6822 9090 6840 9108
rect 6822 9108 6840 9126
rect 6822 9126 6840 9144
rect 6822 9144 6840 9162
rect 6822 9162 6840 9180
rect 6822 9180 6840 9198
rect 6822 9198 6840 9216
rect 6822 9216 6840 9234
rect 6822 9234 6840 9252
rect 6822 9252 6840 9270
rect 6822 9270 6840 9288
rect 6822 9288 6840 9306
rect 6822 9306 6840 9324
rect 6822 9324 6840 9342
rect 6822 9342 6840 9360
rect 6822 9360 6840 9378
rect 6822 9378 6840 9396
rect 6822 9396 6840 9414
rect 6822 9414 6840 9432
rect 6822 9432 6840 9450
rect 6822 9450 6840 9468
rect 6822 9468 6840 9486
rect 6822 9486 6840 9504
rect 6822 9504 6840 9522
rect 6822 9522 6840 9540
rect 6822 9540 6840 9558
rect 6822 9558 6840 9576
rect 6822 9576 6840 9594
rect 6822 9594 6840 9612
rect 6822 9612 6840 9630
rect 6822 9630 6840 9648
rect 6822 9648 6840 9666
rect 6822 9666 6840 9684
rect 6822 9684 6840 9702
rect 6822 9702 6840 9720
rect 6822 9720 6840 9738
rect 6822 9738 6840 9756
rect 6822 9756 6840 9774
rect 6822 9774 6840 9792
rect 6822 9792 6840 9810
rect 6822 9810 6840 9828
rect 6822 9828 6840 9846
rect 6822 9846 6840 9864
rect 6822 9864 6840 9882
rect 6822 9882 6840 9900
rect 6822 9900 6840 9918
rect 6822 9918 6840 9936
rect 6822 9936 6840 9954
rect 6822 9954 6840 9972
rect 6822 9972 6840 9990
rect 6822 9990 6840 10008
rect 6822 10008 6840 10026
rect 6822 10026 6840 10044
rect 6822 10044 6840 10062
rect 6822 10062 6840 10080
rect 6822 10080 6840 10098
rect 6822 10098 6840 10116
rect 6822 10116 6840 10134
rect 6822 10134 6840 10152
rect 6822 10152 6840 10170
rect 6822 10170 6840 10188
rect 6822 10188 6840 10206
rect 6822 10206 6840 10224
rect 6822 10224 6840 10242
rect 6822 10242 6840 10260
rect 6840 1692 6858 1710
rect 6840 1710 6858 1728
rect 6840 1728 6858 1746
rect 6840 1746 6858 1764
rect 6840 1764 6858 1782
rect 6840 1782 6858 1800
rect 6840 1800 6858 1818
rect 6840 1818 6858 1836
rect 6840 1836 6858 1854
rect 6840 1854 6858 1872
rect 6840 1872 6858 1890
rect 6840 1890 6858 1908
rect 6840 1908 6858 1926
rect 6840 1926 6858 1944
rect 6840 1944 6858 1962
rect 6840 1962 6858 1980
rect 6840 1980 6858 1998
rect 6840 1998 6858 2016
rect 6840 2016 6858 2034
rect 6840 2034 6858 2052
rect 6840 2052 6858 2070
rect 6840 2070 6858 2088
rect 6840 2088 6858 2106
rect 6840 2106 6858 2124
rect 6840 2124 6858 2142
rect 6840 2142 6858 2160
rect 6840 2160 6858 2178
rect 6840 2178 6858 2196
rect 6840 2196 6858 2214
rect 6840 2214 6858 2232
rect 6840 2232 6858 2250
rect 6840 2250 6858 2268
rect 6840 2268 6858 2286
rect 6840 2286 6858 2304
rect 6840 2304 6858 2322
rect 6840 2322 6858 2340
rect 6840 2340 6858 2358
rect 6840 2358 6858 2376
rect 6840 2376 6858 2394
rect 6840 2394 6858 2412
rect 6840 2412 6858 2430
rect 6840 2430 6858 2448
rect 6840 2448 6858 2466
rect 6840 2466 6858 2484
rect 6840 2484 6858 2502
rect 6840 2502 6858 2520
rect 6840 2520 6858 2538
rect 6840 2538 6858 2556
rect 6840 2556 6858 2574
rect 6840 2574 6858 2592
rect 6840 2592 6858 2610
rect 6840 2610 6858 2628
rect 6840 2628 6858 2646
rect 6840 2646 6858 2664
rect 6840 2664 6858 2682
rect 6840 2682 6858 2700
rect 6840 2700 6858 2718
rect 6840 2718 6858 2736
rect 6840 2736 6858 2754
rect 6840 2754 6858 2772
rect 6840 2772 6858 2790
rect 6840 2790 6858 2808
rect 6840 2808 6858 2826
rect 6840 2826 6858 2844
rect 6840 2844 6858 2862
rect 6840 2862 6858 2880
rect 6840 2880 6858 2898
rect 6840 2898 6858 2916
rect 6840 2916 6858 2934
rect 6840 2934 6858 2952
rect 6840 2952 6858 2970
rect 6840 2970 6858 2988
rect 6840 2988 6858 3006
rect 6840 3006 6858 3024
rect 6840 3024 6858 3042
rect 6840 3222 6858 3240
rect 6840 3240 6858 3258
rect 6840 3258 6858 3276
rect 6840 3276 6858 3294
rect 6840 3294 6858 3312
rect 6840 3312 6858 3330
rect 6840 3330 6858 3348
rect 6840 3348 6858 3366
rect 6840 3366 6858 3384
rect 6840 3384 6858 3402
rect 6840 3402 6858 3420
rect 6840 3420 6858 3438
rect 6840 3438 6858 3456
rect 6840 3456 6858 3474
rect 6840 3474 6858 3492
rect 6840 3492 6858 3510
rect 6840 3510 6858 3528
rect 6840 3528 6858 3546
rect 6840 3546 6858 3564
rect 6840 3564 6858 3582
rect 6840 3582 6858 3600
rect 6840 3600 6858 3618
rect 6840 3618 6858 3636
rect 6840 3834 6858 3852
rect 6840 3852 6858 3870
rect 6840 3870 6858 3888
rect 6840 3888 6858 3906
rect 6840 3906 6858 3924
rect 6840 3924 6858 3942
rect 6840 3942 6858 3960
rect 6840 3960 6858 3978
rect 6840 3978 6858 3996
rect 6840 3996 6858 4014
rect 6840 4014 6858 4032
rect 6840 4032 6858 4050
rect 6840 4050 6858 4068
rect 6840 4068 6858 4086
rect 6840 4086 6858 4104
rect 6840 4104 6858 4122
rect 6840 4122 6858 4140
rect 6840 4140 6858 4158
rect 6840 4158 6858 4176
rect 6840 4176 6858 4194
rect 6840 4194 6858 4212
rect 6840 4212 6858 4230
rect 6840 4230 6858 4248
rect 6840 4248 6858 4266
rect 6840 4266 6858 4284
rect 6840 4284 6858 4302
rect 6840 4302 6858 4320
rect 6840 4320 6858 4338
rect 6840 4338 6858 4356
rect 6840 4356 6858 4374
rect 6840 4374 6858 4392
rect 6840 4392 6858 4410
rect 6840 4410 6858 4428
rect 6840 4428 6858 4446
rect 6840 4446 6858 4464
rect 6840 4464 6858 4482
rect 6840 4482 6858 4500
rect 6840 4500 6858 4518
rect 6840 4518 6858 4536
rect 6840 4536 6858 4554
rect 6840 4554 6858 4572
rect 6840 4572 6858 4590
rect 6840 4590 6858 4608
rect 6840 4608 6858 4626
rect 6840 4626 6858 4644
rect 6840 4644 6858 4662
rect 6840 4662 6858 4680
rect 6840 4680 6858 4698
rect 6840 4698 6858 4716
rect 6840 4716 6858 4734
rect 6840 4734 6858 4752
rect 6840 4752 6858 4770
rect 6840 4770 6858 4788
rect 6840 4788 6858 4806
rect 6840 4806 6858 4824
rect 6840 4824 6858 4842
rect 6840 4842 6858 4860
rect 6840 4860 6858 4878
rect 6840 4878 6858 4896
rect 6840 4896 6858 4914
rect 6840 4914 6858 4932
rect 6840 4932 6858 4950
rect 6840 4950 6858 4968
rect 6840 4968 6858 4986
rect 6840 4986 6858 5004
rect 6840 5004 6858 5022
rect 6840 5022 6858 5040
rect 6840 5040 6858 5058
rect 6840 5058 6858 5076
rect 6840 5076 6858 5094
rect 6840 5094 6858 5112
rect 6840 5112 6858 5130
rect 6840 5130 6858 5148
rect 6840 5148 6858 5166
rect 6840 5166 6858 5184
rect 6840 5184 6858 5202
rect 6840 5202 6858 5220
rect 6840 5220 6858 5238
rect 6840 5238 6858 5256
rect 6840 5256 6858 5274
rect 6840 5274 6858 5292
rect 6840 5292 6858 5310
rect 6840 5310 6858 5328
rect 6840 5328 6858 5346
rect 6840 5346 6858 5364
rect 6840 5364 6858 5382
rect 6840 5382 6858 5400
rect 6840 5400 6858 5418
rect 6840 5418 6858 5436
rect 6840 5436 6858 5454
rect 6840 5454 6858 5472
rect 6840 5472 6858 5490
rect 6840 5490 6858 5508
rect 6840 5508 6858 5526
rect 6840 5526 6858 5544
rect 6840 5544 6858 5562
rect 6840 5562 6858 5580
rect 6840 5580 6858 5598
rect 6840 5598 6858 5616
rect 6840 5616 6858 5634
rect 6840 5634 6858 5652
rect 6840 5652 6858 5670
rect 6840 5670 6858 5688
rect 6840 5688 6858 5706
rect 6840 5706 6858 5724
rect 6840 5724 6858 5742
rect 6840 5742 6858 5760
rect 6840 5760 6858 5778
rect 6840 5778 6858 5796
rect 6840 5796 6858 5814
rect 6840 5814 6858 5832
rect 6840 5832 6858 5850
rect 6840 5850 6858 5868
rect 6840 5868 6858 5886
rect 6840 5886 6858 5904
rect 6840 5904 6858 5922
rect 6840 5922 6858 5940
rect 6840 5940 6858 5958
rect 6840 5958 6858 5976
rect 6840 5976 6858 5994
rect 6840 5994 6858 6012
rect 6840 6012 6858 6030
rect 6840 6030 6858 6048
rect 6840 6048 6858 6066
rect 6840 6066 6858 6084
rect 6840 6084 6858 6102
rect 6840 6102 6858 6120
rect 6840 6120 6858 6138
rect 6840 7434 6858 7452
rect 6840 7452 6858 7470
rect 6840 7470 6858 7488
rect 6840 7488 6858 7506
rect 6840 7506 6858 7524
rect 6840 7524 6858 7542
rect 6840 7542 6858 7560
rect 6840 7560 6858 7578
rect 6840 7578 6858 7596
rect 6840 7596 6858 7614
rect 6840 7614 6858 7632
rect 6840 7632 6858 7650
rect 6840 7650 6858 7668
rect 6840 7668 6858 7686
rect 6840 7686 6858 7704
rect 6840 7704 6858 7722
rect 6840 7722 6858 7740
rect 6840 7740 6858 7758
rect 6840 7758 6858 7776
rect 6840 7776 6858 7794
rect 6840 7794 6858 7812
rect 6840 7812 6858 7830
rect 6840 7830 6858 7848
rect 6840 7848 6858 7866
rect 6840 7866 6858 7884
rect 6840 7884 6858 7902
rect 6840 7902 6858 7920
rect 6840 7920 6858 7938
rect 6840 7938 6858 7956
rect 6840 7956 6858 7974
rect 6840 7974 6858 7992
rect 6840 7992 6858 8010
rect 6840 8010 6858 8028
rect 6840 8028 6858 8046
rect 6840 8046 6858 8064
rect 6840 8064 6858 8082
rect 6840 8082 6858 8100
rect 6840 8100 6858 8118
rect 6840 8118 6858 8136
rect 6840 8136 6858 8154
rect 6840 8154 6858 8172
rect 6840 8172 6858 8190
rect 6840 8190 6858 8208
rect 6840 8208 6858 8226
rect 6840 8226 6858 8244
rect 6840 8244 6858 8262
rect 6840 8262 6858 8280
rect 6840 8280 6858 8298
rect 6840 8298 6858 8316
rect 6840 8316 6858 8334
rect 6840 8334 6858 8352
rect 6840 8352 6858 8370
rect 6840 8370 6858 8388
rect 6840 8388 6858 8406
rect 6840 8406 6858 8424
rect 6840 8424 6858 8442
rect 6840 8442 6858 8460
rect 6840 8460 6858 8478
rect 6840 8478 6858 8496
rect 6840 8496 6858 8514
rect 6840 8514 6858 8532
rect 6840 8532 6858 8550
rect 6840 8550 6858 8568
rect 6840 8568 6858 8586
rect 6840 8586 6858 8604
rect 6840 8604 6858 8622
rect 6840 8622 6858 8640
rect 6840 8640 6858 8658
rect 6840 8658 6858 8676
rect 6840 8676 6858 8694
rect 6840 8694 6858 8712
rect 6840 8712 6858 8730
rect 6840 8730 6858 8748
rect 6840 8748 6858 8766
rect 6840 8766 6858 8784
rect 6840 8784 6858 8802
rect 6840 8802 6858 8820
rect 6840 8820 6858 8838
rect 6840 8838 6858 8856
rect 6840 8856 6858 8874
rect 6840 8874 6858 8892
rect 6840 8892 6858 8910
rect 6840 8910 6858 8928
rect 6840 8928 6858 8946
rect 6840 8946 6858 8964
rect 6840 8964 6858 8982
rect 6840 8982 6858 9000
rect 6840 9000 6858 9018
rect 6840 9018 6858 9036
rect 6840 9036 6858 9054
rect 6840 9054 6858 9072
rect 6840 9072 6858 9090
rect 6840 9090 6858 9108
rect 6840 9108 6858 9126
rect 6840 9126 6858 9144
rect 6840 9144 6858 9162
rect 6840 9162 6858 9180
rect 6840 9180 6858 9198
rect 6840 9198 6858 9216
rect 6840 9216 6858 9234
rect 6840 9234 6858 9252
rect 6840 9252 6858 9270
rect 6840 9270 6858 9288
rect 6840 9288 6858 9306
rect 6840 9306 6858 9324
rect 6840 9324 6858 9342
rect 6840 9342 6858 9360
rect 6840 9360 6858 9378
rect 6840 9378 6858 9396
rect 6840 9396 6858 9414
rect 6840 9414 6858 9432
rect 6840 9432 6858 9450
rect 6840 9450 6858 9468
rect 6840 9468 6858 9486
rect 6840 9486 6858 9504
rect 6840 9504 6858 9522
rect 6840 9522 6858 9540
rect 6840 9540 6858 9558
rect 6840 9558 6858 9576
rect 6840 9576 6858 9594
rect 6840 9594 6858 9612
rect 6840 9612 6858 9630
rect 6840 9630 6858 9648
rect 6840 9648 6858 9666
rect 6840 9666 6858 9684
rect 6840 9684 6858 9702
rect 6840 9702 6858 9720
rect 6840 9720 6858 9738
rect 6840 9738 6858 9756
rect 6840 9756 6858 9774
rect 6840 9774 6858 9792
rect 6840 9792 6858 9810
rect 6840 9810 6858 9828
rect 6840 9828 6858 9846
rect 6840 9846 6858 9864
rect 6840 9864 6858 9882
rect 6840 9882 6858 9900
rect 6840 9900 6858 9918
rect 6840 9918 6858 9936
rect 6840 9936 6858 9954
rect 6840 9954 6858 9972
rect 6840 9972 6858 9990
rect 6840 9990 6858 10008
rect 6840 10008 6858 10026
rect 6840 10026 6858 10044
rect 6840 10044 6858 10062
rect 6840 10062 6858 10080
rect 6840 10080 6858 10098
rect 6840 10098 6858 10116
rect 6840 10116 6858 10134
rect 6840 10134 6858 10152
rect 6840 10152 6858 10170
rect 6840 10170 6858 10188
rect 6840 10188 6858 10206
rect 6840 10206 6858 10224
rect 6840 10224 6858 10242
rect 6840 10242 6858 10260
rect 6840 10260 6858 10278
rect 6858 1710 6876 1728
rect 6858 1728 6876 1746
rect 6858 1746 6876 1764
rect 6858 1764 6876 1782
rect 6858 1782 6876 1800
rect 6858 1800 6876 1818
rect 6858 1818 6876 1836
rect 6858 1836 6876 1854
rect 6858 1854 6876 1872
rect 6858 1872 6876 1890
rect 6858 1890 6876 1908
rect 6858 1908 6876 1926
rect 6858 1926 6876 1944
rect 6858 1944 6876 1962
rect 6858 1962 6876 1980
rect 6858 1980 6876 1998
rect 6858 1998 6876 2016
rect 6858 2016 6876 2034
rect 6858 2034 6876 2052
rect 6858 2052 6876 2070
rect 6858 2070 6876 2088
rect 6858 2088 6876 2106
rect 6858 2106 6876 2124
rect 6858 2124 6876 2142
rect 6858 2142 6876 2160
rect 6858 2160 6876 2178
rect 6858 2178 6876 2196
rect 6858 2196 6876 2214
rect 6858 2214 6876 2232
rect 6858 2232 6876 2250
rect 6858 2250 6876 2268
rect 6858 2268 6876 2286
rect 6858 2286 6876 2304
rect 6858 2304 6876 2322
rect 6858 2322 6876 2340
rect 6858 2340 6876 2358
rect 6858 2358 6876 2376
rect 6858 2376 6876 2394
rect 6858 2394 6876 2412
rect 6858 2412 6876 2430
rect 6858 2430 6876 2448
rect 6858 2448 6876 2466
rect 6858 2466 6876 2484
rect 6858 2484 6876 2502
rect 6858 2502 6876 2520
rect 6858 2520 6876 2538
rect 6858 2538 6876 2556
rect 6858 2556 6876 2574
rect 6858 2574 6876 2592
rect 6858 2592 6876 2610
rect 6858 2610 6876 2628
rect 6858 2628 6876 2646
rect 6858 2646 6876 2664
rect 6858 2664 6876 2682
rect 6858 2682 6876 2700
rect 6858 2700 6876 2718
rect 6858 2718 6876 2736
rect 6858 2736 6876 2754
rect 6858 2754 6876 2772
rect 6858 2772 6876 2790
rect 6858 2790 6876 2808
rect 6858 2808 6876 2826
rect 6858 2826 6876 2844
rect 6858 2844 6876 2862
rect 6858 2862 6876 2880
rect 6858 2880 6876 2898
rect 6858 2898 6876 2916
rect 6858 2916 6876 2934
rect 6858 2934 6876 2952
rect 6858 2952 6876 2970
rect 6858 2970 6876 2988
rect 6858 2988 6876 3006
rect 6858 3006 6876 3024
rect 6858 3024 6876 3042
rect 6858 3042 6876 3060
rect 6858 3222 6876 3240
rect 6858 3240 6876 3258
rect 6858 3258 6876 3276
rect 6858 3276 6876 3294
rect 6858 3294 6876 3312
rect 6858 3312 6876 3330
rect 6858 3330 6876 3348
rect 6858 3348 6876 3366
rect 6858 3366 6876 3384
rect 6858 3384 6876 3402
rect 6858 3402 6876 3420
rect 6858 3420 6876 3438
rect 6858 3438 6876 3456
rect 6858 3456 6876 3474
rect 6858 3474 6876 3492
rect 6858 3492 6876 3510
rect 6858 3510 6876 3528
rect 6858 3528 6876 3546
rect 6858 3546 6876 3564
rect 6858 3564 6876 3582
rect 6858 3582 6876 3600
rect 6858 3600 6876 3618
rect 6858 3618 6876 3636
rect 6858 3636 6876 3654
rect 6858 3852 6876 3870
rect 6858 3870 6876 3888
rect 6858 3888 6876 3906
rect 6858 3906 6876 3924
rect 6858 3924 6876 3942
rect 6858 3942 6876 3960
rect 6858 3960 6876 3978
rect 6858 3978 6876 3996
rect 6858 3996 6876 4014
rect 6858 4014 6876 4032
rect 6858 4032 6876 4050
rect 6858 4050 6876 4068
rect 6858 4068 6876 4086
rect 6858 4086 6876 4104
rect 6858 4104 6876 4122
rect 6858 4122 6876 4140
rect 6858 4140 6876 4158
rect 6858 4158 6876 4176
rect 6858 4176 6876 4194
rect 6858 4194 6876 4212
rect 6858 4212 6876 4230
rect 6858 4230 6876 4248
rect 6858 4248 6876 4266
rect 6858 4266 6876 4284
rect 6858 4284 6876 4302
rect 6858 4302 6876 4320
rect 6858 4320 6876 4338
rect 6858 4338 6876 4356
rect 6858 4356 6876 4374
rect 6858 4374 6876 4392
rect 6858 4392 6876 4410
rect 6858 4410 6876 4428
rect 6858 4428 6876 4446
rect 6858 4446 6876 4464
rect 6858 4464 6876 4482
rect 6858 4482 6876 4500
rect 6858 4500 6876 4518
rect 6858 4518 6876 4536
rect 6858 4536 6876 4554
rect 6858 4554 6876 4572
rect 6858 4572 6876 4590
rect 6858 4590 6876 4608
rect 6858 4608 6876 4626
rect 6858 4626 6876 4644
rect 6858 4644 6876 4662
rect 6858 4662 6876 4680
rect 6858 4680 6876 4698
rect 6858 4698 6876 4716
rect 6858 4716 6876 4734
rect 6858 4734 6876 4752
rect 6858 4752 6876 4770
rect 6858 4770 6876 4788
rect 6858 4788 6876 4806
rect 6858 4806 6876 4824
rect 6858 4824 6876 4842
rect 6858 4842 6876 4860
rect 6858 4860 6876 4878
rect 6858 4878 6876 4896
rect 6858 4896 6876 4914
rect 6858 4914 6876 4932
rect 6858 4932 6876 4950
rect 6858 4950 6876 4968
rect 6858 4968 6876 4986
rect 6858 4986 6876 5004
rect 6858 5004 6876 5022
rect 6858 5022 6876 5040
rect 6858 5040 6876 5058
rect 6858 5058 6876 5076
rect 6858 5076 6876 5094
rect 6858 5094 6876 5112
rect 6858 5112 6876 5130
rect 6858 5130 6876 5148
rect 6858 5148 6876 5166
rect 6858 5166 6876 5184
rect 6858 5184 6876 5202
rect 6858 5202 6876 5220
rect 6858 5220 6876 5238
rect 6858 5238 6876 5256
rect 6858 5256 6876 5274
rect 6858 5274 6876 5292
rect 6858 5292 6876 5310
rect 6858 5310 6876 5328
rect 6858 5328 6876 5346
rect 6858 5346 6876 5364
rect 6858 5364 6876 5382
rect 6858 5382 6876 5400
rect 6858 5400 6876 5418
rect 6858 5418 6876 5436
rect 6858 5436 6876 5454
rect 6858 5454 6876 5472
rect 6858 5472 6876 5490
rect 6858 5490 6876 5508
rect 6858 5508 6876 5526
rect 6858 5526 6876 5544
rect 6858 5544 6876 5562
rect 6858 5562 6876 5580
rect 6858 5580 6876 5598
rect 6858 5598 6876 5616
rect 6858 5616 6876 5634
rect 6858 5634 6876 5652
rect 6858 5652 6876 5670
rect 6858 5670 6876 5688
rect 6858 5688 6876 5706
rect 6858 5706 6876 5724
rect 6858 5724 6876 5742
rect 6858 5742 6876 5760
rect 6858 5760 6876 5778
rect 6858 5778 6876 5796
rect 6858 5796 6876 5814
rect 6858 5814 6876 5832
rect 6858 5832 6876 5850
rect 6858 5850 6876 5868
rect 6858 5868 6876 5886
rect 6858 5886 6876 5904
rect 6858 5904 6876 5922
rect 6858 5922 6876 5940
rect 6858 5940 6876 5958
rect 6858 5958 6876 5976
rect 6858 5976 6876 5994
rect 6858 5994 6876 6012
rect 6858 6012 6876 6030
rect 6858 6030 6876 6048
rect 6858 6048 6876 6066
rect 6858 6066 6876 6084
rect 6858 6084 6876 6102
rect 6858 6102 6876 6120
rect 6858 6120 6876 6138
rect 6858 7488 6876 7506
rect 6858 7506 6876 7524
rect 6858 7524 6876 7542
rect 6858 7542 6876 7560
rect 6858 7560 6876 7578
rect 6858 7578 6876 7596
rect 6858 7596 6876 7614
rect 6858 7614 6876 7632
rect 6858 7632 6876 7650
rect 6858 7650 6876 7668
rect 6858 7668 6876 7686
rect 6858 7686 6876 7704
rect 6858 7704 6876 7722
rect 6858 7722 6876 7740
rect 6858 7740 6876 7758
rect 6858 7758 6876 7776
rect 6858 7776 6876 7794
rect 6858 7794 6876 7812
rect 6858 7812 6876 7830
rect 6858 7830 6876 7848
rect 6858 7848 6876 7866
rect 6858 7866 6876 7884
rect 6858 7884 6876 7902
rect 6858 7902 6876 7920
rect 6858 7920 6876 7938
rect 6858 7938 6876 7956
rect 6858 7956 6876 7974
rect 6858 7974 6876 7992
rect 6858 7992 6876 8010
rect 6858 8010 6876 8028
rect 6858 8028 6876 8046
rect 6858 8046 6876 8064
rect 6858 8064 6876 8082
rect 6858 8082 6876 8100
rect 6858 8100 6876 8118
rect 6858 8118 6876 8136
rect 6858 8136 6876 8154
rect 6858 8154 6876 8172
rect 6858 8172 6876 8190
rect 6858 8190 6876 8208
rect 6858 8208 6876 8226
rect 6858 8226 6876 8244
rect 6858 8244 6876 8262
rect 6858 8262 6876 8280
rect 6858 8280 6876 8298
rect 6858 8298 6876 8316
rect 6858 8316 6876 8334
rect 6858 8334 6876 8352
rect 6858 8352 6876 8370
rect 6858 8370 6876 8388
rect 6858 8388 6876 8406
rect 6858 8406 6876 8424
rect 6858 8424 6876 8442
rect 6858 8442 6876 8460
rect 6858 8460 6876 8478
rect 6858 8478 6876 8496
rect 6858 8496 6876 8514
rect 6858 8514 6876 8532
rect 6858 8532 6876 8550
rect 6858 8550 6876 8568
rect 6858 8568 6876 8586
rect 6858 8586 6876 8604
rect 6858 8604 6876 8622
rect 6858 8622 6876 8640
rect 6858 8640 6876 8658
rect 6858 8658 6876 8676
rect 6858 8676 6876 8694
rect 6858 8694 6876 8712
rect 6858 8712 6876 8730
rect 6858 8730 6876 8748
rect 6858 8748 6876 8766
rect 6858 8766 6876 8784
rect 6858 8784 6876 8802
rect 6858 8802 6876 8820
rect 6858 8820 6876 8838
rect 6858 8838 6876 8856
rect 6858 8856 6876 8874
rect 6858 8874 6876 8892
rect 6858 8892 6876 8910
rect 6858 8910 6876 8928
rect 6858 8928 6876 8946
rect 6858 8946 6876 8964
rect 6858 8964 6876 8982
rect 6858 8982 6876 9000
rect 6858 9000 6876 9018
rect 6858 9018 6876 9036
rect 6858 9036 6876 9054
rect 6858 9054 6876 9072
rect 6858 9072 6876 9090
rect 6858 9090 6876 9108
rect 6858 9108 6876 9126
rect 6858 9126 6876 9144
rect 6858 9144 6876 9162
rect 6858 9162 6876 9180
rect 6858 9180 6876 9198
rect 6858 9198 6876 9216
rect 6858 9216 6876 9234
rect 6858 9234 6876 9252
rect 6858 9252 6876 9270
rect 6858 9270 6876 9288
rect 6858 9288 6876 9306
rect 6858 9306 6876 9324
rect 6858 9324 6876 9342
rect 6858 9342 6876 9360
rect 6858 9360 6876 9378
rect 6858 9378 6876 9396
rect 6858 9396 6876 9414
rect 6858 9414 6876 9432
rect 6858 9432 6876 9450
rect 6858 9450 6876 9468
rect 6858 9468 6876 9486
rect 6858 9486 6876 9504
rect 6858 9504 6876 9522
rect 6858 9522 6876 9540
rect 6858 9540 6876 9558
rect 6858 9558 6876 9576
rect 6858 9576 6876 9594
rect 6858 9594 6876 9612
rect 6858 9612 6876 9630
rect 6858 9630 6876 9648
rect 6858 9648 6876 9666
rect 6858 9666 6876 9684
rect 6858 9684 6876 9702
rect 6858 9702 6876 9720
rect 6858 9720 6876 9738
rect 6858 9738 6876 9756
rect 6858 9756 6876 9774
rect 6858 9774 6876 9792
rect 6858 9792 6876 9810
rect 6858 9810 6876 9828
rect 6858 9828 6876 9846
rect 6858 9846 6876 9864
rect 6858 9864 6876 9882
rect 6858 9882 6876 9900
rect 6858 9900 6876 9918
rect 6858 9918 6876 9936
rect 6858 9936 6876 9954
rect 6858 9954 6876 9972
rect 6858 9972 6876 9990
rect 6858 9990 6876 10008
rect 6858 10008 6876 10026
rect 6858 10026 6876 10044
rect 6858 10044 6876 10062
rect 6858 10062 6876 10080
rect 6858 10080 6876 10098
rect 6858 10098 6876 10116
rect 6858 10116 6876 10134
rect 6858 10134 6876 10152
rect 6858 10152 6876 10170
rect 6858 10170 6876 10188
rect 6858 10188 6876 10206
rect 6858 10206 6876 10224
rect 6858 10224 6876 10242
rect 6858 10242 6876 10260
rect 6858 10260 6876 10278
rect 6858 10278 6876 10296
rect 6858 10296 6876 10314
rect 6876 1710 6894 1728
rect 6876 1728 6894 1746
rect 6876 1746 6894 1764
rect 6876 1764 6894 1782
rect 6876 1782 6894 1800
rect 6876 1800 6894 1818
rect 6876 1818 6894 1836
rect 6876 1836 6894 1854
rect 6876 1854 6894 1872
rect 6876 1872 6894 1890
rect 6876 1890 6894 1908
rect 6876 1908 6894 1926
rect 6876 1926 6894 1944
rect 6876 1944 6894 1962
rect 6876 1962 6894 1980
rect 6876 1980 6894 1998
rect 6876 1998 6894 2016
rect 6876 2016 6894 2034
rect 6876 2034 6894 2052
rect 6876 2052 6894 2070
rect 6876 2070 6894 2088
rect 6876 2088 6894 2106
rect 6876 2106 6894 2124
rect 6876 2124 6894 2142
rect 6876 2142 6894 2160
rect 6876 2160 6894 2178
rect 6876 2178 6894 2196
rect 6876 2196 6894 2214
rect 6876 2214 6894 2232
rect 6876 2232 6894 2250
rect 6876 2250 6894 2268
rect 6876 2268 6894 2286
rect 6876 2286 6894 2304
rect 6876 2304 6894 2322
rect 6876 2322 6894 2340
rect 6876 2340 6894 2358
rect 6876 2358 6894 2376
rect 6876 2376 6894 2394
rect 6876 2394 6894 2412
rect 6876 2412 6894 2430
rect 6876 2430 6894 2448
rect 6876 2448 6894 2466
rect 6876 2466 6894 2484
rect 6876 2484 6894 2502
rect 6876 2502 6894 2520
rect 6876 2520 6894 2538
rect 6876 2538 6894 2556
rect 6876 2556 6894 2574
rect 6876 2574 6894 2592
rect 6876 2592 6894 2610
rect 6876 2610 6894 2628
rect 6876 2628 6894 2646
rect 6876 2646 6894 2664
rect 6876 2664 6894 2682
rect 6876 2682 6894 2700
rect 6876 2700 6894 2718
rect 6876 2718 6894 2736
rect 6876 2736 6894 2754
rect 6876 2754 6894 2772
rect 6876 2772 6894 2790
rect 6876 2790 6894 2808
rect 6876 2808 6894 2826
rect 6876 2826 6894 2844
rect 6876 2844 6894 2862
rect 6876 2862 6894 2880
rect 6876 2880 6894 2898
rect 6876 2898 6894 2916
rect 6876 2916 6894 2934
rect 6876 2934 6894 2952
rect 6876 2952 6894 2970
rect 6876 2970 6894 2988
rect 6876 2988 6894 3006
rect 6876 3006 6894 3024
rect 6876 3024 6894 3042
rect 6876 3042 6894 3060
rect 6876 3222 6894 3240
rect 6876 3240 6894 3258
rect 6876 3258 6894 3276
rect 6876 3276 6894 3294
rect 6876 3294 6894 3312
rect 6876 3312 6894 3330
rect 6876 3330 6894 3348
rect 6876 3348 6894 3366
rect 6876 3366 6894 3384
rect 6876 3384 6894 3402
rect 6876 3402 6894 3420
rect 6876 3420 6894 3438
rect 6876 3438 6894 3456
rect 6876 3456 6894 3474
rect 6876 3474 6894 3492
rect 6876 3492 6894 3510
rect 6876 3510 6894 3528
rect 6876 3528 6894 3546
rect 6876 3546 6894 3564
rect 6876 3564 6894 3582
rect 6876 3582 6894 3600
rect 6876 3600 6894 3618
rect 6876 3618 6894 3636
rect 6876 3636 6894 3654
rect 6876 3654 6894 3672
rect 6876 3870 6894 3888
rect 6876 3888 6894 3906
rect 6876 3906 6894 3924
rect 6876 3924 6894 3942
rect 6876 3942 6894 3960
rect 6876 3960 6894 3978
rect 6876 3978 6894 3996
rect 6876 3996 6894 4014
rect 6876 4014 6894 4032
rect 6876 4032 6894 4050
rect 6876 4050 6894 4068
rect 6876 4068 6894 4086
rect 6876 4086 6894 4104
rect 6876 4104 6894 4122
rect 6876 4122 6894 4140
rect 6876 4140 6894 4158
rect 6876 4158 6894 4176
rect 6876 4176 6894 4194
rect 6876 4194 6894 4212
rect 6876 4212 6894 4230
rect 6876 4230 6894 4248
rect 6876 4248 6894 4266
rect 6876 4266 6894 4284
rect 6876 4284 6894 4302
rect 6876 4302 6894 4320
rect 6876 4320 6894 4338
rect 6876 4338 6894 4356
rect 6876 4356 6894 4374
rect 6876 4374 6894 4392
rect 6876 4392 6894 4410
rect 6876 4410 6894 4428
rect 6876 4428 6894 4446
rect 6876 4446 6894 4464
rect 6876 4464 6894 4482
rect 6876 4482 6894 4500
rect 6876 4500 6894 4518
rect 6876 4518 6894 4536
rect 6876 4536 6894 4554
rect 6876 4554 6894 4572
rect 6876 4572 6894 4590
rect 6876 4590 6894 4608
rect 6876 4608 6894 4626
rect 6876 4626 6894 4644
rect 6876 4644 6894 4662
rect 6876 4662 6894 4680
rect 6876 4680 6894 4698
rect 6876 4698 6894 4716
rect 6876 4716 6894 4734
rect 6876 4734 6894 4752
rect 6876 4752 6894 4770
rect 6876 4770 6894 4788
rect 6876 4788 6894 4806
rect 6876 4806 6894 4824
rect 6876 4824 6894 4842
rect 6876 4842 6894 4860
rect 6876 4860 6894 4878
rect 6876 4878 6894 4896
rect 6876 4896 6894 4914
rect 6876 4914 6894 4932
rect 6876 4932 6894 4950
rect 6876 4950 6894 4968
rect 6876 4968 6894 4986
rect 6876 4986 6894 5004
rect 6876 5004 6894 5022
rect 6876 5022 6894 5040
rect 6876 5040 6894 5058
rect 6876 5058 6894 5076
rect 6876 5076 6894 5094
rect 6876 5094 6894 5112
rect 6876 5112 6894 5130
rect 6876 5130 6894 5148
rect 6876 5148 6894 5166
rect 6876 5166 6894 5184
rect 6876 5184 6894 5202
rect 6876 5202 6894 5220
rect 6876 5220 6894 5238
rect 6876 5238 6894 5256
rect 6876 5256 6894 5274
rect 6876 5274 6894 5292
rect 6876 5292 6894 5310
rect 6876 5310 6894 5328
rect 6876 5328 6894 5346
rect 6876 5346 6894 5364
rect 6876 5364 6894 5382
rect 6876 5382 6894 5400
rect 6876 5400 6894 5418
rect 6876 5418 6894 5436
rect 6876 5436 6894 5454
rect 6876 5454 6894 5472
rect 6876 5472 6894 5490
rect 6876 5490 6894 5508
rect 6876 5508 6894 5526
rect 6876 5526 6894 5544
rect 6876 5544 6894 5562
rect 6876 5562 6894 5580
rect 6876 5580 6894 5598
rect 6876 5598 6894 5616
rect 6876 5616 6894 5634
rect 6876 5634 6894 5652
rect 6876 5652 6894 5670
rect 6876 5670 6894 5688
rect 6876 5688 6894 5706
rect 6876 5706 6894 5724
rect 6876 5724 6894 5742
rect 6876 5742 6894 5760
rect 6876 5760 6894 5778
rect 6876 5778 6894 5796
rect 6876 5796 6894 5814
rect 6876 5814 6894 5832
rect 6876 5832 6894 5850
rect 6876 5850 6894 5868
rect 6876 5868 6894 5886
rect 6876 5886 6894 5904
rect 6876 5904 6894 5922
rect 6876 5922 6894 5940
rect 6876 5940 6894 5958
rect 6876 5958 6894 5976
rect 6876 5976 6894 5994
rect 6876 5994 6894 6012
rect 6876 6012 6894 6030
rect 6876 6030 6894 6048
rect 6876 6048 6894 6066
rect 6876 6066 6894 6084
rect 6876 6084 6894 6102
rect 6876 6102 6894 6120
rect 6876 6120 6894 6138
rect 6876 6138 6894 6156
rect 6876 7524 6894 7542
rect 6876 7542 6894 7560
rect 6876 7560 6894 7578
rect 6876 7578 6894 7596
rect 6876 7596 6894 7614
rect 6876 7614 6894 7632
rect 6876 7632 6894 7650
rect 6876 7650 6894 7668
rect 6876 7668 6894 7686
rect 6876 7686 6894 7704
rect 6876 7704 6894 7722
rect 6876 7722 6894 7740
rect 6876 7740 6894 7758
rect 6876 7758 6894 7776
rect 6876 7776 6894 7794
rect 6876 7794 6894 7812
rect 6876 7812 6894 7830
rect 6876 7830 6894 7848
rect 6876 7848 6894 7866
rect 6876 7866 6894 7884
rect 6876 7884 6894 7902
rect 6876 7902 6894 7920
rect 6876 7920 6894 7938
rect 6876 7938 6894 7956
rect 6876 7956 6894 7974
rect 6876 7974 6894 7992
rect 6876 7992 6894 8010
rect 6876 8010 6894 8028
rect 6876 8028 6894 8046
rect 6876 8046 6894 8064
rect 6876 8064 6894 8082
rect 6876 8082 6894 8100
rect 6876 8100 6894 8118
rect 6876 8118 6894 8136
rect 6876 8136 6894 8154
rect 6876 8154 6894 8172
rect 6876 8172 6894 8190
rect 6876 8190 6894 8208
rect 6876 8208 6894 8226
rect 6876 8226 6894 8244
rect 6876 8244 6894 8262
rect 6876 8262 6894 8280
rect 6876 8280 6894 8298
rect 6876 8298 6894 8316
rect 6876 8316 6894 8334
rect 6876 8334 6894 8352
rect 6876 8352 6894 8370
rect 6876 8370 6894 8388
rect 6876 8388 6894 8406
rect 6876 8406 6894 8424
rect 6876 8424 6894 8442
rect 6876 8442 6894 8460
rect 6876 8460 6894 8478
rect 6876 8478 6894 8496
rect 6876 8496 6894 8514
rect 6876 8514 6894 8532
rect 6876 8532 6894 8550
rect 6876 8550 6894 8568
rect 6876 8568 6894 8586
rect 6876 8586 6894 8604
rect 6876 8604 6894 8622
rect 6876 8622 6894 8640
rect 6876 8640 6894 8658
rect 6876 8658 6894 8676
rect 6876 8676 6894 8694
rect 6876 8694 6894 8712
rect 6876 8712 6894 8730
rect 6876 8730 6894 8748
rect 6876 8748 6894 8766
rect 6876 8766 6894 8784
rect 6876 8784 6894 8802
rect 6876 8802 6894 8820
rect 6876 8820 6894 8838
rect 6876 8838 6894 8856
rect 6876 8856 6894 8874
rect 6876 8874 6894 8892
rect 6876 8892 6894 8910
rect 6876 8910 6894 8928
rect 6876 8928 6894 8946
rect 6876 8946 6894 8964
rect 6876 8964 6894 8982
rect 6876 8982 6894 9000
rect 6876 9000 6894 9018
rect 6876 9018 6894 9036
rect 6876 9036 6894 9054
rect 6876 9054 6894 9072
rect 6876 9072 6894 9090
rect 6876 9090 6894 9108
rect 6876 9108 6894 9126
rect 6876 9126 6894 9144
rect 6876 9144 6894 9162
rect 6876 9162 6894 9180
rect 6876 9180 6894 9198
rect 6876 9198 6894 9216
rect 6876 9216 6894 9234
rect 6876 9234 6894 9252
rect 6876 9252 6894 9270
rect 6876 9270 6894 9288
rect 6876 9288 6894 9306
rect 6876 9306 6894 9324
rect 6876 9324 6894 9342
rect 6876 9342 6894 9360
rect 6876 9360 6894 9378
rect 6876 9378 6894 9396
rect 6876 9396 6894 9414
rect 6876 9414 6894 9432
rect 6876 9432 6894 9450
rect 6876 9450 6894 9468
rect 6876 9468 6894 9486
rect 6876 9486 6894 9504
rect 6876 9504 6894 9522
rect 6876 9522 6894 9540
rect 6876 9540 6894 9558
rect 6876 9558 6894 9576
rect 6876 9576 6894 9594
rect 6876 9594 6894 9612
rect 6876 9612 6894 9630
rect 6876 9630 6894 9648
rect 6876 9648 6894 9666
rect 6876 9666 6894 9684
rect 6876 9684 6894 9702
rect 6876 9702 6894 9720
rect 6876 9720 6894 9738
rect 6876 9738 6894 9756
rect 6876 9756 6894 9774
rect 6876 9774 6894 9792
rect 6876 9792 6894 9810
rect 6876 9810 6894 9828
rect 6876 9828 6894 9846
rect 6876 9846 6894 9864
rect 6876 9864 6894 9882
rect 6876 9882 6894 9900
rect 6876 9900 6894 9918
rect 6876 9918 6894 9936
rect 6876 9936 6894 9954
rect 6876 9954 6894 9972
rect 6876 9972 6894 9990
rect 6876 9990 6894 10008
rect 6876 10008 6894 10026
rect 6876 10026 6894 10044
rect 6876 10044 6894 10062
rect 6876 10062 6894 10080
rect 6876 10080 6894 10098
rect 6876 10098 6894 10116
rect 6876 10116 6894 10134
rect 6876 10134 6894 10152
rect 6876 10152 6894 10170
rect 6876 10170 6894 10188
rect 6876 10188 6894 10206
rect 6876 10206 6894 10224
rect 6876 10224 6894 10242
rect 6876 10242 6894 10260
rect 6876 10260 6894 10278
rect 6876 10278 6894 10296
rect 6876 10296 6894 10314
rect 6876 10314 6894 10332
rect 6894 1728 6912 1746
rect 6894 1746 6912 1764
rect 6894 1764 6912 1782
rect 6894 1782 6912 1800
rect 6894 1800 6912 1818
rect 6894 1818 6912 1836
rect 6894 1836 6912 1854
rect 6894 1854 6912 1872
rect 6894 1872 6912 1890
rect 6894 1890 6912 1908
rect 6894 1908 6912 1926
rect 6894 1926 6912 1944
rect 6894 1944 6912 1962
rect 6894 1962 6912 1980
rect 6894 1980 6912 1998
rect 6894 1998 6912 2016
rect 6894 2016 6912 2034
rect 6894 2034 6912 2052
rect 6894 2052 6912 2070
rect 6894 2070 6912 2088
rect 6894 2088 6912 2106
rect 6894 2106 6912 2124
rect 6894 2124 6912 2142
rect 6894 2142 6912 2160
rect 6894 2160 6912 2178
rect 6894 2178 6912 2196
rect 6894 2196 6912 2214
rect 6894 2214 6912 2232
rect 6894 2232 6912 2250
rect 6894 2250 6912 2268
rect 6894 2268 6912 2286
rect 6894 2286 6912 2304
rect 6894 2304 6912 2322
rect 6894 2322 6912 2340
rect 6894 2340 6912 2358
rect 6894 2358 6912 2376
rect 6894 2376 6912 2394
rect 6894 2394 6912 2412
rect 6894 2412 6912 2430
rect 6894 2430 6912 2448
rect 6894 2448 6912 2466
rect 6894 2466 6912 2484
rect 6894 2484 6912 2502
rect 6894 2502 6912 2520
rect 6894 2520 6912 2538
rect 6894 2538 6912 2556
rect 6894 2556 6912 2574
rect 6894 2574 6912 2592
rect 6894 2592 6912 2610
rect 6894 2610 6912 2628
rect 6894 2628 6912 2646
rect 6894 2646 6912 2664
rect 6894 2664 6912 2682
rect 6894 2682 6912 2700
rect 6894 2700 6912 2718
rect 6894 2718 6912 2736
rect 6894 2736 6912 2754
rect 6894 2754 6912 2772
rect 6894 2772 6912 2790
rect 6894 2790 6912 2808
rect 6894 2808 6912 2826
rect 6894 2826 6912 2844
rect 6894 2844 6912 2862
rect 6894 2862 6912 2880
rect 6894 2880 6912 2898
rect 6894 2898 6912 2916
rect 6894 2916 6912 2934
rect 6894 2934 6912 2952
rect 6894 2952 6912 2970
rect 6894 2970 6912 2988
rect 6894 2988 6912 3006
rect 6894 3006 6912 3024
rect 6894 3024 6912 3042
rect 6894 3042 6912 3060
rect 6894 3240 6912 3258
rect 6894 3258 6912 3276
rect 6894 3276 6912 3294
rect 6894 3294 6912 3312
rect 6894 3312 6912 3330
rect 6894 3330 6912 3348
rect 6894 3348 6912 3366
rect 6894 3366 6912 3384
rect 6894 3384 6912 3402
rect 6894 3402 6912 3420
rect 6894 3420 6912 3438
rect 6894 3438 6912 3456
rect 6894 3456 6912 3474
rect 6894 3474 6912 3492
rect 6894 3492 6912 3510
rect 6894 3510 6912 3528
rect 6894 3528 6912 3546
rect 6894 3546 6912 3564
rect 6894 3564 6912 3582
rect 6894 3582 6912 3600
rect 6894 3600 6912 3618
rect 6894 3618 6912 3636
rect 6894 3636 6912 3654
rect 6894 3654 6912 3672
rect 6894 3672 6912 3690
rect 6894 3906 6912 3924
rect 6894 3924 6912 3942
rect 6894 3942 6912 3960
rect 6894 3960 6912 3978
rect 6894 3978 6912 3996
rect 6894 3996 6912 4014
rect 6894 4014 6912 4032
rect 6894 4032 6912 4050
rect 6894 4050 6912 4068
rect 6894 4068 6912 4086
rect 6894 4086 6912 4104
rect 6894 4104 6912 4122
rect 6894 4122 6912 4140
rect 6894 4140 6912 4158
rect 6894 4158 6912 4176
rect 6894 4176 6912 4194
rect 6894 4194 6912 4212
rect 6894 4212 6912 4230
rect 6894 4230 6912 4248
rect 6894 4248 6912 4266
rect 6894 4266 6912 4284
rect 6894 4284 6912 4302
rect 6894 4302 6912 4320
rect 6894 4320 6912 4338
rect 6894 4338 6912 4356
rect 6894 4356 6912 4374
rect 6894 4374 6912 4392
rect 6894 4392 6912 4410
rect 6894 4410 6912 4428
rect 6894 4428 6912 4446
rect 6894 4446 6912 4464
rect 6894 4464 6912 4482
rect 6894 4482 6912 4500
rect 6894 4500 6912 4518
rect 6894 4518 6912 4536
rect 6894 4536 6912 4554
rect 6894 4554 6912 4572
rect 6894 4572 6912 4590
rect 6894 4590 6912 4608
rect 6894 4608 6912 4626
rect 6894 4626 6912 4644
rect 6894 4644 6912 4662
rect 6894 4662 6912 4680
rect 6894 4680 6912 4698
rect 6894 4698 6912 4716
rect 6894 4716 6912 4734
rect 6894 4734 6912 4752
rect 6894 4752 6912 4770
rect 6894 4770 6912 4788
rect 6894 4788 6912 4806
rect 6894 4806 6912 4824
rect 6894 4824 6912 4842
rect 6894 4842 6912 4860
rect 6894 4860 6912 4878
rect 6894 4878 6912 4896
rect 6894 4896 6912 4914
rect 6894 4914 6912 4932
rect 6894 4932 6912 4950
rect 6894 4950 6912 4968
rect 6894 4968 6912 4986
rect 6894 4986 6912 5004
rect 6894 5004 6912 5022
rect 6894 5022 6912 5040
rect 6894 5040 6912 5058
rect 6894 5058 6912 5076
rect 6894 5076 6912 5094
rect 6894 5094 6912 5112
rect 6894 5112 6912 5130
rect 6894 5130 6912 5148
rect 6894 5148 6912 5166
rect 6894 5166 6912 5184
rect 6894 5184 6912 5202
rect 6894 5202 6912 5220
rect 6894 5220 6912 5238
rect 6894 5238 6912 5256
rect 6894 5256 6912 5274
rect 6894 5274 6912 5292
rect 6894 5292 6912 5310
rect 6894 5310 6912 5328
rect 6894 5328 6912 5346
rect 6894 5346 6912 5364
rect 6894 5364 6912 5382
rect 6894 5382 6912 5400
rect 6894 5400 6912 5418
rect 6894 5418 6912 5436
rect 6894 5436 6912 5454
rect 6894 5454 6912 5472
rect 6894 5472 6912 5490
rect 6894 5490 6912 5508
rect 6894 5508 6912 5526
rect 6894 5526 6912 5544
rect 6894 5544 6912 5562
rect 6894 5562 6912 5580
rect 6894 5580 6912 5598
rect 6894 5598 6912 5616
rect 6894 5616 6912 5634
rect 6894 5634 6912 5652
rect 6894 5652 6912 5670
rect 6894 5670 6912 5688
rect 6894 5688 6912 5706
rect 6894 5706 6912 5724
rect 6894 5724 6912 5742
rect 6894 5742 6912 5760
rect 6894 5760 6912 5778
rect 6894 5778 6912 5796
rect 6894 5796 6912 5814
rect 6894 5814 6912 5832
rect 6894 5832 6912 5850
rect 6894 5850 6912 5868
rect 6894 5868 6912 5886
rect 6894 5886 6912 5904
rect 6894 5904 6912 5922
rect 6894 5922 6912 5940
rect 6894 5940 6912 5958
rect 6894 5958 6912 5976
rect 6894 5976 6912 5994
rect 6894 5994 6912 6012
rect 6894 6012 6912 6030
rect 6894 6030 6912 6048
rect 6894 6048 6912 6066
rect 6894 6066 6912 6084
rect 6894 6084 6912 6102
rect 6894 6102 6912 6120
rect 6894 6120 6912 6138
rect 6894 6138 6912 6156
rect 6894 6156 6912 6174
rect 6894 7578 6912 7596
rect 6894 7596 6912 7614
rect 6894 7614 6912 7632
rect 6894 7632 6912 7650
rect 6894 7650 6912 7668
rect 6894 7668 6912 7686
rect 6894 7686 6912 7704
rect 6894 7704 6912 7722
rect 6894 7722 6912 7740
rect 6894 7740 6912 7758
rect 6894 7758 6912 7776
rect 6894 7776 6912 7794
rect 6894 7794 6912 7812
rect 6894 7812 6912 7830
rect 6894 7830 6912 7848
rect 6894 7848 6912 7866
rect 6894 7866 6912 7884
rect 6894 7884 6912 7902
rect 6894 7902 6912 7920
rect 6894 7920 6912 7938
rect 6894 7938 6912 7956
rect 6894 7956 6912 7974
rect 6894 7974 6912 7992
rect 6894 7992 6912 8010
rect 6894 8010 6912 8028
rect 6894 8028 6912 8046
rect 6894 8046 6912 8064
rect 6894 8064 6912 8082
rect 6894 8082 6912 8100
rect 6894 8100 6912 8118
rect 6894 8118 6912 8136
rect 6894 8136 6912 8154
rect 6894 8154 6912 8172
rect 6894 8172 6912 8190
rect 6894 8190 6912 8208
rect 6894 8208 6912 8226
rect 6894 8226 6912 8244
rect 6894 8244 6912 8262
rect 6894 8262 6912 8280
rect 6894 8280 6912 8298
rect 6894 8298 6912 8316
rect 6894 8316 6912 8334
rect 6894 8334 6912 8352
rect 6894 8352 6912 8370
rect 6894 8370 6912 8388
rect 6894 8388 6912 8406
rect 6894 8406 6912 8424
rect 6894 8424 6912 8442
rect 6894 8442 6912 8460
rect 6894 8460 6912 8478
rect 6894 8478 6912 8496
rect 6894 8496 6912 8514
rect 6894 8514 6912 8532
rect 6894 8532 6912 8550
rect 6894 8550 6912 8568
rect 6894 8568 6912 8586
rect 6894 8586 6912 8604
rect 6894 8604 6912 8622
rect 6894 8622 6912 8640
rect 6894 8640 6912 8658
rect 6894 8658 6912 8676
rect 6894 8676 6912 8694
rect 6894 8694 6912 8712
rect 6894 8712 6912 8730
rect 6894 8730 6912 8748
rect 6894 8748 6912 8766
rect 6894 8766 6912 8784
rect 6894 8784 6912 8802
rect 6894 8802 6912 8820
rect 6894 8820 6912 8838
rect 6894 8838 6912 8856
rect 6894 8856 6912 8874
rect 6894 8874 6912 8892
rect 6894 8892 6912 8910
rect 6894 8910 6912 8928
rect 6894 8928 6912 8946
rect 6894 8946 6912 8964
rect 6894 8964 6912 8982
rect 6894 8982 6912 9000
rect 6894 9000 6912 9018
rect 6894 9018 6912 9036
rect 6894 9036 6912 9054
rect 6894 9054 6912 9072
rect 6894 9072 6912 9090
rect 6894 9090 6912 9108
rect 6894 9108 6912 9126
rect 6894 9126 6912 9144
rect 6894 9144 6912 9162
rect 6894 9162 6912 9180
rect 6894 9180 6912 9198
rect 6894 9198 6912 9216
rect 6894 9216 6912 9234
rect 6894 9234 6912 9252
rect 6894 9252 6912 9270
rect 6894 9270 6912 9288
rect 6894 9288 6912 9306
rect 6894 9306 6912 9324
rect 6894 9324 6912 9342
rect 6894 9342 6912 9360
rect 6894 9360 6912 9378
rect 6894 9378 6912 9396
rect 6894 9396 6912 9414
rect 6894 9414 6912 9432
rect 6894 9432 6912 9450
rect 6894 9450 6912 9468
rect 6894 9468 6912 9486
rect 6894 9486 6912 9504
rect 6894 9504 6912 9522
rect 6894 9522 6912 9540
rect 6894 9540 6912 9558
rect 6894 9558 6912 9576
rect 6894 9576 6912 9594
rect 6894 9594 6912 9612
rect 6894 9612 6912 9630
rect 6894 9630 6912 9648
rect 6894 9648 6912 9666
rect 6894 9666 6912 9684
rect 6894 9684 6912 9702
rect 6894 9702 6912 9720
rect 6894 9720 6912 9738
rect 6894 9738 6912 9756
rect 6894 9756 6912 9774
rect 6894 9774 6912 9792
rect 6894 9792 6912 9810
rect 6894 9810 6912 9828
rect 6894 9828 6912 9846
rect 6894 9846 6912 9864
rect 6894 9864 6912 9882
rect 6894 9882 6912 9900
rect 6894 9900 6912 9918
rect 6894 9918 6912 9936
rect 6894 9936 6912 9954
rect 6894 9954 6912 9972
rect 6894 9972 6912 9990
rect 6894 9990 6912 10008
rect 6894 10008 6912 10026
rect 6894 10026 6912 10044
rect 6894 10044 6912 10062
rect 6894 10062 6912 10080
rect 6894 10080 6912 10098
rect 6894 10098 6912 10116
rect 6894 10116 6912 10134
rect 6894 10134 6912 10152
rect 6894 10152 6912 10170
rect 6894 10170 6912 10188
rect 6894 10188 6912 10206
rect 6894 10206 6912 10224
rect 6894 10224 6912 10242
rect 6894 10242 6912 10260
rect 6894 10260 6912 10278
rect 6894 10278 6912 10296
rect 6894 10296 6912 10314
rect 6894 10314 6912 10332
rect 6894 10332 6912 10350
rect 6912 1728 6930 1746
rect 6912 1746 6930 1764
rect 6912 1764 6930 1782
rect 6912 1782 6930 1800
rect 6912 1800 6930 1818
rect 6912 1818 6930 1836
rect 6912 1836 6930 1854
rect 6912 1854 6930 1872
rect 6912 1872 6930 1890
rect 6912 1890 6930 1908
rect 6912 1908 6930 1926
rect 6912 1926 6930 1944
rect 6912 1944 6930 1962
rect 6912 1962 6930 1980
rect 6912 1980 6930 1998
rect 6912 1998 6930 2016
rect 6912 2016 6930 2034
rect 6912 2034 6930 2052
rect 6912 2052 6930 2070
rect 6912 2070 6930 2088
rect 6912 2088 6930 2106
rect 6912 2106 6930 2124
rect 6912 2124 6930 2142
rect 6912 2142 6930 2160
rect 6912 2160 6930 2178
rect 6912 2178 6930 2196
rect 6912 2196 6930 2214
rect 6912 2214 6930 2232
rect 6912 2232 6930 2250
rect 6912 2250 6930 2268
rect 6912 2268 6930 2286
rect 6912 2286 6930 2304
rect 6912 2304 6930 2322
rect 6912 2322 6930 2340
rect 6912 2340 6930 2358
rect 6912 2358 6930 2376
rect 6912 2376 6930 2394
rect 6912 2394 6930 2412
rect 6912 2412 6930 2430
rect 6912 2430 6930 2448
rect 6912 2448 6930 2466
rect 6912 2466 6930 2484
rect 6912 2484 6930 2502
rect 6912 2502 6930 2520
rect 6912 2520 6930 2538
rect 6912 2538 6930 2556
rect 6912 2556 6930 2574
rect 6912 2574 6930 2592
rect 6912 2592 6930 2610
rect 6912 2610 6930 2628
rect 6912 2628 6930 2646
rect 6912 2646 6930 2664
rect 6912 2664 6930 2682
rect 6912 2682 6930 2700
rect 6912 2700 6930 2718
rect 6912 2718 6930 2736
rect 6912 2736 6930 2754
rect 6912 2754 6930 2772
rect 6912 2772 6930 2790
rect 6912 2790 6930 2808
rect 6912 2808 6930 2826
rect 6912 2826 6930 2844
rect 6912 2844 6930 2862
rect 6912 2862 6930 2880
rect 6912 2880 6930 2898
rect 6912 2898 6930 2916
rect 6912 2916 6930 2934
rect 6912 2934 6930 2952
rect 6912 2952 6930 2970
rect 6912 2970 6930 2988
rect 6912 2988 6930 3006
rect 6912 3006 6930 3024
rect 6912 3024 6930 3042
rect 6912 3042 6930 3060
rect 6912 3240 6930 3258
rect 6912 3258 6930 3276
rect 6912 3276 6930 3294
rect 6912 3294 6930 3312
rect 6912 3312 6930 3330
rect 6912 3330 6930 3348
rect 6912 3348 6930 3366
rect 6912 3366 6930 3384
rect 6912 3384 6930 3402
rect 6912 3402 6930 3420
rect 6912 3420 6930 3438
rect 6912 3438 6930 3456
rect 6912 3456 6930 3474
rect 6912 3474 6930 3492
rect 6912 3492 6930 3510
rect 6912 3510 6930 3528
rect 6912 3528 6930 3546
rect 6912 3546 6930 3564
rect 6912 3564 6930 3582
rect 6912 3582 6930 3600
rect 6912 3600 6930 3618
rect 6912 3618 6930 3636
rect 6912 3636 6930 3654
rect 6912 3654 6930 3672
rect 6912 3672 6930 3690
rect 6912 3690 6930 3708
rect 6912 3708 6930 3726
rect 6912 3924 6930 3942
rect 6912 3942 6930 3960
rect 6912 3960 6930 3978
rect 6912 3978 6930 3996
rect 6912 3996 6930 4014
rect 6912 4014 6930 4032
rect 6912 4032 6930 4050
rect 6912 4050 6930 4068
rect 6912 4068 6930 4086
rect 6912 4086 6930 4104
rect 6912 4104 6930 4122
rect 6912 4122 6930 4140
rect 6912 4140 6930 4158
rect 6912 4158 6930 4176
rect 6912 4176 6930 4194
rect 6912 4194 6930 4212
rect 6912 4212 6930 4230
rect 6912 4230 6930 4248
rect 6912 4248 6930 4266
rect 6912 4266 6930 4284
rect 6912 4284 6930 4302
rect 6912 4302 6930 4320
rect 6912 4320 6930 4338
rect 6912 4338 6930 4356
rect 6912 4356 6930 4374
rect 6912 4374 6930 4392
rect 6912 4392 6930 4410
rect 6912 4410 6930 4428
rect 6912 4428 6930 4446
rect 6912 4446 6930 4464
rect 6912 4464 6930 4482
rect 6912 4482 6930 4500
rect 6912 4500 6930 4518
rect 6912 4518 6930 4536
rect 6912 4536 6930 4554
rect 6912 4554 6930 4572
rect 6912 4572 6930 4590
rect 6912 4590 6930 4608
rect 6912 4608 6930 4626
rect 6912 4626 6930 4644
rect 6912 4644 6930 4662
rect 6912 4662 6930 4680
rect 6912 4680 6930 4698
rect 6912 4698 6930 4716
rect 6912 4716 6930 4734
rect 6912 4734 6930 4752
rect 6912 4752 6930 4770
rect 6912 4770 6930 4788
rect 6912 4788 6930 4806
rect 6912 4806 6930 4824
rect 6912 4824 6930 4842
rect 6912 4842 6930 4860
rect 6912 4860 6930 4878
rect 6912 4878 6930 4896
rect 6912 4896 6930 4914
rect 6912 4914 6930 4932
rect 6912 4932 6930 4950
rect 6912 4950 6930 4968
rect 6912 4968 6930 4986
rect 6912 4986 6930 5004
rect 6912 5004 6930 5022
rect 6912 5022 6930 5040
rect 6912 5040 6930 5058
rect 6912 5058 6930 5076
rect 6912 5076 6930 5094
rect 6912 5094 6930 5112
rect 6912 5112 6930 5130
rect 6912 5130 6930 5148
rect 6912 5148 6930 5166
rect 6912 5166 6930 5184
rect 6912 5184 6930 5202
rect 6912 5202 6930 5220
rect 6912 5220 6930 5238
rect 6912 5238 6930 5256
rect 6912 5256 6930 5274
rect 6912 5274 6930 5292
rect 6912 5292 6930 5310
rect 6912 5310 6930 5328
rect 6912 5328 6930 5346
rect 6912 5346 6930 5364
rect 6912 5364 6930 5382
rect 6912 5382 6930 5400
rect 6912 5400 6930 5418
rect 6912 5418 6930 5436
rect 6912 5436 6930 5454
rect 6912 5454 6930 5472
rect 6912 5472 6930 5490
rect 6912 5490 6930 5508
rect 6912 5508 6930 5526
rect 6912 5526 6930 5544
rect 6912 5544 6930 5562
rect 6912 5562 6930 5580
rect 6912 5580 6930 5598
rect 6912 5598 6930 5616
rect 6912 5616 6930 5634
rect 6912 5634 6930 5652
rect 6912 5652 6930 5670
rect 6912 5670 6930 5688
rect 6912 5688 6930 5706
rect 6912 5706 6930 5724
rect 6912 5724 6930 5742
rect 6912 5742 6930 5760
rect 6912 5760 6930 5778
rect 6912 5778 6930 5796
rect 6912 5796 6930 5814
rect 6912 5814 6930 5832
rect 6912 5832 6930 5850
rect 6912 5850 6930 5868
rect 6912 5868 6930 5886
rect 6912 5886 6930 5904
rect 6912 5904 6930 5922
rect 6912 5922 6930 5940
rect 6912 5940 6930 5958
rect 6912 5958 6930 5976
rect 6912 5976 6930 5994
rect 6912 5994 6930 6012
rect 6912 6012 6930 6030
rect 6912 6030 6930 6048
rect 6912 6048 6930 6066
rect 6912 6066 6930 6084
rect 6912 6084 6930 6102
rect 6912 6102 6930 6120
rect 6912 6120 6930 6138
rect 6912 6138 6930 6156
rect 6912 6156 6930 6174
rect 6912 6174 6930 6192
rect 6912 7632 6930 7650
rect 6912 7650 6930 7668
rect 6912 7668 6930 7686
rect 6912 7686 6930 7704
rect 6912 7704 6930 7722
rect 6912 7722 6930 7740
rect 6912 7740 6930 7758
rect 6912 7758 6930 7776
rect 6912 7776 6930 7794
rect 6912 7794 6930 7812
rect 6912 7812 6930 7830
rect 6912 7830 6930 7848
rect 6912 7848 6930 7866
rect 6912 7866 6930 7884
rect 6912 7884 6930 7902
rect 6912 7902 6930 7920
rect 6912 7920 6930 7938
rect 6912 7938 6930 7956
rect 6912 7956 6930 7974
rect 6912 7974 6930 7992
rect 6912 7992 6930 8010
rect 6912 8010 6930 8028
rect 6912 8028 6930 8046
rect 6912 8046 6930 8064
rect 6912 8064 6930 8082
rect 6912 8082 6930 8100
rect 6912 8100 6930 8118
rect 6912 8118 6930 8136
rect 6912 8136 6930 8154
rect 6912 8154 6930 8172
rect 6912 8172 6930 8190
rect 6912 8190 6930 8208
rect 6912 8208 6930 8226
rect 6912 8226 6930 8244
rect 6912 8244 6930 8262
rect 6912 8262 6930 8280
rect 6912 8280 6930 8298
rect 6912 8298 6930 8316
rect 6912 8316 6930 8334
rect 6912 8334 6930 8352
rect 6912 8352 6930 8370
rect 6912 8370 6930 8388
rect 6912 8388 6930 8406
rect 6912 8406 6930 8424
rect 6912 8424 6930 8442
rect 6912 8442 6930 8460
rect 6912 8460 6930 8478
rect 6912 8478 6930 8496
rect 6912 8496 6930 8514
rect 6912 8514 6930 8532
rect 6912 8532 6930 8550
rect 6912 8550 6930 8568
rect 6912 8568 6930 8586
rect 6912 8586 6930 8604
rect 6912 8604 6930 8622
rect 6912 8622 6930 8640
rect 6912 8640 6930 8658
rect 6912 8658 6930 8676
rect 6912 8676 6930 8694
rect 6912 8694 6930 8712
rect 6912 8712 6930 8730
rect 6912 8730 6930 8748
rect 6912 8748 6930 8766
rect 6912 8766 6930 8784
rect 6912 8784 6930 8802
rect 6912 8802 6930 8820
rect 6912 8820 6930 8838
rect 6912 8838 6930 8856
rect 6912 8856 6930 8874
rect 6912 8874 6930 8892
rect 6912 8892 6930 8910
rect 6912 8910 6930 8928
rect 6912 8928 6930 8946
rect 6912 8946 6930 8964
rect 6912 8964 6930 8982
rect 6912 8982 6930 9000
rect 6912 9000 6930 9018
rect 6912 9018 6930 9036
rect 6912 9036 6930 9054
rect 6912 9054 6930 9072
rect 6912 9072 6930 9090
rect 6912 9090 6930 9108
rect 6912 9108 6930 9126
rect 6912 9126 6930 9144
rect 6912 9144 6930 9162
rect 6912 9162 6930 9180
rect 6912 9180 6930 9198
rect 6912 9198 6930 9216
rect 6912 9216 6930 9234
rect 6912 9234 6930 9252
rect 6912 9252 6930 9270
rect 6912 9270 6930 9288
rect 6912 9288 6930 9306
rect 6912 9306 6930 9324
rect 6912 9324 6930 9342
rect 6912 9342 6930 9360
rect 6912 9360 6930 9378
rect 6912 9378 6930 9396
rect 6912 9396 6930 9414
rect 6912 9414 6930 9432
rect 6912 9432 6930 9450
rect 6912 9450 6930 9468
rect 6912 9468 6930 9486
rect 6912 9486 6930 9504
rect 6912 9504 6930 9522
rect 6912 9522 6930 9540
rect 6912 9540 6930 9558
rect 6912 9558 6930 9576
rect 6912 9576 6930 9594
rect 6912 9594 6930 9612
rect 6912 9612 6930 9630
rect 6912 9630 6930 9648
rect 6912 9648 6930 9666
rect 6912 9666 6930 9684
rect 6912 9684 6930 9702
rect 6912 9702 6930 9720
rect 6912 9720 6930 9738
rect 6912 9738 6930 9756
rect 6912 9756 6930 9774
rect 6912 9774 6930 9792
rect 6912 9792 6930 9810
rect 6912 9810 6930 9828
rect 6912 9828 6930 9846
rect 6912 9846 6930 9864
rect 6912 9864 6930 9882
rect 6912 9882 6930 9900
rect 6912 9900 6930 9918
rect 6912 9918 6930 9936
rect 6912 9936 6930 9954
rect 6912 9954 6930 9972
rect 6912 9972 6930 9990
rect 6912 9990 6930 10008
rect 6912 10008 6930 10026
rect 6912 10026 6930 10044
rect 6912 10044 6930 10062
rect 6912 10062 6930 10080
rect 6912 10080 6930 10098
rect 6912 10098 6930 10116
rect 6912 10116 6930 10134
rect 6912 10134 6930 10152
rect 6912 10152 6930 10170
rect 6912 10170 6930 10188
rect 6912 10188 6930 10206
rect 6912 10206 6930 10224
rect 6912 10224 6930 10242
rect 6912 10242 6930 10260
rect 6912 10260 6930 10278
rect 6912 10278 6930 10296
rect 6912 10296 6930 10314
rect 6912 10314 6930 10332
rect 6912 10332 6930 10350
rect 6912 10350 6930 10368
rect 6930 1746 6948 1764
rect 6930 1764 6948 1782
rect 6930 1782 6948 1800
rect 6930 1800 6948 1818
rect 6930 1818 6948 1836
rect 6930 1836 6948 1854
rect 6930 1854 6948 1872
rect 6930 1872 6948 1890
rect 6930 1890 6948 1908
rect 6930 1908 6948 1926
rect 6930 1926 6948 1944
rect 6930 1944 6948 1962
rect 6930 1962 6948 1980
rect 6930 1980 6948 1998
rect 6930 1998 6948 2016
rect 6930 2016 6948 2034
rect 6930 2034 6948 2052
rect 6930 2052 6948 2070
rect 6930 2070 6948 2088
rect 6930 2088 6948 2106
rect 6930 2106 6948 2124
rect 6930 2124 6948 2142
rect 6930 2142 6948 2160
rect 6930 2160 6948 2178
rect 6930 2178 6948 2196
rect 6930 2196 6948 2214
rect 6930 2214 6948 2232
rect 6930 2232 6948 2250
rect 6930 2250 6948 2268
rect 6930 2268 6948 2286
rect 6930 2286 6948 2304
rect 6930 2304 6948 2322
rect 6930 2322 6948 2340
rect 6930 2340 6948 2358
rect 6930 2358 6948 2376
rect 6930 2376 6948 2394
rect 6930 2394 6948 2412
rect 6930 2412 6948 2430
rect 6930 2430 6948 2448
rect 6930 2448 6948 2466
rect 6930 2466 6948 2484
rect 6930 2484 6948 2502
rect 6930 2502 6948 2520
rect 6930 2520 6948 2538
rect 6930 2538 6948 2556
rect 6930 2556 6948 2574
rect 6930 2574 6948 2592
rect 6930 2592 6948 2610
rect 6930 2610 6948 2628
rect 6930 2628 6948 2646
rect 6930 2646 6948 2664
rect 6930 2664 6948 2682
rect 6930 2682 6948 2700
rect 6930 2700 6948 2718
rect 6930 2718 6948 2736
rect 6930 2736 6948 2754
rect 6930 2754 6948 2772
rect 6930 2772 6948 2790
rect 6930 2790 6948 2808
rect 6930 2808 6948 2826
rect 6930 2826 6948 2844
rect 6930 2844 6948 2862
rect 6930 2862 6948 2880
rect 6930 2880 6948 2898
rect 6930 2898 6948 2916
rect 6930 2916 6948 2934
rect 6930 2934 6948 2952
rect 6930 2952 6948 2970
rect 6930 2970 6948 2988
rect 6930 2988 6948 3006
rect 6930 3006 6948 3024
rect 6930 3024 6948 3042
rect 6930 3042 6948 3060
rect 6930 3060 6948 3078
rect 6930 3240 6948 3258
rect 6930 3258 6948 3276
rect 6930 3276 6948 3294
rect 6930 3294 6948 3312
rect 6930 3312 6948 3330
rect 6930 3330 6948 3348
rect 6930 3348 6948 3366
rect 6930 3366 6948 3384
rect 6930 3384 6948 3402
rect 6930 3402 6948 3420
rect 6930 3420 6948 3438
rect 6930 3438 6948 3456
rect 6930 3456 6948 3474
rect 6930 3474 6948 3492
rect 6930 3492 6948 3510
rect 6930 3510 6948 3528
rect 6930 3528 6948 3546
rect 6930 3546 6948 3564
rect 6930 3564 6948 3582
rect 6930 3582 6948 3600
rect 6930 3600 6948 3618
rect 6930 3618 6948 3636
rect 6930 3636 6948 3654
rect 6930 3654 6948 3672
rect 6930 3672 6948 3690
rect 6930 3690 6948 3708
rect 6930 3708 6948 3726
rect 6930 3726 6948 3744
rect 6930 3942 6948 3960
rect 6930 3960 6948 3978
rect 6930 3978 6948 3996
rect 6930 3996 6948 4014
rect 6930 4014 6948 4032
rect 6930 4032 6948 4050
rect 6930 4050 6948 4068
rect 6930 4068 6948 4086
rect 6930 4086 6948 4104
rect 6930 4104 6948 4122
rect 6930 4122 6948 4140
rect 6930 4140 6948 4158
rect 6930 4158 6948 4176
rect 6930 4176 6948 4194
rect 6930 4194 6948 4212
rect 6930 4212 6948 4230
rect 6930 4230 6948 4248
rect 6930 4248 6948 4266
rect 6930 4266 6948 4284
rect 6930 4284 6948 4302
rect 6930 4302 6948 4320
rect 6930 4320 6948 4338
rect 6930 4338 6948 4356
rect 6930 4356 6948 4374
rect 6930 4374 6948 4392
rect 6930 4392 6948 4410
rect 6930 4410 6948 4428
rect 6930 4428 6948 4446
rect 6930 4446 6948 4464
rect 6930 4464 6948 4482
rect 6930 4482 6948 4500
rect 6930 4500 6948 4518
rect 6930 4518 6948 4536
rect 6930 4536 6948 4554
rect 6930 4554 6948 4572
rect 6930 4572 6948 4590
rect 6930 4590 6948 4608
rect 6930 4608 6948 4626
rect 6930 4626 6948 4644
rect 6930 4644 6948 4662
rect 6930 4662 6948 4680
rect 6930 4680 6948 4698
rect 6930 4698 6948 4716
rect 6930 4716 6948 4734
rect 6930 4734 6948 4752
rect 6930 4752 6948 4770
rect 6930 4770 6948 4788
rect 6930 4788 6948 4806
rect 6930 4806 6948 4824
rect 6930 4824 6948 4842
rect 6930 4842 6948 4860
rect 6930 4860 6948 4878
rect 6930 4878 6948 4896
rect 6930 4896 6948 4914
rect 6930 4914 6948 4932
rect 6930 4932 6948 4950
rect 6930 4950 6948 4968
rect 6930 4968 6948 4986
rect 6930 4986 6948 5004
rect 6930 5004 6948 5022
rect 6930 5022 6948 5040
rect 6930 5040 6948 5058
rect 6930 5058 6948 5076
rect 6930 5076 6948 5094
rect 6930 5094 6948 5112
rect 6930 5112 6948 5130
rect 6930 5130 6948 5148
rect 6930 5148 6948 5166
rect 6930 5166 6948 5184
rect 6930 5184 6948 5202
rect 6930 5202 6948 5220
rect 6930 5220 6948 5238
rect 6930 5238 6948 5256
rect 6930 5256 6948 5274
rect 6930 5274 6948 5292
rect 6930 5292 6948 5310
rect 6930 5310 6948 5328
rect 6930 5328 6948 5346
rect 6930 5346 6948 5364
rect 6930 5364 6948 5382
rect 6930 5382 6948 5400
rect 6930 5400 6948 5418
rect 6930 5418 6948 5436
rect 6930 5436 6948 5454
rect 6930 5454 6948 5472
rect 6930 5472 6948 5490
rect 6930 5490 6948 5508
rect 6930 5508 6948 5526
rect 6930 5526 6948 5544
rect 6930 5544 6948 5562
rect 6930 5562 6948 5580
rect 6930 5580 6948 5598
rect 6930 5598 6948 5616
rect 6930 5616 6948 5634
rect 6930 5634 6948 5652
rect 6930 5652 6948 5670
rect 6930 5670 6948 5688
rect 6930 5688 6948 5706
rect 6930 5706 6948 5724
rect 6930 5724 6948 5742
rect 6930 5742 6948 5760
rect 6930 5760 6948 5778
rect 6930 5778 6948 5796
rect 6930 5796 6948 5814
rect 6930 5814 6948 5832
rect 6930 5832 6948 5850
rect 6930 5850 6948 5868
rect 6930 5868 6948 5886
rect 6930 5886 6948 5904
rect 6930 5904 6948 5922
rect 6930 5922 6948 5940
rect 6930 5940 6948 5958
rect 6930 5958 6948 5976
rect 6930 5976 6948 5994
rect 6930 5994 6948 6012
rect 6930 6012 6948 6030
rect 6930 6030 6948 6048
rect 6930 6048 6948 6066
rect 6930 6066 6948 6084
rect 6930 6084 6948 6102
rect 6930 6102 6948 6120
rect 6930 6120 6948 6138
rect 6930 6138 6948 6156
rect 6930 6156 6948 6174
rect 6930 6174 6948 6192
rect 6930 6192 6948 6210
rect 6930 7668 6948 7686
rect 6930 7686 6948 7704
rect 6930 7704 6948 7722
rect 6930 7722 6948 7740
rect 6930 7740 6948 7758
rect 6930 7758 6948 7776
rect 6930 7776 6948 7794
rect 6930 7794 6948 7812
rect 6930 7812 6948 7830
rect 6930 7830 6948 7848
rect 6930 7848 6948 7866
rect 6930 7866 6948 7884
rect 6930 7884 6948 7902
rect 6930 7902 6948 7920
rect 6930 7920 6948 7938
rect 6930 7938 6948 7956
rect 6930 7956 6948 7974
rect 6930 7974 6948 7992
rect 6930 7992 6948 8010
rect 6930 8010 6948 8028
rect 6930 8028 6948 8046
rect 6930 8046 6948 8064
rect 6930 8064 6948 8082
rect 6930 8082 6948 8100
rect 6930 8100 6948 8118
rect 6930 8118 6948 8136
rect 6930 8136 6948 8154
rect 6930 8154 6948 8172
rect 6930 8172 6948 8190
rect 6930 8190 6948 8208
rect 6930 8208 6948 8226
rect 6930 8226 6948 8244
rect 6930 8244 6948 8262
rect 6930 8262 6948 8280
rect 6930 8280 6948 8298
rect 6930 8298 6948 8316
rect 6930 8316 6948 8334
rect 6930 8334 6948 8352
rect 6930 8352 6948 8370
rect 6930 8370 6948 8388
rect 6930 8388 6948 8406
rect 6930 8406 6948 8424
rect 6930 8424 6948 8442
rect 6930 8442 6948 8460
rect 6930 8460 6948 8478
rect 6930 8478 6948 8496
rect 6930 8496 6948 8514
rect 6930 8514 6948 8532
rect 6930 8532 6948 8550
rect 6930 8550 6948 8568
rect 6930 8568 6948 8586
rect 6930 8586 6948 8604
rect 6930 8604 6948 8622
rect 6930 8622 6948 8640
rect 6930 8640 6948 8658
rect 6930 8658 6948 8676
rect 6930 8676 6948 8694
rect 6930 8694 6948 8712
rect 6930 8712 6948 8730
rect 6930 8730 6948 8748
rect 6930 8748 6948 8766
rect 6930 8766 6948 8784
rect 6930 8784 6948 8802
rect 6930 8802 6948 8820
rect 6930 8820 6948 8838
rect 6930 8838 6948 8856
rect 6930 8856 6948 8874
rect 6930 8874 6948 8892
rect 6930 8892 6948 8910
rect 6930 8910 6948 8928
rect 6930 8928 6948 8946
rect 6930 8946 6948 8964
rect 6930 8964 6948 8982
rect 6930 8982 6948 9000
rect 6930 9000 6948 9018
rect 6930 9018 6948 9036
rect 6930 9036 6948 9054
rect 6930 9054 6948 9072
rect 6930 9072 6948 9090
rect 6930 9090 6948 9108
rect 6930 9108 6948 9126
rect 6930 9126 6948 9144
rect 6930 9144 6948 9162
rect 6930 9162 6948 9180
rect 6930 9180 6948 9198
rect 6930 9198 6948 9216
rect 6930 9216 6948 9234
rect 6930 9234 6948 9252
rect 6930 9252 6948 9270
rect 6930 9270 6948 9288
rect 6930 9288 6948 9306
rect 6930 9306 6948 9324
rect 6930 9324 6948 9342
rect 6930 9342 6948 9360
rect 6930 9360 6948 9378
rect 6930 9378 6948 9396
rect 6930 9396 6948 9414
rect 6930 9414 6948 9432
rect 6930 9432 6948 9450
rect 6930 9450 6948 9468
rect 6930 9468 6948 9486
rect 6930 9486 6948 9504
rect 6930 9504 6948 9522
rect 6930 9522 6948 9540
rect 6930 9540 6948 9558
rect 6930 9558 6948 9576
rect 6930 9576 6948 9594
rect 6930 9594 6948 9612
rect 6930 9612 6948 9630
rect 6930 9630 6948 9648
rect 6930 9648 6948 9666
rect 6930 9666 6948 9684
rect 6930 9684 6948 9702
rect 6930 9702 6948 9720
rect 6930 9720 6948 9738
rect 6930 9738 6948 9756
rect 6930 9756 6948 9774
rect 6930 9774 6948 9792
rect 6930 9792 6948 9810
rect 6930 9810 6948 9828
rect 6930 9828 6948 9846
rect 6930 9846 6948 9864
rect 6930 9864 6948 9882
rect 6930 9882 6948 9900
rect 6930 9900 6948 9918
rect 6930 9918 6948 9936
rect 6930 9936 6948 9954
rect 6930 9954 6948 9972
rect 6930 9972 6948 9990
rect 6930 9990 6948 10008
rect 6930 10008 6948 10026
rect 6930 10026 6948 10044
rect 6930 10044 6948 10062
rect 6930 10062 6948 10080
rect 6930 10080 6948 10098
rect 6930 10098 6948 10116
rect 6930 10116 6948 10134
rect 6930 10134 6948 10152
rect 6930 10152 6948 10170
rect 6930 10170 6948 10188
rect 6930 10188 6948 10206
rect 6930 10206 6948 10224
rect 6930 10224 6948 10242
rect 6930 10242 6948 10260
rect 6930 10260 6948 10278
rect 6930 10278 6948 10296
rect 6930 10296 6948 10314
rect 6930 10314 6948 10332
rect 6930 10332 6948 10350
rect 6930 10350 6948 10368
rect 6930 10368 6948 10386
rect 6930 10386 6948 10404
rect 6948 1764 6966 1782
rect 6948 1782 6966 1800
rect 6948 1800 6966 1818
rect 6948 1818 6966 1836
rect 6948 1836 6966 1854
rect 6948 1854 6966 1872
rect 6948 1872 6966 1890
rect 6948 1890 6966 1908
rect 6948 1908 6966 1926
rect 6948 1926 6966 1944
rect 6948 1944 6966 1962
rect 6948 1962 6966 1980
rect 6948 1980 6966 1998
rect 6948 1998 6966 2016
rect 6948 2016 6966 2034
rect 6948 2034 6966 2052
rect 6948 2052 6966 2070
rect 6948 2070 6966 2088
rect 6948 2088 6966 2106
rect 6948 2106 6966 2124
rect 6948 2124 6966 2142
rect 6948 2142 6966 2160
rect 6948 2160 6966 2178
rect 6948 2178 6966 2196
rect 6948 2196 6966 2214
rect 6948 2214 6966 2232
rect 6948 2232 6966 2250
rect 6948 2250 6966 2268
rect 6948 2268 6966 2286
rect 6948 2286 6966 2304
rect 6948 2304 6966 2322
rect 6948 2322 6966 2340
rect 6948 2340 6966 2358
rect 6948 2358 6966 2376
rect 6948 2376 6966 2394
rect 6948 2394 6966 2412
rect 6948 2412 6966 2430
rect 6948 2430 6966 2448
rect 6948 2448 6966 2466
rect 6948 2466 6966 2484
rect 6948 2484 6966 2502
rect 6948 2502 6966 2520
rect 6948 2520 6966 2538
rect 6948 2538 6966 2556
rect 6948 2556 6966 2574
rect 6948 2574 6966 2592
rect 6948 2592 6966 2610
rect 6948 2610 6966 2628
rect 6948 2628 6966 2646
rect 6948 2646 6966 2664
rect 6948 2664 6966 2682
rect 6948 2682 6966 2700
rect 6948 2700 6966 2718
rect 6948 2718 6966 2736
rect 6948 2736 6966 2754
rect 6948 2754 6966 2772
rect 6948 2772 6966 2790
rect 6948 2790 6966 2808
rect 6948 2808 6966 2826
rect 6948 2826 6966 2844
rect 6948 2844 6966 2862
rect 6948 2862 6966 2880
rect 6948 2880 6966 2898
rect 6948 2898 6966 2916
rect 6948 2916 6966 2934
rect 6948 2934 6966 2952
rect 6948 2952 6966 2970
rect 6948 2970 6966 2988
rect 6948 2988 6966 3006
rect 6948 3006 6966 3024
rect 6948 3024 6966 3042
rect 6948 3042 6966 3060
rect 6948 3060 6966 3078
rect 6948 3258 6966 3276
rect 6948 3276 6966 3294
rect 6948 3294 6966 3312
rect 6948 3312 6966 3330
rect 6948 3330 6966 3348
rect 6948 3348 6966 3366
rect 6948 3366 6966 3384
rect 6948 3384 6966 3402
rect 6948 3402 6966 3420
rect 6948 3420 6966 3438
rect 6948 3438 6966 3456
rect 6948 3456 6966 3474
rect 6948 3474 6966 3492
rect 6948 3492 6966 3510
rect 6948 3510 6966 3528
rect 6948 3528 6966 3546
rect 6948 3546 6966 3564
rect 6948 3564 6966 3582
rect 6948 3582 6966 3600
rect 6948 3600 6966 3618
rect 6948 3618 6966 3636
rect 6948 3636 6966 3654
rect 6948 3654 6966 3672
rect 6948 3672 6966 3690
rect 6948 3690 6966 3708
rect 6948 3708 6966 3726
rect 6948 3726 6966 3744
rect 6948 3744 6966 3762
rect 6948 3960 6966 3978
rect 6948 3978 6966 3996
rect 6948 3996 6966 4014
rect 6948 4014 6966 4032
rect 6948 4032 6966 4050
rect 6948 4050 6966 4068
rect 6948 4068 6966 4086
rect 6948 4086 6966 4104
rect 6948 4104 6966 4122
rect 6948 4122 6966 4140
rect 6948 4140 6966 4158
rect 6948 4158 6966 4176
rect 6948 4176 6966 4194
rect 6948 4194 6966 4212
rect 6948 4212 6966 4230
rect 6948 4230 6966 4248
rect 6948 4248 6966 4266
rect 6948 4266 6966 4284
rect 6948 4284 6966 4302
rect 6948 4302 6966 4320
rect 6948 4320 6966 4338
rect 6948 4338 6966 4356
rect 6948 4356 6966 4374
rect 6948 4374 6966 4392
rect 6948 4392 6966 4410
rect 6948 4410 6966 4428
rect 6948 4428 6966 4446
rect 6948 4446 6966 4464
rect 6948 4464 6966 4482
rect 6948 4482 6966 4500
rect 6948 4500 6966 4518
rect 6948 4518 6966 4536
rect 6948 4536 6966 4554
rect 6948 4554 6966 4572
rect 6948 4572 6966 4590
rect 6948 4590 6966 4608
rect 6948 4608 6966 4626
rect 6948 4626 6966 4644
rect 6948 4644 6966 4662
rect 6948 4662 6966 4680
rect 6948 4680 6966 4698
rect 6948 4698 6966 4716
rect 6948 4716 6966 4734
rect 6948 4734 6966 4752
rect 6948 4752 6966 4770
rect 6948 4770 6966 4788
rect 6948 4788 6966 4806
rect 6948 4806 6966 4824
rect 6948 4824 6966 4842
rect 6948 4842 6966 4860
rect 6948 4860 6966 4878
rect 6948 4878 6966 4896
rect 6948 4896 6966 4914
rect 6948 4914 6966 4932
rect 6948 4932 6966 4950
rect 6948 4950 6966 4968
rect 6948 4968 6966 4986
rect 6948 4986 6966 5004
rect 6948 5004 6966 5022
rect 6948 5022 6966 5040
rect 6948 5040 6966 5058
rect 6948 5058 6966 5076
rect 6948 5076 6966 5094
rect 6948 5094 6966 5112
rect 6948 5112 6966 5130
rect 6948 5130 6966 5148
rect 6948 5148 6966 5166
rect 6948 5166 6966 5184
rect 6948 5184 6966 5202
rect 6948 5202 6966 5220
rect 6948 5220 6966 5238
rect 6948 5238 6966 5256
rect 6948 5256 6966 5274
rect 6948 5274 6966 5292
rect 6948 5292 6966 5310
rect 6948 5310 6966 5328
rect 6948 5328 6966 5346
rect 6948 5346 6966 5364
rect 6948 5364 6966 5382
rect 6948 5382 6966 5400
rect 6948 5400 6966 5418
rect 6948 5418 6966 5436
rect 6948 5436 6966 5454
rect 6948 5454 6966 5472
rect 6948 5472 6966 5490
rect 6948 5490 6966 5508
rect 6948 5508 6966 5526
rect 6948 5526 6966 5544
rect 6948 5544 6966 5562
rect 6948 5562 6966 5580
rect 6948 5580 6966 5598
rect 6948 5598 6966 5616
rect 6948 5616 6966 5634
rect 6948 5634 6966 5652
rect 6948 5652 6966 5670
rect 6948 5670 6966 5688
rect 6948 5688 6966 5706
rect 6948 5706 6966 5724
rect 6948 5724 6966 5742
rect 6948 5742 6966 5760
rect 6948 5760 6966 5778
rect 6948 5778 6966 5796
rect 6948 5796 6966 5814
rect 6948 5814 6966 5832
rect 6948 5832 6966 5850
rect 6948 5850 6966 5868
rect 6948 5868 6966 5886
rect 6948 5886 6966 5904
rect 6948 5904 6966 5922
rect 6948 5922 6966 5940
rect 6948 5940 6966 5958
rect 6948 5958 6966 5976
rect 6948 5976 6966 5994
rect 6948 5994 6966 6012
rect 6948 6012 6966 6030
rect 6948 6030 6966 6048
rect 6948 6048 6966 6066
rect 6948 6066 6966 6084
rect 6948 6084 6966 6102
rect 6948 6102 6966 6120
rect 6948 6120 6966 6138
rect 6948 6138 6966 6156
rect 6948 6156 6966 6174
rect 6948 6174 6966 6192
rect 6948 6192 6966 6210
rect 6948 6210 6966 6228
rect 6948 7722 6966 7740
rect 6948 7740 6966 7758
rect 6948 7758 6966 7776
rect 6948 7776 6966 7794
rect 6948 7794 6966 7812
rect 6948 7812 6966 7830
rect 6948 7830 6966 7848
rect 6948 7848 6966 7866
rect 6948 7866 6966 7884
rect 6948 7884 6966 7902
rect 6948 7902 6966 7920
rect 6948 7920 6966 7938
rect 6948 7938 6966 7956
rect 6948 7956 6966 7974
rect 6948 7974 6966 7992
rect 6948 7992 6966 8010
rect 6948 8010 6966 8028
rect 6948 8028 6966 8046
rect 6948 8046 6966 8064
rect 6948 8064 6966 8082
rect 6948 8082 6966 8100
rect 6948 8100 6966 8118
rect 6948 8118 6966 8136
rect 6948 8136 6966 8154
rect 6948 8154 6966 8172
rect 6948 8172 6966 8190
rect 6948 8190 6966 8208
rect 6948 8208 6966 8226
rect 6948 8226 6966 8244
rect 6948 8244 6966 8262
rect 6948 8262 6966 8280
rect 6948 8280 6966 8298
rect 6948 8298 6966 8316
rect 6948 8316 6966 8334
rect 6948 8334 6966 8352
rect 6948 8352 6966 8370
rect 6948 8370 6966 8388
rect 6948 8388 6966 8406
rect 6948 8406 6966 8424
rect 6948 8424 6966 8442
rect 6948 8442 6966 8460
rect 6948 8460 6966 8478
rect 6948 8478 6966 8496
rect 6948 8496 6966 8514
rect 6948 8514 6966 8532
rect 6948 8532 6966 8550
rect 6948 8550 6966 8568
rect 6948 8568 6966 8586
rect 6948 8586 6966 8604
rect 6948 8604 6966 8622
rect 6948 8622 6966 8640
rect 6948 8640 6966 8658
rect 6948 8658 6966 8676
rect 6948 8676 6966 8694
rect 6948 8694 6966 8712
rect 6948 8712 6966 8730
rect 6948 8730 6966 8748
rect 6948 8748 6966 8766
rect 6948 8766 6966 8784
rect 6948 8784 6966 8802
rect 6948 8802 6966 8820
rect 6948 8820 6966 8838
rect 6948 8838 6966 8856
rect 6948 8856 6966 8874
rect 6948 8874 6966 8892
rect 6948 8892 6966 8910
rect 6948 8910 6966 8928
rect 6948 8928 6966 8946
rect 6948 8946 6966 8964
rect 6948 8964 6966 8982
rect 6948 8982 6966 9000
rect 6948 9000 6966 9018
rect 6948 9018 6966 9036
rect 6948 9036 6966 9054
rect 6948 9054 6966 9072
rect 6948 9072 6966 9090
rect 6948 9090 6966 9108
rect 6948 9108 6966 9126
rect 6948 9126 6966 9144
rect 6948 9144 6966 9162
rect 6948 9162 6966 9180
rect 6948 9180 6966 9198
rect 6948 9198 6966 9216
rect 6948 9216 6966 9234
rect 6948 9234 6966 9252
rect 6948 9252 6966 9270
rect 6948 9270 6966 9288
rect 6948 9288 6966 9306
rect 6948 9306 6966 9324
rect 6948 9324 6966 9342
rect 6948 9342 6966 9360
rect 6948 9360 6966 9378
rect 6948 9378 6966 9396
rect 6948 9396 6966 9414
rect 6948 9414 6966 9432
rect 6948 9432 6966 9450
rect 6948 9450 6966 9468
rect 6948 9468 6966 9486
rect 6948 9486 6966 9504
rect 6948 9504 6966 9522
rect 6948 9522 6966 9540
rect 6948 9540 6966 9558
rect 6948 9558 6966 9576
rect 6948 9576 6966 9594
rect 6948 9594 6966 9612
rect 6948 9612 6966 9630
rect 6948 9630 6966 9648
rect 6948 9648 6966 9666
rect 6948 9666 6966 9684
rect 6948 9684 6966 9702
rect 6948 9702 6966 9720
rect 6948 9720 6966 9738
rect 6948 9738 6966 9756
rect 6948 9756 6966 9774
rect 6948 9774 6966 9792
rect 6948 9792 6966 9810
rect 6948 9810 6966 9828
rect 6948 9828 6966 9846
rect 6948 9846 6966 9864
rect 6948 9864 6966 9882
rect 6948 9882 6966 9900
rect 6948 9900 6966 9918
rect 6948 9918 6966 9936
rect 6948 9936 6966 9954
rect 6948 9954 6966 9972
rect 6948 9972 6966 9990
rect 6948 9990 6966 10008
rect 6948 10008 6966 10026
rect 6948 10026 6966 10044
rect 6948 10044 6966 10062
rect 6948 10062 6966 10080
rect 6948 10080 6966 10098
rect 6948 10098 6966 10116
rect 6948 10116 6966 10134
rect 6948 10134 6966 10152
rect 6948 10152 6966 10170
rect 6948 10170 6966 10188
rect 6948 10188 6966 10206
rect 6948 10206 6966 10224
rect 6948 10224 6966 10242
rect 6948 10242 6966 10260
rect 6948 10260 6966 10278
rect 6948 10278 6966 10296
rect 6948 10296 6966 10314
rect 6948 10314 6966 10332
rect 6948 10332 6966 10350
rect 6948 10350 6966 10368
rect 6948 10368 6966 10386
rect 6948 10386 6966 10404
rect 6948 10404 6966 10422
rect 6966 1764 6984 1782
rect 6966 1782 6984 1800
rect 6966 1800 6984 1818
rect 6966 1818 6984 1836
rect 6966 1836 6984 1854
rect 6966 1854 6984 1872
rect 6966 1872 6984 1890
rect 6966 1890 6984 1908
rect 6966 1908 6984 1926
rect 6966 1926 6984 1944
rect 6966 1944 6984 1962
rect 6966 1962 6984 1980
rect 6966 1980 6984 1998
rect 6966 1998 6984 2016
rect 6966 2016 6984 2034
rect 6966 2034 6984 2052
rect 6966 2052 6984 2070
rect 6966 2070 6984 2088
rect 6966 2088 6984 2106
rect 6966 2106 6984 2124
rect 6966 2124 6984 2142
rect 6966 2142 6984 2160
rect 6966 2160 6984 2178
rect 6966 2178 6984 2196
rect 6966 2196 6984 2214
rect 6966 2214 6984 2232
rect 6966 2232 6984 2250
rect 6966 2250 6984 2268
rect 6966 2268 6984 2286
rect 6966 2286 6984 2304
rect 6966 2304 6984 2322
rect 6966 2322 6984 2340
rect 6966 2340 6984 2358
rect 6966 2358 6984 2376
rect 6966 2376 6984 2394
rect 6966 2394 6984 2412
rect 6966 2412 6984 2430
rect 6966 2430 6984 2448
rect 6966 2448 6984 2466
rect 6966 2466 6984 2484
rect 6966 2484 6984 2502
rect 6966 2502 6984 2520
rect 6966 2520 6984 2538
rect 6966 2538 6984 2556
rect 6966 2556 6984 2574
rect 6966 2574 6984 2592
rect 6966 2592 6984 2610
rect 6966 2610 6984 2628
rect 6966 2628 6984 2646
rect 6966 2646 6984 2664
rect 6966 2664 6984 2682
rect 6966 2682 6984 2700
rect 6966 2700 6984 2718
rect 6966 2718 6984 2736
rect 6966 2736 6984 2754
rect 6966 2754 6984 2772
rect 6966 2772 6984 2790
rect 6966 2790 6984 2808
rect 6966 2808 6984 2826
rect 6966 2826 6984 2844
rect 6966 2844 6984 2862
rect 6966 2862 6984 2880
rect 6966 2880 6984 2898
rect 6966 2898 6984 2916
rect 6966 2916 6984 2934
rect 6966 2934 6984 2952
rect 6966 2952 6984 2970
rect 6966 2970 6984 2988
rect 6966 2988 6984 3006
rect 6966 3006 6984 3024
rect 6966 3024 6984 3042
rect 6966 3042 6984 3060
rect 6966 3060 6984 3078
rect 6966 3258 6984 3276
rect 6966 3276 6984 3294
rect 6966 3294 6984 3312
rect 6966 3312 6984 3330
rect 6966 3330 6984 3348
rect 6966 3348 6984 3366
rect 6966 3366 6984 3384
rect 6966 3384 6984 3402
rect 6966 3402 6984 3420
rect 6966 3420 6984 3438
rect 6966 3438 6984 3456
rect 6966 3456 6984 3474
rect 6966 3474 6984 3492
rect 6966 3492 6984 3510
rect 6966 3510 6984 3528
rect 6966 3528 6984 3546
rect 6966 3546 6984 3564
rect 6966 3564 6984 3582
rect 6966 3582 6984 3600
rect 6966 3600 6984 3618
rect 6966 3618 6984 3636
rect 6966 3636 6984 3654
rect 6966 3654 6984 3672
rect 6966 3672 6984 3690
rect 6966 3690 6984 3708
rect 6966 3708 6984 3726
rect 6966 3726 6984 3744
rect 6966 3744 6984 3762
rect 6966 3762 6984 3780
rect 6966 3978 6984 3996
rect 6966 3996 6984 4014
rect 6966 4014 6984 4032
rect 6966 4032 6984 4050
rect 6966 4050 6984 4068
rect 6966 4068 6984 4086
rect 6966 4086 6984 4104
rect 6966 4104 6984 4122
rect 6966 4122 6984 4140
rect 6966 4140 6984 4158
rect 6966 4158 6984 4176
rect 6966 4176 6984 4194
rect 6966 4194 6984 4212
rect 6966 4212 6984 4230
rect 6966 4230 6984 4248
rect 6966 4248 6984 4266
rect 6966 4266 6984 4284
rect 6966 4284 6984 4302
rect 6966 4302 6984 4320
rect 6966 4320 6984 4338
rect 6966 4338 6984 4356
rect 6966 4356 6984 4374
rect 6966 4374 6984 4392
rect 6966 4392 6984 4410
rect 6966 4410 6984 4428
rect 6966 4428 6984 4446
rect 6966 4446 6984 4464
rect 6966 4464 6984 4482
rect 6966 4482 6984 4500
rect 6966 4500 6984 4518
rect 6966 4518 6984 4536
rect 6966 4536 6984 4554
rect 6966 4554 6984 4572
rect 6966 4572 6984 4590
rect 6966 4590 6984 4608
rect 6966 4608 6984 4626
rect 6966 4626 6984 4644
rect 6966 4644 6984 4662
rect 6966 4662 6984 4680
rect 6966 4680 6984 4698
rect 6966 4698 6984 4716
rect 6966 4716 6984 4734
rect 6966 4734 6984 4752
rect 6966 4752 6984 4770
rect 6966 4770 6984 4788
rect 6966 4788 6984 4806
rect 6966 4806 6984 4824
rect 6966 4824 6984 4842
rect 6966 4842 6984 4860
rect 6966 4860 6984 4878
rect 6966 4878 6984 4896
rect 6966 4896 6984 4914
rect 6966 4914 6984 4932
rect 6966 4932 6984 4950
rect 6966 4950 6984 4968
rect 6966 4968 6984 4986
rect 6966 4986 6984 5004
rect 6966 5004 6984 5022
rect 6966 5022 6984 5040
rect 6966 5040 6984 5058
rect 6966 5058 6984 5076
rect 6966 5076 6984 5094
rect 6966 5094 6984 5112
rect 6966 5112 6984 5130
rect 6966 5130 6984 5148
rect 6966 5148 6984 5166
rect 6966 5166 6984 5184
rect 6966 5184 6984 5202
rect 6966 5202 6984 5220
rect 6966 5220 6984 5238
rect 6966 5238 6984 5256
rect 6966 5256 6984 5274
rect 6966 5274 6984 5292
rect 6966 5292 6984 5310
rect 6966 5310 6984 5328
rect 6966 5328 6984 5346
rect 6966 5346 6984 5364
rect 6966 5364 6984 5382
rect 6966 5382 6984 5400
rect 6966 5400 6984 5418
rect 6966 5418 6984 5436
rect 6966 5436 6984 5454
rect 6966 5454 6984 5472
rect 6966 5472 6984 5490
rect 6966 5490 6984 5508
rect 6966 5508 6984 5526
rect 6966 5526 6984 5544
rect 6966 5544 6984 5562
rect 6966 5562 6984 5580
rect 6966 5580 6984 5598
rect 6966 5598 6984 5616
rect 6966 5616 6984 5634
rect 6966 5634 6984 5652
rect 6966 5652 6984 5670
rect 6966 5670 6984 5688
rect 6966 5688 6984 5706
rect 6966 5706 6984 5724
rect 6966 5724 6984 5742
rect 6966 5742 6984 5760
rect 6966 5760 6984 5778
rect 6966 5778 6984 5796
rect 6966 5796 6984 5814
rect 6966 5814 6984 5832
rect 6966 5832 6984 5850
rect 6966 5850 6984 5868
rect 6966 5868 6984 5886
rect 6966 5886 6984 5904
rect 6966 5904 6984 5922
rect 6966 5922 6984 5940
rect 6966 5940 6984 5958
rect 6966 5958 6984 5976
rect 6966 5976 6984 5994
rect 6966 5994 6984 6012
rect 6966 6012 6984 6030
rect 6966 6030 6984 6048
rect 6966 6048 6984 6066
rect 6966 6066 6984 6084
rect 6966 6084 6984 6102
rect 6966 6102 6984 6120
rect 6966 6120 6984 6138
rect 6966 6138 6984 6156
rect 6966 6156 6984 6174
rect 6966 6174 6984 6192
rect 6966 6192 6984 6210
rect 6966 6210 6984 6228
rect 6966 7776 6984 7794
rect 6966 7794 6984 7812
rect 6966 7812 6984 7830
rect 6966 7830 6984 7848
rect 6966 7848 6984 7866
rect 6966 7866 6984 7884
rect 6966 7884 6984 7902
rect 6966 7902 6984 7920
rect 6966 7920 6984 7938
rect 6966 7938 6984 7956
rect 6966 7956 6984 7974
rect 6966 7974 6984 7992
rect 6966 7992 6984 8010
rect 6966 8010 6984 8028
rect 6966 8028 6984 8046
rect 6966 8046 6984 8064
rect 6966 8064 6984 8082
rect 6966 8082 6984 8100
rect 6966 8100 6984 8118
rect 6966 8118 6984 8136
rect 6966 8136 6984 8154
rect 6966 8154 6984 8172
rect 6966 8172 6984 8190
rect 6966 8190 6984 8208
rect 6966 8208 6984 8226
rect 6966 8226 6984 8244
rect 6966 8244 6984 8262
rect 6966 8262 6984 8280
rect 6966 8280 6984 8298
rect 6966 8298 6984 8316
rect 6966 8316 6984 8334
rect 6966 8334 6984 8352
rect 6966 8352 6984 8370
rect 6966 8370 6984 8388
rect 6966 8388 6984 8406
rect 6966 8406 6984 8424
rect 6966 8424 6984 8442
rect 6966 8442 6984 8460
rect 6966 8460 6984 8478
rect 6966 8478 6984 8496
rect 6966 8496 6984 8514
rect 6966 8514 6984 8532
rect 6966 8532 6984 8550
rect 6966 8550 6984 8568
rect 6966 8568 6984 8586
rect 6966 8586 6984 8604
rect 6966 8604 6984 8622
rect 6966 8622 6984 8640
rect 6966 8640 6984 8658
rect 6966 8658 6984 8676
rect 6966 8676 6984 8694
rect 6966 8694 6984 8712
rect 6966 8712 6984 8730
rect 6966 8730 6984 8748
rect 6966 8748 6984 8766
rect 6966 8766 6984 8784
rect 6966 8784 6984 8802
rect 6966 8802 6984 8820
rect 6966 8820 6984 8838
rect 6966 8838 6984 8856
rect 6966 8856 6984 8874
rect 6966 8874 6984 8892
rect 6966 8892 6984 8910
rect 6966 8910 6984 8928
rect 6966 8928 6984 8946
rect 6966 8946 6984 8964
rect 6966 8964 6984 8982
rect 6966 8982 6984 9000
rect 6966 9000 6984 9018
rect 6966 9018 6984 9036
rect 6966 9036 6984 9054
rect 6966 9054 6984 9072
rect 6966 9072 6984 9090
rect 6966 9090 6984 9108
rect 6966 9108 6984 9126
rect 6966 9126 6984 9144
rect 6966 9144 6984 9162
rect 6966 9162 6984 9180
rect 6966 9180 6984 9198
rect 6966 9198 6984 9216
rect 6966 9216 6984 9234
rect 6966 9234 6984 9252
rect 6966 9252 6984 9270
rect 6966 9270 6984 9288
rect 6966 9288 6984 9306
rect 6966 9306 6984 9324
rect 6966 9324 6984 9342
rect 6966 9342 6984 9360
rect 6966 9360 6984 9378
rect 6966 9378 6984 9396
rect 6966 9396 6984 9414
rect 6966 9414 6984 9432
rect 6966 9432 6984 9450
rect 6966 9450 6984 9468
rect 6966 9468 6984 9486
rect 6966 9486 6984 9504
rect 6966 9504 6984 9522
rect 6966 9522 6984 9540
rect 6966 9540 6984 9558
rect 6966 9558 6984 9576
rect 6966 9576 6984 9594
rect 6966 9594 6984 9612
rect 6966 9612 6984 9630
rect 6966 9630 6984 9648
rect 6966 9648 6984 9666
rect 6966 9666 6984 9684
rect 6966 9684 6984 9702
rect 6966 9702 6984 9720
rect 6966 9720 6984 9738
rect 6966 9738 6984 9756
rect 6966 9756 6984 9774
rect 6966 9774 6984 9792
rect 6966 9792 6984 9810
rect 6966 9810 6984 9828
rect 6966 9828 6984 9846
rect 6966 9846 6984 9864
rect 6966 9864 6984 9882
rect 6966 9882 6984 9900
rect 6966 9900 6984 9918
rect 6966 9918 6984 9936
rect 6966 9936 6984 9954
rect 6966 9954 6984 9972
rect 6966 9972 6984 9990
rect 6966 9990 6984 10008
rect 6966 10008 6984 10026
rect 6966 10026 6984 10044
rect 6966 10044 6984 10062
rect 6966 10062 6984 10080
rect 6966 10080 6984 10098
rect 6966 10098 6984 10116
rect 6966 10116 6984 10134
rect 6966 10134 6984 10152
rect 6966 10152 6984 10170
rect 6966 10170 6984 10188
rect 6966 10188 6984 10206
rect 6966 10206 6984 10224
rect 6966 10224 6984 10242
rect 6966 10242 6984 10260
rect 6966 10260 6984 10278
rect 6966 10278 6984 10296
rect 6966 10296 6984 10314
rect 6966 10314 6984 10332
rect 6966 10332 6984 10350
rect 6966 10350 6984 10368
rect 6966 10368 6984 10386
rect 6966 10386 6984 10404
rect 6966 10404 6984 10422
rect 6966 10422 6984 10440
rect 6984 1782 7002 1800
rect 6984 1800 7002 1818
rect 6984 1818 7002 1836
rect 6984 1836 7002 1854
rect 6984 1854 7002 1872
rect 6984 1872 7002 1890
rect 6984 1890 7002 1908
rect 6984 1908 7002 1926
rect 6984 1926 7002 1944
rect 6984 1944 7002 1962
rect 6984 1962 7002 1980
rect 6984 1980 7002 1998
rect 6984 1998 7002 2016
rect 6984 2016 7002 2034
rect 6984 2034 7002 2052
rect 6984 2052 7002 2070
rect 6984 2070 7002 2088
rect 6984 2088 7002 2106
rect 6984 2106 7002 2124
rect 6984 2124 7002 2142
rect 6984 2142 7002 2160
rect 6984 2160 7002 2178
rect 6984 2178 7002 2196
rect 6984 2196 7002 2214
rect 6984 2214 7002 2232
rect 6984 2232 7002 2250
rect 6984 2250 7002 2268
rect 6984 2268 7002 2286
rect 6984 2286 7002 2304
rect 6984 2304 7002 2322
rect 6984 2322 7002 2340
rect 6984 2340 7002 2358
rect 6984 2358 7002 2376
rect 6984 2376 7002 2394
rect 6984 2394 7002 2412
rect 6984 2412 7002 2430
rect 6984 2430 7002 2448
rect 6984 2448 7002 2466
rect 6984 2466 7002 2484
rect 6984 2484 7002 2502
rect 6984 2502 7002 2520
rect 6984 2520 7002 2538
rect 6984 2538 7002 2556
rect 6984 2556 7002 2574
rect 6984 2574 7002 2592
rect 6984 2592 7002 2610
rect 6984 2610 7002 2628
rect 6984 2628 7002 2646
rect 6984 2646 7002 2664
rect 6984 2664 7002 2682
rect 6984 2682 7002 2700
rect 6984 2700 7002 2718
rect 6984 2718 7002 2736
rect 6984 2736 7002 2754
rect 6984 2754 7002 2772
rect 6984 2772 7002 2790
rect 6984 2790 7002 2808
rect 6984 2808 7002 2826
rect 6984 2826 7002 2844
rect 6984 2844 7002 2862
rect 6984 2862 7002 2880
rect 6984 2880 7002 2898
rect 6984 2898 7002 2916
rect 6984 2916 7002 2934
rect 6984 2934 7002 2952
rect 6984 2952 7002 2970
rect 6984 2970 7002 2988
rect 6984 2988 7002 3006
rect 6984 3006 7002 3024
rect 6984 3024 7002 3042
rect 6984 3042 7002 3060
rect 6984 3060 7002 3078
rect 6984 3078 7002 3096
rect 6984 3258 7002 3276
rect 6984 3276 7002 3294
rect 6984 3294 7002 3312
rect 6984 3312 7002 3330
rect 6984 3330 7002 3348
rect 6984 3348 7002 3366
rect 6984 3366 7002 3384
rect 6984 3384 7002 3402
rect 6984 3402 7002 3420
rect 6984 3420 7002 3438
rect 6984 3438 7002 3456
rect 6984 3456 7002 3474
rect 6984 3474 7002 3492
rect 6984 3492 7002 3510
rect 6984 3510 7002 3528
rect 6984 3528 7002 3546
rect 6984 3546 7002 3564
rect 6984 3564 7002 3582
rect 6984 3582 7002 3600
rect 6984 3600 7002 3618
rect 6984 3618 7002 3636
rect 6984 3636 7002 3654
rect 6984 3654 7002 3672
rect 6984 3672 7002 3690
rect 6984 3690 7002 3708
rect 6984 3708 7002 3726
rect 6984 3726 7002 3744
rect 6984 3744 7002 3762
rect 6984 3762 7002 3780
rect 6984 3780 7002 3798
rect 6984 4014 7002 4032
rect 6984 4032 7002 4050
rect 6984 4050 7002 4068
rect 6984 4068 7002 4086
rect 6984 4086 7002 4104
rect 6984 4104 7002 4122
rect 6984 4122 7002 4140
rect 6984 4140 7002 4158
rect 6984 4158 7002 4176
rect 6984 4176 7002 4194
rect 6984 4194 7002 4212
rect 6984 4212 7002 4230
rect 6984 4230 7002 4248
rect 6984 4248 7002 4266
rect 6984 4266 7002 4284
rect 6984 4284 7002 4302
rect 6984 4302 7002 4320
rect 6984 4320 7002 4338
rect 6984 4338 7002 4356
rect 6984 4356 7002 4374
rect 6984 4374 7002 4392
rect 6984 4392 7002 4410
rect 6984 4410 7002 4428
rect 6984 4428 7002 4446
rect 6984 4446 7002 4464
rect 6984 4464 7002 4482
rect 6984 4482 7002 4500
rect 6984 4500 7002 4518
rect 6984 4518 7002 4536
rect 6984 4536 7002 4554
rect 6984 4554 7002 4572
rect 6984 4572 7002 4590
rect 6984 4590 7002 4608
rect 6984 4608 7002 4626
rect 6984 4626 7002 4644
rect 6984 4644 7002 4662
rect 6984 4662 7002 4680
rect 6984 4680 7002 4698
rect 6984 4698 7002 4716
rect 6984 4716 7002 4734
rect 6984 4734 7002 4752
rect 6984 4752 7002 4770
rect 6984 4770 7002 4788
rect 6984 4788 7002 4806
rect 6984 4806 7002 4824
rect 6984 4824 7002 4842
rect 6984 4842 7002 4860
rect 6984 4860 7002 4878
rect 6984 4878 7002 4896
rect 6984 4896 7002 4914
rect 6984 4914 7002 4932
rect 6984 4932 7002 4950
rect 6984 4950 7002 4968
rect 6984 4968 7002 4986
rect 6984 4986 7002 5004
rect 6984 5004 7002 5022
rect 6984 5022 7002 5040
rect 6984 5040 7002 5058
rect 6984 5058 7002 5076
rect 6984 5076 7002 5094
rect 6984 5094 7002 5112
rect 6984 5112 7002 5130
rect 6984 5130 7002 5148
rect 6984 5148 7002 5166
rect 6984 5166 7002 5184
rect 6984 5184 7002 5202
rect 6984 5202 7002 5220
rect 6984 5220 7002 5238
rect 6984 5238 7002 5256
rect 6984 5256 7002 5274
rect 6984 5274 7002 5292
rect 6984 5292 7002 5310
rect 6984 5310 7002 5328
rect 6984 5328 7002 5346
rect 6984 5346 7002 5364
rect 6984 5364 7002 5382
rect 6984 5382 7002 5400
rect 6984 5400 7002 5418
rect 6984 5418 7002 5436
rect 6984 5436 7002 5454
rect 6984 5454 7002 5472
rect 6984 5472 7002 5490
rect 6984 5490 7002 5508
rect 6984 5508 7002 5526
rect 6984 5526 7002 5544
rect 6984 5544 7002 5562
rect 6984 5562 7002 5580
rect 6984 5580 7002 5598
rect 6984 5598 7002 5616
rect 6984 5616 7002 5634
rect 6984 5634 7002 5652
rect 6984 5652 7002 5670
rect 6984 5670 7002 5688
rect 6984 5688 7002 5706
rect 6984 5706 7002 5724
rect 6984 5724 7002 5742
rect 6984 5742 7002 5760
rect 6984 5760 7002 5778
rect 6984 5778 7002 5796
rect 6984 5796 7002 5814
rect 6984 5814 7002 5832
rect 6984 5832 7002 5850
rect 6984 5850 7002 5868
rect 6984 5868 7002 5886
rect 6984 5886 7002 5904
rect 6984 5904 7002 5922
rect 6984 5922 7002 5940
rect 6984 5940 7002 5958
rect 6984 5958 7002 5976
rect 6984 5976 7002 5994
rect 6984 5994 7002 6012
rect 6984 6012 7002 6030
rect 6984 6030 7002 6048
rect 6984 6048 7002 6066
rect 6984 6066 7002 6084
rect 6984 6084 7002 6102
rect 6984 6102 7002 6120
rect 6984 6120 7002 6138
rect 6984 6138 7002 6156
rect 6984 6156 7002 6174
rect 6984 6174 7002 6192
rect 6984 6192 7002 6210
rect 6984 6210 7002 6228
rect 6984 6228 7002 6246
rect 6984 7812 7002 7830
rect 6984 7830 7002 7848
rect 6984 7848 7002 7866
rect 6984 7866 7002 7884
rect 6984 7884 7002 7902
rect 6984 7902 7002 7920
rect 6984 7920 7002 7938
rect 6984 7938 7002 7956
rect 6984 7956 7002 7974
rect 6984 7974 7002 7992
rect 6984 7992 7002 8010
rect 6984 8010 7002 8028
rect 6984 8028 7002 8046
rect 6984 8046 7002 8064
rect 6984 8064 7002 8082
rect 6984 8082 7002 8100
rect 6984 8100 7002 8118
rect 6984 8118 7002 8136
rect 6984 8136 7002 8154
rect 6984 8154 7002 8172
rect 6984 8172 7002 8190
rect 6984 8190 7002 8208
rect 6984 8208 7002 8226
rect 6984 8226 7002 8244
rect 6984 8244 7002 8262
rect 6984 8262 7002 8280
rect 6984 8280 7002 8298
rect 6984 8298 7002 8316
rect 6984 8316 7002 8334
rect 6984 8334 7002 8352
rect 6984 8352 7002 8370
rect 6984 8370 7002 8388
rect 6984 8388 7002 8406
rect 6984 8406 7002 8424
rect 6984 8424 7002 8442
rect 6984 8442 7002 8460
rect 6984 8460 7002 8478
rect 6984 8478 7002 8496
rect 6984 8496 7002 8514
rect 6984 8514 7002 8532
rect 6984 8532 7002 8550
rect 6984 8550 7002 8568
rect 6984 8568 7002 8586
rect 6984 8586 7002 8604
rect 6984 8604 7002 8622
rect 6984 8622 7002 8640
rect 6984 8640 7002 8658
rect 6984 8658 7002 8676
rect 6984 8676 7002 8694
rect 6984 8694 7002 8712
rect 6984 8712 7002 8730
rect 6984 8730 7002 8748
rect 6984 8748 7002 8766
rect 6984 8766 7002 8784
rect 6984 8784 7002 8802
rect 6984 8802 7002 8820
rect 6984 8820 7002 8838
rect 6984 8838 7002 8856
rect 6984 8856 7002 8874
rect 6984 8874 7002 8892
rect 6984 8892 7002 8910
rect 6984 8910 7002 8928
rect 6984 8928 7002 8946
rect 6984 8946 7002 8964
rect 6984 8964 7002 8982
rect 6984 8982 7002 9000
rect 6984 9000 7002 9018
rect 6984 9018 7002 9036
rect 6984 9036 7002 9054
rect 6984 9054 7002 9072
rect 6984 9072 7002 9090
rect 6984 9090 7002 9108
rect 6984 9108 7002 9126
rect 6984 9126 7002 9144
rect 6984 9144 7002 9162
rect 6984 9162 7002 9180
rect 6984 9180 7002 9198
rect 6984 9198 7002 9216
rect 6984 9216 7002 9234
rect 6984 9234 7002 9252
rect 6984 9252 7002 9270
rect 6984 9270 7002 9288
rect 6984 9288 7002 9306
rect 6984 9306 7002 9324
rect 6984 9324 7002 9342
rect 6984 9342 7002 9360
rect 6984 9360 7002 9378
rect 6984 9378 7002 9396
rect 6984 9396 7002 9414
rect 6984 9414 7002 9432
rect 6984 9432 7002 9450
rect 6984 9450 7002 9468
rect 6984 9468 7002 9486
rect 6984 9486 7002 9504
rect 6984 9504 7002 9522
rect 6984 9522 7002 9540
rect 6984 9540 7002 9558
rect 6984 9558 7002 9576
rect 6984 9576 7002 9594
rect 6984 9594 7002 9612
rect 6984 9612 7002 9630
rect 6984 9630 7002 9648
rect 6984 9648 7002 9666
rect 6984 9666 7002 9684
rect 6984 9684 7002 9702
rect 6984 9702 7002 9720
rect 6984 9720 7002 9738
rect 6984 9738 7002 9756
rect 6984 9756 7002 9774
rect 6984 9774 7002 9792
rect 6984 9792 7002 9810
rect 6984 9810 7002 9828
rect 6984 9828 7002 9846
rect 6984 9846 7002 9864
rect 6984 9864 7002 9882
rect 6984 9882 7002 9900
rect 6984 9900 7002 9918
rect 6984 9918 7002 9936
rect 6984 9936 7002 9954
rect 6984 9954 7002 9972
rect 6984 9972 7002 9990
rect 6984 9990 7002 10008
rect 6984 10008 7002 10026
rect 6984 10026 7002 10044
rect 6984 10044 7002 10062
rect 6984 10062 7002 10080
rect 6984 10080 7002 10098
rect 6984 10098 7002 10116
rect 6984 10116 7002 10134
rect 6984 10134 7002 10152
rect 6984 10152 7002 10170
rect 6984 10170 7002 10188
rect 6984 10188 7002 10206
rect 6984 10206 7002 10224
rect 6984 10224 7002 10242
rect 6984 10242 7002 10260
rect 6984 10260 7002 10278
rect 6984 10278 7002 10296
rect 6984 10296 7002 10314
rect 6984 10314 7002 10332
rect 6984 10332 7002 10350
rect 6984 10350 7002 10368
rect 6984 10368 7002 10386
rect 6984 10386 7002 10404
rect 6984 10404 7002 10422
rect 6984 10422 7002 10440
rect 6984 10440 7002 10458
rect 7002 1782 7020 1800
rect 7002 1800 7020 1818
rect 7002 1818 7020 1836
rect 7002 1836 7020 1854
rect 7002 1854 7020 1872
rect 7002 1872 7020 1890
rect 7002 1890 7020 1908
rect 7002 1908 7020 1926
rect 7002 1926 7020 1944
rect 7002 1944 7020 1962
rect 7002 1962 7020 1980
rect 7002 1980 7020 1998
rect 7002 1998 7020 2016
rect 7002 2016 7020 2034
rect 7002 2034 7020 2052
rect 7002 2052 7020 2070
rect 7002 2070 7020 2088
rect 7002 2088 7020 2106
rect 7002 2106 7020 2124
rect 7002 2124 7020 2142
rect 7002 2142 7020 2160
rect 7002 2160 7020 2178
rect 7002 2178 7020 2196
rect 7002 2196 7020 2214
rect 7002 2214 7020 2232
rect 7002 2232 7020 2250
rect 7002 2250 7020 2268
rect 7002 2268 7020 2286
rect 7002 2286 7020 2304
rect 7002 2304 7020 2322
rect 7002 2322 7020 2340
rect 7002 2340 7020 2358
rect 7002 2358 7020 2376
rect 7002 2376 7020 2394
rect 7002 2394 7020 2412
rect 7002 2412 7020 2430
rect 7002 2430 7020 2448
rect 7002 2448 7020 2466
rect 7002 2466 7020 2484
rect 7002 2484 7020 2502
rect 7002 2502 7020 2520
rect 7002 2520 7020 2538
rect 7002 2538 7020 2556
rect 7002 2556 7020 2574
rect 7002 2574 7020 2592
rect 7002 2592 7020 2610
rect 7002 2610 7020 2628
rect 7002 2628 7020 2646
rect 7002 2646 7020 2664
rect 7002 2664 7020 2682
rect 7002 2682 7020 2700
rect 7002 2700 7020 2718
rect 7002 2718 7020 2736
rect 7002 2736 7020 2754
rect 7002 2754 7020 2772
rect 7002 2772 7020 2790
rect 7002 2790 7020 2808
rect 7002 2808 7020 2826
rect 7002 2826 7020 2844
rect 7002 2844 7020 2862
rect 7002 2862 7020 2880
rect 7002 2880 7020 2898
rect 7002 2898 7020 2916
rect 7002 2916 7020 2934
rect 7002 2934 7020 2952
rect 7002 2952 7020 2970
rect 7002 2970 7020 2988
rect 7002 2988 7020 3006
rect 7002 3006 7020 3024
rect 7002 3024 7020 3042
rect 7002 3042 7020 3060
rect 7002 3060 7020 3078
rect 7002 3078 7020 3096
rect 7002 3276 7020 3294
rect 7002 3294 7020 3312
rect 7002 3312 7020 3330
rect 7002 3330 7020 3348
rect 7002 3348 7020 3366
rect 7002 3366 7020 3384
rect 7002 3384 7020 3402
rect 7002 3402 7020 3420
rect 7002 3420 7020 3438
rect 7002 3438 7020 3456
rect 7002 3456 7020 3474
rect 7002 3474 7020 3492
rect 7002 3492 7020 3510
rect 7002 3510 7020 3528
rect 7002 3528 7020 3546
rect 7002 3546 7020 3564
rect 7002 3564 7020 3582
rect 7002 3582 7020 3600
rect 7002 3600 7020 3618
rect 7002 3618 7020 3636
rect 7002 3636 7020 3654
rect 7002 3654 7020 3672
rect 7002 3672 7020 3690
rect 7002 3690 7020 3708
rect 7002 3708 7020 3726
rect 7002 3726 7020 3744
rect 7002 3744 7020 3762
rect 7002 3762 7020 3780
rect 7002 3780 7020 3798
rect 7002 3798 7020 3816
rect 7002 4032 7020 4050
rect 7002 4050 7020 4068
rect 7002 4068 7020 4086
rect 7002 4086 7020 4104
rect 7002 4104 7020 4122
rect 7002 4122 7020 4140
rect 7002 4140 7020 4158
rect 7002 4158 7020 4176
rect 7002 4176 7020 4194
rect 7002 4194 7020 4212
rect 7002 4212 7020 4230
rect 7002 4230 7020 4248
rect 7002 4248 7020 4266
rect 7002 4266 7020 4284
rect 7002 4284 7020 4302
rect 7002 4302 7020 4320
rect 7002 4320 7020 4338
rect 7002 4338 7020 4356
rect 7002 4356 7020 4374
rect 7002 4374 7020 4392
rect 7002 4392 7020 4410
rect 7002 4410 7020 4428
rect 7002 4428 7020 4446
rect 7002 4446 7020 4464
rect 7002 4464 7020 4482
rect 7002 4482 7020 4500
rect 7002 4500 7020 4518
rect 7002 4518 7020 4536
rect 7002 4536 7020 4554
rect 7002 4554 7020 4572
rect 7002 4572 7020 4590
rect 7002 4590 7020 4608
rect 7002 4608 7020 4626
rect 7002 4626 7020 4644
rect 7002 4644 7020 4662
rect 7002 4662 7020 4680
rect 7002 4680 7020 4698
rect 7002 4698 7020 4716
rect 7002 4716 7020 4734
rect 7002 4734 7020 4752
rect 7002 4752 7020 4770
rect 7002 4770 7020 4788
rect 7002 4788 7020 4806
rect 7002 4806 7020 4824
rect 7002 4824 7020 4842
rect 7002 4842 7020 4860
rect 7002 4860 7020 4878
rect 7002 4878 7020 4896
rect 7002 4896 7020 4914
rect 7002 4914 7020 4932
rect 7002 4932 7020 4950
rect 7002 4950 7020 4968
rect 7002 4968 7020 4986
rect 7002 4986 7020 5004
rect 7002 5004 7020 5022
rect 7002 5022 7020 5040
rect 7002 5040 7020 5058
rect 7002 5058 7020 5076
rect 7002 5076 7020 5094
rect 7002 5094 7020 5112
rect 7002 5112 7020 5130
rect 7002 5130 7020 5148
rect 7002 5148 7020 5166
rect 7002 5166 7020 5184
rect 7002 5184 7020 5202
rect 7002 5202 7020 5220
rect 7002 5220 7020 5238
rect 7002 5238 7020 5256
rect 7002 5256 7020 5274
rect 7002 5274 7020 5292
rect 7002 5292 7020 5310
rect 7002 5310 7020 5328
rect 7002 5328 7020 5346
rect 7002 5346 7020 5364
rect 7002 5364 7020 5382
rect 7002 5382 7020 5400
rect 7002 5400 7020 5418
rect 7002 5418 7020 5436
rect 7002 5436 7020 5454
rect 7002 5454 7020 5472
rect 7002 5472 7020 5490
rect 7002 5490 7020 5508
rect 7002 5508 7020 5526
rect 7002 5526 7020 5544
rect 7002 5544 7020 5562
rect 7002 5562 7020 5580
rect 7002 5580 7020 5598
rect 7002 5598 7020 5616
rect 7002 5616 7020 5634
rect 7002 5634 7020 5652
rect 7002 5652 7020 5670
rect 7002 5670 7020 5688
rect 7002 5688 7020 5706
rect 7002 5706 7020 5724
rect 7002 5724 7020 5742
rect 7002 5742 7020 5760
rect 7002 5760 7020 5778
rect 7002 5778 7020 5796
rect 7002 5796 7020 5814
rect 7002 5814 7020 5832
rect 7002 5832 7020 5850
rect 7002 5850 7020 5868
rect 7002 5868 7020 5886
rect 7002 5886 7020 5904
rect 7002 5904 7020 5922
rect 7002 5922 7020 5940
rect 7002 5940 7020 5958
rect 7002 5958 7020 5976
rect 7002 5976 7020 5994
rect 7002 5994 7020 6012
rect 7002 6012 7020 6030
rect 7002 6030 7020 6048
rect 7002 6048 7020 6066
rect 7002 6066 7020 6084
rect 7002 6084 7020 6102
rect 7002 6102 7020 6120
rect 7002 6120 7020 6138
rect 7002 6138 7020 6156
rect 7002 6156 7020 6174
rect 7002 6174 7020 6192
rect 7002 6192 7020 6210
rect 7002 6210 7020 6228
rect 7002 6228 7020 6246
rect 7002 6246 7020 6264
rect 7002 7866 7020 7884
rect 7002 7884 7020 7902
rect 7002 7902 7020 7920
rect 7002 7920 7020 7938
rect 7002 7938 7020 7956
rect 7002 7956 7020 7974
rect 7002 7974 7020 7992
rect 7002 7992 7020 8010
rect 7002 8010 7020 8028
rect 7002 8028 7020 8046
rect 7002 8046 7020 8064
rect 7002 8064 7020 8082
rect 7002 8082 7020 8100
rect 7002 8100 7020 8118
rect 7002 8118 7020 8136
rect 7002 8136 7020 8154
rect 7002 8154 7020 8172
rect 7002 8172 7020 8190
rect 7002 8190 7020 8208
rect 7002 8208 7020 8226
rect 7002 8226 7020 8244
rect 7002 8244 7020 8262
rect 7002 8262 7020 8280
rect 7002 8280 7020 8298
rect 7002 8298 7020 8316
rect 7002 8316 7020 8334
rect 7002 8334 7020 8352
rect 7002 8352 7020 8370
rect 7002 8370 7020 8388
rect 7002 8388 7020 8406
rect 7002 8406 7020 8424
rect 7002 8424 7020 8442
rect 7002 8442 7020 8460
rect 7002 8460 7020 8478
rect 7002 8478 7020 8496
rect 7002 8496 7020 8514
rect 7002 8514 7020 8532
rect 7002 8532 7020 8550
rect 7002 8550 7020 8568
rect 7002 8568 7020 8586
rect 7002 8586 7020 8604
rect 7002 8604 7020 8622
rect 7002 8622 7020 8640
rect 7002 8640 7020 8658
rect 7002 8658 7020 8676
rect 7002 8676 7020 8694
rect 7002 8694 7020 8712
rect 7002 8712 7020 8730
rect 7002 8730 7020 8748
rect 7002 8748 7020 8766
rect 7002 8766 7020 8784
rect 7002 8784 7020 8802
rect 7002 8802 7020 8820
rect 7002 8820 7020 8838
rect 7002 8838 7020 8856
rect 7002 8856 7020 8874
rect 7002 8874 7020 8892
rect 7002 8892 7020 8910
rect 7002 8910 7020 8928
rect 7002 8928 7020 8946
rect 7002 8946 7020 8964
rect 7002 8964 7020 8982
rect 7002 8982 7020 9000
rect 7002 9000 7020 9018
rect 7002 9018 7020 9036
rect 7002 9036 7020 9054
rect 7002 9054 7020 9072
rect 7002 9072 7020 9090
rect 7002 9090 7020 9108
rect 7002 9108 7020 9126
rect 7002 9126 7020 9144
rect 7002 9144 7020 9162
rect 7002 9162 7020 9180
rect 7002 9180 7020 9198
rect 7002 9198 7020 9216
rect 7002 9216 7020 9234
rect 7002 9234 7020 9252
rect 7002 9252 7020 9270
rect 7002 9270 7020 9288
rect 7002 9288 7020 9306
rect 7002 9306 7020 9324
rect 7002 9324 7020 9342
rect 7002 9342 7020 9360
rect 7002 9360 7020 9378
rect 7002 9378 7020 9396
rect 7002 9396 7020 9414
rect 7002 9414 7020 9432
rect 7002 9432 7020 9450
rect 7002 9450 7020 9468
rect 7002 9468 7020 9486
rect 7002 9486 7020 9504
rect 7002 9504 7020 9522
rect 7002 9522 7020 9540
rect 7002 9540 7020 9558
rect 7002 9558 7020 9576
rect 7002 9576 7020 9594
rect 7002 9594 7020 9612
rect 7002 9612 7020 9630
rect 7002 9630 7020 9648
rect 7002 9648 7020 9666
rect 7002 9666 7020 9684
rect 7002 9684 7020 9702
rect 7002 9702 7020 9720
rect 7002 9720 7020 9738
rect 7002 9738 7020 9756
rect 7002 9756 7020 9774
rect 7002 9774 7020 9792
rect 7002 9792 7020 9810
rect 7002 9810 7020 9828
rect 7002 9828 7020 9846
rect 7002 9846 7020 9864
rect 7002 9864 7020 9882
rect 7002 9882 7020 9900
rect 7002 9900 7020 9918
rect 7002 9918 7020 9936
rect 7002 9936 7020 9954
rect 7002 9954 7020 9972
rect 7002 9972 7020 9990
rect 7002 9990 7020 10008
rect 7002 10008 7020 10026
rect 7002 10026 7020 10044
rect 7002 10044 7020 10062
rect 7002 10062 7020 10080
rect 7002 10080 7020 10098
rect 7002 10098 7020 10116
rect 7002 10116 7020 10134
rect 7002 10134 7020 10152
rect 7002 10152 7020 10170
rect 7002 10170 7020 10188
rect 7002 10188 7020 10206
rect 7002 10206 7020 10224
rect 7002 10224 7020 10242
rect 7002 10242 7020 10260
rect 7002 10260 7020 10278
rect 7002 10278 7020 10296
rect 7002 10296 7020 10314
rect 7002 10314 7020 10332
rect 7002 10332 7020 10350
rect 7002 10350 7020 10368
rect 7002 10368 7020 10386
rect 7002 10386 7020 10404
rect 7002 10404 7020 10422
rect 7002 10422 7020 10440
rect 7002 10440 7020 10458
rect 7002 10458 7020 10476
rect 7020 1800 7038 1818
rect 7020 1818 7038 1836
rect 7020 1836 7038 1854
rect 7020 1854 7038 1872
rect 7020 1872 7038 1890
rect 7020 1890 7038 1908
rect 7020 1908 7038 1926
rect 7020 1926 7038 1944
rect 7020 1944 7038 1962
rect 7020 1962 7038 1980
rect 7020 1980 7038 1998
rect 7020 1998 7038 2016
rect 7020 2016 7038 2034
rect 7020 2034 7038 2052
rect 7020 2052 7038 2070
rect 7020 2070 7038 2088
rect 7020 2088 7038 2106
rect 7020 2106 7038 2124
rect 7020 2124 7038 2142
rect 7020 2142 7038 2160
rect 7020 2160 7038 2178
rect 7020 2178 7038 2196
rect 7020 2196 7038 2214
rect 7020 2214 7038 2232
rect 7020 2232 7038 2250
rect 7020 2250 7038 2268
rect 7020 2268 7038 2286
rect 7020 2286 7038 2304
rect 7020 2304 7038 2322
rect 7020 2322 7038 2340
rect 7020 2340 7038 2358
rect 7020 2358 7038 2376
rect 7020 2376 7038 2394
rect 7020 2394 7038 2412
rect 7020 2412 7038 2430
rect 7020 2430 7038 2448
rect 7020 2448 7038 2466
rect 7020 2466 7038 2484
rect 7020 2484 7038 2502
rect 7020 2502 7038 2520
rect 7020 2520 7038 2538
rect 7020 2538 7038 2556
rect 7020 2556 7038 2574
rect 7020 2574 7038 2592
rect 7020 2592 7038 2610
rect 7020 2610 7038 2628
rect 7020 2628 7038 2646
rect 7020 2646 7038 2664
rect 7020 2664 7038 2682
rect 7020 2682 7038 2700
rect 7020 2700 7038 2718
rect 7020 2718 7038 2736
rect 7020 2736 7038 2754
rect 7020 2754 7038 2772
rect 7020 2772 7038 2790
rect 7020 2790 7038 2808
rect 7020 2808 7038 2826
rect 7020 2826 7038 2844
rect 7020 2844 7038 2862
rect 7020 2862 7038 2880
rect 7020 2880 7038 2898
rect 7020 2898 7038 2916
rect 7020 2916 7038 2934
rect 7020 2934 7038 2952
rect 7020 2952 7038 2970
rect 7020 2970 7038 2988
rect 7020 2988 7038 3006
rect 7020 3006 7038 3024
rect 7020 3024 7038 3042
rect 7020 3042 7038 3060
rect 7020 3060 7038 3078
rect 7020 3078 7038 3096
rect 7020 3276 7038 3294
rect 7020 3294 7038 3312
rect 7020 3312 7038 3330
rect 7020 3330 7038 3348
rect 7020 3348 7038 3366
rect 7020 3366 7038 3384
rect 7020 3384 7038 3402
rect 7020 3402 7038 3420
rect 7020 3420 7038 3438
rect 7020 3438 7038 3456
rect 7020 3456 7038 3474
rect 7020 3474 7038 3492
rect 7020 3492 7038 3510
rect 7020 3510 7038 3528
rect 7020 3528 7038 3546
rect 7020 3546 7038 3564
rect 7020 3564 7038 3582
rect 7020 3582 7038 3600
rect 7020 3600 7038 3618
rect 7020 3618 7038 3636
rect 7020 3636 7038 3654
rect 7020 3654 7038 3672
rect 7020 3672 7038 3690
rect 7020 3690 7038 3708
rect 7020 3708 7038 3726
rect 7020 3726 7038 3744
rect 7020 3744 7038 3762
rect 7020 3762 7038 3780
rect 7020 3780 7038 3798
rect 7020 3798 7038 3816
rect 7020 3816 7038 3834
rect 7020 4050 7038 4068
rect 7020 4068 7038 4086
rect 7020 4086 7038 4104
rect 7020 4104 7038 4122
rect 7020 4122 7038 4140
rect 7020 4140 7038 4158
rect 7020 4158 7038 4176
rect 7020 4176 7038 4194
rect 7020 4194 7038 4212
rect 7020 4212 7038 4230
rect 7020 4230 7038 4248
rect 7020 4248 7038 4266
rect 7020 4266 7038 4284
rect 7020 4284 7038 4302
rect 7020 4302 7038 4320
rect 7020 4320 7038 4338
rect 7020 4338 7038 4356
rect 7020 4356 7038 4374
rect 7020 4374 7038 4392
rect 7020 4392 7038 4410
rect 7020 4410 7038 4428
rect 7020 4428 7038 4446
rect 7020 4446 7038 4464
rect 7020 4464 7038 4482
rect 7020 4482 7038 4500
rect 7020 4500 7038 4518
rect 7020 4518 7038 4536
rect 7020 4536 7038 4554
rect 7020 4554 7038 4572
rect 7020 4572 7038 4590
rect 7020 4590 7038 4608
rect 7020 4608 7038 4626
rect 7020 4626 7038 4644
rect 7020 4644 7038 4662
rect 7020 4662 7038 4680
rect 7020 4680 7038 4698
rect 7020 4698 7038 4716
rect 7020 4716 7038 4734
rect 7020 4734 7038 4752
rect 7020 4752 7038 4770
rect 7020 4770 7038 4788
rect 7020 4788 7038 4806
rect 7020 4806 7038 4824
rect 7020 4824 7038 4842
rect 7020 4842 7038 4860
rect 7020 4860 7038 4878
rect 7020 4878 7038 4896
rect 7020 4896 7038 4914
rect 7020 4914 7038 4932
rect 7020 4932 7038 4950
rect 7020 4950 7038 4968
rect 7020 4968 7038 4986
rect 7020 4986 7038 5004
rect 7020 5004 7038 5022
rect 7020 5022 7038 5040
rect 7020 5040 7038 5058
rect 7020 5058 7038 5076
rect 7020 5076 7038 5094
rect 7020 5094 7038 5112
rect 7020 5112 7038 5130
rect 7020 5130 7038 5148
rect 7020 5148 7038 5166
rect 7020 5166 7038 5184
rect 7020 5184 7038 5202
rect 7020 5202 7038 5220
rect 7020 5220 7038 5238
rect 7020 5238 7038 5256
rect 7020 5256 7038 5274
rect 7020 5274 7038 5292
rect 7020 5292 7038 5310
rect 7020 5310 7038 5328
rect 7020 5328 7038 5346
rect 7020 5346 7038 5364
rect 7020 5364 7038 5382
rect 7020 5382 7038 5400
rect 7020 5400 7038 5418
rect 7020 5418 7038 5436
rect 7020 5436 7038 5454
rect 7020 5454 7038 5472
rect 7020 5472 7038 5490
rect 7020 5490 7038 5508
rect 7020 5508 7038 5526
rect 7020 5526 7038 5544
rect 7020 5544 7038 5562
rect 7020 5562 7038 5580
rect 7020 5580 7038 5598
rect 7020 5598 7038 5616
rect 7020 5616 7038 5634
rect 7020 5634 7038 5652
rect 7020 5652 7038 5670
rect 7020 5670 7038 5688
rect 7020 5688 7038 5706
rect 7020 5706 7038 5724
rect 7020 5724 7038 5742
rect 7020 5742 7038 5760
rect 7020 5760 7038 5778
rect 7020 5778 7038 5796
rect 7020 5796 7038 5814
rect 7020 5814 7038 5832
rect 7020 5832 7038 5850
rect 7020 5850 7038 5868
rect 7020 5868 7038 5886
rect 7020 5886 7038 5904
rect 7020 5904 7038 5922
rect 7020 5922 7038 5940
rect 7020 5940 7038 5958
rect 7020 5958 7038 5976
rect 7020 5976 7038 5994
rect 7020 5994 7038 6012
rect 7020 6012 7038 6030
rect 7020 6030 7038 6048
rect 7020 6048 7038 6066
rect 7020 6066 7038 6084
rect 7020 6084 7038 6102
rect 7020 6102 7038 6120
rect 7020 6120 7038 6138
rect 7020 6138 7038 6156
rect 7020 6156 7038 6174
rect 7020 6174 7038 6192
rect 7020 6192 7038 6210
rect 7020 6210 7038 6228
rect 7020 6228 7038 6246
rect 7020 6246 7038 6264
rect 7020 6264 7038 6282
rect 7020 7920 7038 7938
rect 7020 7938 7038 7956
rect 7020 7956 7038 7974
rect 7020 7974 7038 7992
rect 7020 7992 7038 8010
rect 7020 8010 7038 8028
rect 7020 8028 7038 8046
rect 7020 8046 7038 8064
rect 7020 8064 7038 8082
rect 7020 8082 7038 8100
rect 7020 8100 7038 8118
rect 7020 8118 7038 8136
rect 7020 8136 7038 8154
rect 7020 8154 7038 8172
rect 7020 8172 7038 8190
rect 7020 8190 7038 8208
rect 7020 8208 7038 8226
rect 7020 8226 7038 8244
rect 7020 8244 7038 8262
rect 7020 8262 7038 8280
rect 7020 8280 7038 8298
rect 7020 8298 7038 8316
rect 7020 8316 7038 8334
rect 7020 8334 7038 8352
rect 7020 8352 7038 8370
rect 7020 8370 7038 8388
rect 7020 8388 7038 8406
rect 7020 8406 7038 8424
rect 7020 8424 7038 8442
rect 7020 8442 7038 8460
rect 7020 8460 7038 8478
rect 7020 8478 7038 8496
rect 7020 8496 7038 8514
rect 7020 8514 7038 8532
rect 7020 8532 7038 8550
rect 7020 8550 7038 8568
rect 7020 8568 7038 8586
rect 7020 8586 7038 8604
rect 7020 8604 7038 8622
rect 7020 8622 7038 8640
rect 7020 8640 7038 8658
rect 7020 8658 7038 8676
rect 7020 8676 7038 8694
rect 7020 8694 7038 8712
rect 7020 8712 7038 8730
rect 7020 8730 7038 8748
rect 7020 8748 7038 8766
rect 7020 8766 7038 8784
rect 7020 8784 7038 8802
rect 7020 8802 7038 8820
rect 7020 8820 7038 8838
rect 7020 8838 7038 8856
rect 7020 8856 7038 8874
rect 7020 8874 7038 8892
rect 7020 8892 7038 8910
rect 7020 8910 7038 8928
rect 7020 8928 7038 8946
rect 7020 8946 7038 8964
rect 7020 8964 7038 8982
rect 7020 8982 7038 9000
rect 7020 9000 7038 9018
rect 7020 9018 7038 9036
rect 7020 9036 7038 9054
rect 7020 9054 7038 9072
rect 7020 9072 7038 9090
rect 7020 9090 7038 9108
rect 7020 9108 7038 9126
rect 7020 9126 7038 9144
rect 7020 9144 7038 9162
rect 7020 9162 7038 9180
rect 7020 9180 7038 9198
rect 7020 9198 7038 9216
rect 7020 9216 7038 9234
rect 7020 9234 7038 9252
rect 7020 9252 7038 9270
rect 7020 9270 7038 9288
rect 7020 9288 7038 9306
rect 7020 9306 7038 9324
rect 7020 9324 7038 9342
rect 7020 9342 7038 9360
rect 7020 9360 7038 9378
rect 7020 9378 7038 9396
rect 7020 9396 7038 9414
rect 7020 9414 7038 9432
rect 7020 9432 7038 9450
rect 7020 9450 7038 9468
rect 7020 9468 7038 9486
rect 7020 9486 7038 9504
rect 7020 9504 7038 9522
rect 7020 9522 7038 9540
rect 7020 9540 7038 9558
rect 7020 9558 7038 9576
rect 7020 9576 7038 9594
rect 7020 9594 7038 9612
rect 7020 9612 7038 9630
rect 7020 9630 7038 9648
rect 7020 9648 7038 9666
rect 7020 9666 7038 9684
rect 7020 9684 7038 9702
rect 7020 9702 7038 9720
rect 7020 9720 7038 9738
rect 7020 9738 7038 9756
rect 7020 9756 7038 9774
rect 7020 9774 7038 9792
rect 7020 9792 7038 9810
rect 7020 9810 7038 9828
rect 7020 9828 7038 9846
rect 7020 9846 7038 9864
rect 7020 9864 7038 9882
rect 7020 9882 7038 9900
rect 7020 9900 7038 9918
rect 7020 9918 7038 9936
rect 7020 9936 7038 9954
rect 7020 9954 7038 9972
rect 7020 9972 7038 9990
rect 7020 9990 7038 10008
rect 7020 10008 7038 10026
rect 7020 10026 7038 10044
rect 7020 10044 7038 10062
rect 7020 10062 7038 10080
rect 7020 10080 7038 10098
rect 7020 10098 7038 10116
rect 7020 10116 7038 10134
rect 7020 10134 7038 10152
rect 7020 10152 7038 10170
rect 7020 10170 7038 10188
rect 7020 10188 7038 10206
rect 7020 10206 7038 10224
rect 7020 10224 7038 10242
rect 7020 10242 7038 10260
rect 7020 10260 7038 10278
rect 7020 10278 7038 10296
rect 7020 10296 7038 10314
rect 7020 10314 7038 10332
rect 7020 10332 7038 10350
rect 7020 10350 7038 10368
rect 7020 10368 7038 10386
rect 7020 10386 7038 10404
rect 7020 10404 7038 10422
rect 7020 10422 7038 10440
rect 7020 10440 7038 10458
rect 7020 10458 7038 10476
rect 7020 10476 7038 10494
rect 7020 10494 7038 10512
rect 7038 1818 7056 1836
rect 7038 1836 7056 1854
rect 7038 1854 7056 1872
rect 7038 1872 7056 1890
rect 7038 1890 7056 1908
rect 7038 1908 7056 1926
rect 7038 1926 7056 1944
rect 7038 1944 7056 1962
rect 7038 1962 7056 1980
rect 7038 1980 7056 1998
rect 7038 1998 7056 2016
rect 7038 2016 7056 2034
rect 7038 2034 7056 2052
rect 7038 2052 7056 2070
rect 7038 2070 7056 2088
rect 7038 2088 7056 2106
rect 7038 2106 7056 2124
rect 7038 2124 7056 2142
rect 7038 2142 7056 2160
rect 7038 2160 7056 2178
rect 7038 2178 7056 2196
rect 7038 2196 7056 2214
rect 7038 2214 7056 2232
rect 7038 2232 7056 2250
rect 7038 2250 7056 2268
rect 7038 2268 7056 2286
rect 7038 2286 7056 2304
rect 7038 2304 7056 2322
rect 7038 2322 7056 2340
rect 7038 2340 7056 2358
rect 7038 2358 7056 2376
rect 7038 2376 7056 2394
rect 7038 2394 7056 2412
rect 7038 2412 7056 2430
rect 7038 2430 7056 2448
rect 7038 2448 7056 2466
rect 7038 2466 7056 2484
rect 7038 2484 7056 2502
rect 7038 2502 7056 2520
rect 7038 2520 7056 2538
rect 7038 2538 7056 2556
rect 7038 2556 7056 2574
rect 7038 2574 7056 2592
rect 7038 2592 7056 2610
rect 7038 2610 7056 2628
rect 7038 2628 7056 2646
rect 7038 2646 7056 2664
rect 7038 2664 7056 2682
rect 7038 2682 7056 2700
rect 7038 2700 7056 2718
rect 7038 2718 7056 2736
rect 7038 2736 7056 2754
rect 7038 2754 7056 2772
rect 7038 2772 7056 2790
rect 7038 2790 7056 2808
rect 7038 2808 7056 2826
rect 7038 2826 7056 2844
rect 7038 2844 7056 2862
rect 7038 2862 7056 2880
rect 7038 2880 7056 2898
rect 7038 2898 7056 2916
rect 7038 2916 7056 2934
rect 7038 2934 7056 2952
rect 7038 2952 7056 2970
rect 7038 2970 7056 2988
rect 7038 2988 7056 3006
rect 7038 3006 7056 3024
rect 7038 3024 7056 3042
rect 7038 3042 7056 3060
rect 7038 3060 7056 3078
rect 7038 3078 7056 3096
rect 7038 3294 7056 3312
rect 7038 3312 7056 3330
rect 7038 3330 7056 3348
rect 7038 3348 7056 3366
rect 7038 3366 7056 3384
rect 7038 3384 7056 3402
rect 7038 3402 7056 3420
rect 7038 3420 7056 3438
rect 7038 3438 7056 3456
rect 7038 3456 7056 3474
rect 7038 3474 7056 3492
rect 7038 3492 7056 3510
rect 7038 3510 7056 3528
rect 7038 3528 7056 3546
rect 7038 3546 7056 3564
rect 7038 3564 7056 3582
rect 7038 3582 7056 3600
rect 7038 3600 7056 3618
rect 7038 3618 7056 3636
rect 7038 3636 7056 3654
rect 7038 3654 7056 3672
rect 7038 3672 7056 3690
rect 7038 3690 7056 3708
rect 7038 3708 7056 3726
rect 7038 3726 7056 3744
rect 7038 3744 7056 3762
rect 7038 3762 7056 3780
rect 7038 3780 7056 3798
rect 7038 3798 7056 3816
rect 7038 3816 7056 3834
rect 7038 3834 7056 3852
rect 7038 3852 7056 3870
rect 7038 4068 7056 4086
rect 7038 4086 7056 4104
rect 7038 4104 7056 4122
rect 7038 4122 7056 4140
rect 7038 4140 7056 4158
rect 7038 4158 7056 4176
rect 7038 4176 7056 4194
rect 7038 4194 7056 4212
rect 7038 4212 7056 4230
rect 7038 4230 7056 4248
rect 7038 4248 7056 4266
rect 7038 4266 7056 4284
rect 7038 4284 7056 4302
rect 7038 4302 7056 4320
rect 7038 4320 7056 4338
rect 7038 4338 7056 4356
rect 7038 4356 7056 4374
rect 7038 4374 7056 4392
rect 7038 4392 7056 4410
rect 7038 4410 7056 4428
rect 7038 4428 7056 4446
rect 7038 4446 7056 4464
rect 7038 4464 7056 4482
rect 7038 4482 7056 4500
rect 7038 4500 7056 4518
rect 7038 4518 7056 4536
rect 7038 4536 7056 4554
rect 7038 4554 7056 4572
rect 7038 4572 7056 4590
rect 7038 4590 7056 4608
rect 7038 4608 7056 4626
rect 7038 4626 7056 4644
rect 7038 4644 7056 4662
rect 7038 4662 7056 4680
rect 7038 4680 7056 4698
rect 7038 4698 7056 4716
rect 7038 4716 7056 4734
rect 7038 4734 7056 4752
rect 7038 4752 7056 4770
rect 7038 4770 7056 4788
rect 7038 4788 7056 4806
rect 7038 4806 7056 4824
rect 7038 4824 7056 4842
rect 7038 4842 7056 4860
rect 7038 4860 7056 4878
rect 7038 4878 7056 4896
rect 7038 4896 7056 4914
rect 7038 4914 7056 4932
rect 7038 4932 7056 4950
rect 7038 4950 7056 4968
rect 7038 4968 7056 4986
rect 7038 4986 7056 5004
rect 7038 5004 7056 5022
rect 7038 5022 7056 5040
rect 7038 5040 7056 5058
rect 7038 5058 7056 5076
rect 7038 5076 7056 5094
rect 7038 5094 7056 5112
rect 7038 5112 7056 5130
rect 7038 5130 7056 5148
rect 7038 5148 7056 5166
rect 7038 5166 7056 5184
rect 7038 5184 7056 5202
rect 7038 5202 7056 5220
rect 7038 5220 7056 5238
rect 7038 5238 7056 5256
rect 7038 5256 7056 5274
rect 7038 5274 7056 5292
rect 7038 5292 7056 5310
rect 7038 5310 7056 5328
rect 7038 5328 7056 5346
rect 7038 5346 7056 5364
rect 7038 5364 7056 5382
rect 7038 5382 7056 5400
rect 7038 5400 7056 5418
rect 7038 5418 7056 5436
rect 7038 5436 7056 5454
rect 7038 5454 7056 5472
rect 7038 5472 7056 5490
rect 7038 5490 7056 5508
rect 7038 5508 7056 5526
rect 7038 5526 7056 5544
rect 7038 5544 7056 5562
rect 7038 5562 7056 5580
rect 7038 5580 7056 5598
rect 7038 5598 7056 5616
rect 7038 5616 7056 5634
rect 7038 5634 7056 5652
rect 7038 5652 7056 5670
rect 7038 5670 7056 5688
rect 7038 5688 7056 5706
rect 7038 5706 7056 5724
rect 7038 5724 7056 5742
rect 7038 5742 7056 5760
rect 7038 5760 7056 5778
rect 7038 5778 7056 5796
rect 7038 5796 7056 5814
rect 7038 5814 7056 5832
rect 7038 5832 7056 5850
rect 7038 5850 7056 5868
rect 7038 5868 7056 5886
rect 7038 5886 7056 5904
rect 7038 5904 7056 5922
rect 7038 5922 7056 5940
rect 7038 5940 7056 5958
rect 7038 5958 7056 5976
rect 7038 5976 7056 5994
rect 7038 5994 7056 6012
rect 7038 6012 7056 6030
rect 7038 6030 7056 6048
rect 7038 6048 7056 6066
rect 7038 6066 7056 6084
rect 7038 6084 7056 6102
rect 7038 6102 7056 6120
rect 7038 6120 7056 6138
rect 7038 6138 7056 6156
rect 7038 6156 7056 6174
rect 7038 6174 7056 6192
rect 7038 6192 7056 6210
rect 7038 6210 7056 6228
rect 7038 6228 7056 6246
rect 7038 6246 7056 6264
rect 7038 6264 7056 6282
rect 7038 6282 7056 6300
rect 7038 7974 7056 7992
rect 7038 7992 7056 8010
rect 7038 8010 7056 8028
rect 7038 8028 7056 8046
rect 7038 8046 7056 8064
rect 7038 8064 7056 8082
rect 7038 8082 7056 8100
rect 7038 8100 7056 8118
rect 7038 8118 7056 8136
rect 7038 8136 7056 8154
rect 7038 8154 7056 8172
rect 7038 8172 7056 8190
rect 7038 8190 7056 8208
rect 7038 8208 7056 8226
rect 7038 8226 7056 8244
rect 7038 8244 7056 8262
rect 7038 8262 7056 8280
rect 7038 8280 7056 8298
rect 7038 8298 7056 8316
rect 7038 8316 7056 8334
rect 7038 8334 7056 8352
rect 7038 8352 7056 8370
rect 7038 8370 7056 8388
rect 7038 8388 7056 8406
rect 7038 8406 7056 8424
rect 7038 8424 7056 8442
rect 7038 8442 7056 8460
rect 7038 8460 7056 8478
rect 7038 8478 7056 8496
rect 7038 8496 7056 8514
rect 7038 8514 7056 8532
rect 7038 8532 7056 8550
rect 7038 8550 7056 8568
rect 7038 8568 7056 8586
rect 7038 8586 7056 8604
rect 7038 8604 7056 8622
rect 7038 8622 7056 8640
rect 7038 8640 7056 8658
rect 7038 8658 7056 8676
rect 7038 8676 7056 8694
rect 7038 8694 7056 8712
rect 7038 8712 7056 8730
rect 7038 8730 7056 8748
rect 7038 8748 7056 8766
rect 7038 8766 7056 8784
rect 7038 8784 7056 8802
rect 7038 8802 7056 8820
rect 7038 8820 7056 8838
rect 7038 8838 7056 8856
rect 7038 8856 7056 8874
rect 7038 8874 7056 8892
rect 7038 8892 7056 8910
rect 7038 8910 7056 8928
rect 7038 8928 7056 8946
rect 7038 8946 7056 8964
rect 7038 8964 7056 8982
rect 7038 8982 7056 9000
rect 7038 9000 7056 9018
rect 7038 9018 7056 9036
rect 7038 9036 7056 9054
rect 7038 9054 7056 9072
rect 7038 9072 7056 9090
rect 7038 9090 7056 9108
rect 7038 9108 7056 9126
rect 7038 9126 7056 9144
rect 7038 9144 7056 9162
rect 7038 9162 7056 9180
rect 7038 9180 7056 9198
rect 7038 9198 7056 9216
rect 7038 9216 7056 9234
rect 7038 9234 7056 9252
rect 7038 9252 7056 9270
rect 7038 9270 7056 9288
rect 7038 9288 7056 9306
rect 7038 9306 7056 9324
rect 7038 9324 7056 9342
rect 7038 9342 7056 9360
rect 7038 9360 7056 9378
rect 7038 9378 7056 9396
rect 7038 9396 7056 9414
rect 7038 9414 7056 9432
rect 7038 9432 7056 9450
rect 7038 9450 7056 9468
rect 7038 9468 7056 9486
rect 7038 9486 7056 9504
rect 7038 9504 7056 9522
rect 7038 9522 7056 9540
rect 7038 9540 7056 9558
rect 7038 9558 7056 9576
rect 7038 9576 7056 9594
rect 7038 9594 7056 9612
rect 7038 9612 7056 9630
rect 7038 9630 7056 9648
rect 7038 9648 7056 9666
rect 7038 9666 7056 9684
rect 7038 9684 7056 9702
rect 7038 9702 7056 9720
rect 7038 9720 7056 9738
rect 7038 9738 7056 9756
rect 7038 9756 7056 9774
rect 7038 9774 7056 9792
rect 7038 9792 7056 9810
rect 7038 9810 7056 9828
rect 7038 9828 7056 9846
rect 7038 9846 7056 9864
rect 7038 9864 7056 9882
rect 7038 9882 7056 9900
rect 7038 9900 7056 9918
rect 7038 9918 7056 9936
rect 7038 9936 7056 9954
rect 7038 9954 7056 9972
rect 7038 9972 7056 9990
rect 7038 9990 7056 10008
rect 7038 10008 7056 10026
rect 7038 10026 7056 10044
rect 7038 10044 7056 10062
rect 7038 10062 7056 10080
rect 7038 10080 7056 10098
rect 7038 10098 7056 10116
rect 7038 10116 7056 10134
rect 7038 10134 7056 10152
rect 7038 10152 7056 10170
rect 7038 10170 7056 10188
rect 7038 10188 7056 10206
rect 7038 10206 7056 10224
rect 7038 10224 7056 10242
rect 7038 10242 7056 10260
rect 7038 10260 7056 10278
rect 7038 10278 7056 10296
rect 7038 10296 7056 10314
rect 7038 10314 7056 10332
rect 7038 10332 7056 10350
rect 7038 10350 7056 10368
rect 7038 10368 7056 10386
rect 7038 10386 7056 10404
rect 7038 10404 7056 10422
rect 7038 10422 7056 10440
rect 7038 10440 7056 10458
rect 7038 10458 7056 10476
rect 7038 10476 7056 10494
rect 7038 10494 7056 10512
rect 7038 10512 7056 10530
rect 7056 1818 7074 1836
rect 7056 1836 7074 1854
rect 7056 1854 7074 1872
rect 7056 1872 7074 1890
rect 7056 1890 7074 1908
rect 7056 1908 7074 1926
rect 7056 1926 7074 1944
rect 7056 1944 7074 1962
rect 7056 1962 7074 1980
rect 7056 1980 7074 1998
rect 7056 1998 7074 2016
rect 7056 2016 7074 2034
rect 7056 2034 7074 2052
rect 7056 2052 7074 2070
rect 7056 2070 7074 2088
rect 7056 2088 7074 2106
rect 7056 2106 7074 2124
rect 7056 2124 7074 2142
rect 7056 2142 7074 2160
rect 7056 2160 7074 2178
rect 7056 2178 7074 2196
rect 7056 2196 7074 2214
rect 7056 2214 7074 2232
rect 7056 2232 7074 2250
rect 7056 2250 7074 2268
rect 7056 2268 7074 2286
rect 7056 2286 7074 2304
rect 7056 2304 7074 2322
rect 7056 2322 7074 2340
rect 7056 2340 7074 2358
rect 7056 2358 7074 2376
rect 7056 2376 7074 2394
rect 7056 2394 7074 2412
rect 7056 2412 7074 2430
rect 7056 2430 7074 2448
rect 7056 2448 7074 2466
rect 7056 2466 7074 2484
rect 7056 2484 7074 2502
rect 7056 2502 7074 2520
rect 7056 2520 7074 2538
rect 7056 2538 7074 2556
rect 7056 2556 7074 2574
rect 7056 2574 7074 2592
rect 7056 2592 7074 2610
rect 7056 2610 7074 2628
rect 7056 2628 7074 2646
rect 7056 2646 7074 2664
rect 7056 2664 7074 2682
rect 7056 2682 7074 2700
rect 7056 2700 7074 2718
rect 7056 2718 7074 2736
rect 7056 2736 7074 2754
rect 7056 2754 7074 2772
rect 7056 2772 7074 2790
rect 7056 2790 7074 2808
rect 7056 2808 7074 2826
rect 7056 2826 7074 2844
rect 7056 2844 7074 2862
rect 7056 2862 7074 2880
rect 7056 2880 7074 2898
rect 7056 2898 7074 2916
rect 7056 2916 7074 2934
rect 7056 2934 7074 2952
rect 7056 2952 7074 2970
rect 7056 2970 7074 2988
rect 7056 2988 7074 3006
rect 7056 3006 7074 3024
rect 7056 3024 7074 3042
rect 7056 3042 7074 3060
rect 7056 3060 7074 3078
rect 7056 3078 7074 3096
rect 7056 3096 7074 3114
rect 7056 3294 7074 3312
rect 7056 3312 7074 3330
rect 7056 3330 7074 3348
rect 7056 3348 7074 3366
rect 7056 3366 7074 3384
rect 7056 3384 7074 3402
rect 7056 3402 7074 3420
rect 7056 3420 7074 3438
rect 7056 3438 7074 3456
rect 7056 3456 7074 3474
rect 7056 3474 7074 3492
rect 7056 3492 7074 3510
rect 7056 3510 7074 3528
rect 7056 3528 7074 3546
rect 7056 3546 7074 3564
rect 7056 3564 7074 3582
rect 7056 3582 7074 3600
rect 7056 3600 7074 3618
rect 7056 3618 7074 3636
rect 7056 3636 7074 3654
rect 7056 3654 7074 3672
rect 7056 3672 7074 3690
rect 7056 3690 7074 3708
rect 7056 3708 7074 3726
rect 7056 3726 7074 3744
rect 7056 3744 7074 3762
rect 7056 3762 7074 3780
rect 7056 3780 7074 3798
rect 7056 3798 7074 3816
rect 7056 3816 7074 3834
rect 7056 3834 7074 3852
rect 7056 3852 7074 3870
rect 7056 3870 7074 3888
rect 7056 4104 7074 4122
rect 7056 4122 7074 4140
rect 7056 4140 7074 4158
rect 7056 4158 7074 4176
rect 7056 4176 7074 4194
rect 7056 4194 7074 4212
rect 7056 4212 7074 4230
rect 7056 4230 7074 4248
rect 7056 4248 7074 4266
rect 7056 4266 7074 4284
rect 7056 4284 7074 4302
rect 7056 4302 7074 4320
rect 7056 4320 7074 4338
rect 7056 4338 7074 4356
rect 7056 4356 7074 4374
rect 7056 4374 7074 4392
rect 7056 4392 7074 4410
rect 7056 4410 7074 4428
rect 7056 4428 7074 4446
rect 7056 4446 7074 4464
rect 7056 4464 7074 4482
rect 7056 4482 7074 4500
rect 7056 4500 7074 4518
rect 7056 4518 7074 4536
rect 7056 4536 7074 4554
rect 7056 4554 7074 4572
rect 7056 4572 7074 4590
rect 7056 4590 7074 4608
rect 7056 4608 7074 4626
rect 7056 4626 7074 4644
rect 7056 4644 7074 4662
rect 7056 4662 7074 4680
rect 7056 4680 7074 4698
rect 7056 4698 7074 4716
rect 7056 4716 7074 4734
rect 7056 4734 7074 4752
rect 7056 4752 7074 4770
rect 7056 4770 7074 4788
rect 7056 4788 7074 4806
rect 7056 4806 7074 4824
rect 7056 4824 7074 4842
rect 7056 4842 7074 4860
rect 7056 4860 7074 4878
rect 7056 4878 7074 4896
rect 7056 4896 7074 4914
rect 7056 4914 7074 4932
rect 7056 4932 7074 4950
rect 7056 4950 7074 4968
rect 7056 4968 7074 4986
rect 7056 4986 7074 5004
rect 7056 5004 7074 5022
rect 7056 5022 7074 5040
rect 7056 5040 7074 5058
rect 7056 5058 7074 5076
rect 7056 5076 7074 5094
rect 7056 5094 7074 5112
rect 7056 5112 7074 5130
rect 7056 5130 7074 5148
rect 7056 5148 7074 5166
rect 7056 5166 7074 5184
rect 7056 5184 7074 5202
rect 7056 5202 7074 5220
rect 7056 5220 7074 5238
rect 7056 5238 7074 5256
rect 7056 5256 7074 5274
rect 7056 5274 7074 5292
rect 7056 5292 7074 5310
rect 7056 5310 7074 5328
rect 7056 5328 7074 5346
rect 7056 5346 7074 5364
rect 7056 5364 7074 5382
rect 7056 5382 7074 5400
rect 7056 5400 7074 5418
rect 7056 5418 7074 5436
rect 7056 5436 7074 5454
rect 7056 5454 7074 5472
rect 7056 5472 7074 5490
rect 7056 5490 7074 5508
rect 7056 5508 7074 5526
rect 7056 5526 7074 5544
rect 7056 5544 7074 5562
rect 7056 5562 7074 5580
rect 7056 5580 7074 5598
rect 7056 5598 7074 5616
rect 7056 5616 7074 5634
rect 7056 5634 7074 5652
rect 7056 5652 7074 5670
rect 7056 5670 7074 5688
rect 7056 5688 7074 5706
rect 7056 5706 7074 5724
rect 7056 5724 7074 5742
rect 7056 5742 7074 5760
rect 7056 5760 7074 5778
rect 7056 5778 7074 5796
rect 7056 5796 7074 5814
rect 7056 5814 7074 5832
rect 7056 5832 7074 5850
rect 7056 5850 7074 5868
rect 7056 5868 7074 5886
rect 7056 5886 7074 5904
rect 7056 5904 7074 5922
rect 7056 5922 7074 5940
rect 7056 5940 7074 5958
rect 7056 5958 7074 5976
rect 7056 5976 7074 5994
rect 7056 5994 7074 6012
rect 7056 6012 7074 6030
rect 7056 6030 7074 6048
rect 7056 6048 7074 6066
rect 7056 6066 7074 6084
rect 7056 6084 7074 6102
rect 7056 6102 7074 6120
rect 7056 6120 7074 6138
rect 7056 6138 7074 6156
rect 7056 6156 7074 6174
rect 7056 6174 7074 6192
rect 7056 6192 7074 6210
rect 7056 6210 7074 6228
rect 7056 6228 7074 6246
rect 7056 6246 7074 6264
rect 7056 6264 7074 6282
rect 7056 6282 7074 6300
rect 7056 8028 7074 8046
rect 7056 8046 7074 8064
rect 7056 8064 7074 8082
rect 7056 8082 7074 8100
rect 7056 8100 7074 8118
rect 7056 8118 7074 8136
rect 7056 8136 7074 8154
rect 7056 8154 7074 8172
rect 7056 8172 7074 8190
rect 7056 8190 7074 8208
rect 7056 8208 7074 8226
rect 7056 8226 7074 8244
rect 7056 8244 7074 8262
rect 7056 8262 7074 8280
rect 7056 8280 7074 8298
rect 7056 8298 7074 8316
rect 7056 8316 7074 8334
rect 7056 8334 7074 8352
rect 7056 8352 7074 8370
rect 7056 8370 7074 8388
rect 7056 8388 7074 8406
rect 7056 8406 7074 8424
rect 7056 8424 7074 8442
rect 7056 8442 7074 8460
rect 7056 8460 7074 8478
rect 7056 8478 7074 8496
rect 7056 8496 7074 8514
rect 7056 8514 7074 8532
rect 7056 8532 7074 8550
rect 7056 8550 7074 8568
rect 7056 8568 7074 8586
rect 7056 8586 7074 8604
rect 7056 8604 7074 8622
rect 7056 8622 7074 8640
rect 7056 8640 7074 8658
rect 7056 8658 7074 8676
rect 7056 8676 7074 8694
rect 7056 8694 7074 8712
rect 7056 8712 7074 8730
rect 7056 8730 7074 8748
rect 7056 8748 7074 8766
rect 7056 8766 7074 8784
rect 7056 8784 7074 8802
rect 7056 8802 7074 8820
rect 7056 8820 7074 8838
rect 7056 8838 7074 8856
rect 7056 8856 7074 8874
rect 7056 8874 7074 8892
rect 7056 8892 7074 8910
rect 7056 8910 7074 8928
rect 7056 8928 7074 8946
rect 7056 8946 7074 8964
rect 7056 8964 7074 8982
rect 7056 8982 7074 9000
rect 7056 9000 7074 9018
rect 7056 9018 7074 9036
rect 7056 9036 7074 9054
rect 7056 9054 7074 9072
rect 7056 9072 7074 9090
rect 7056 9090 7074 9108
rect 7056 9108 7074 9126
rect 7056 9126 7074 9144
rect 7056 9144 7074 9162
rect 7056 9162 7074 9180
rect 7056 9180 7074 9198
rect 7056 9198 7074 9216
rect 7056 9216 7074 9234
rect 7056 9234 7074 9252
rect 7056 9252 7074 9270
rect 7056 9270 7074 9288
rect 7056 9288 7074 9306
rect 7056 9306 7074 9324
rect 7056 9324 7074 9342
rect 7056 9342 7074 9360
rect 7056 9360 7074 9378
rect 7056 9378 7074 9396
rect 7056 9396 7074 9414
rect 7056 9414 7074 9432
rect 7056 9432 7074 9450
rect 7056 9450 7074 9468
rect 7056 9468 7074 9486
rect 7056 9486 7074 9504
rect 7056 9504 7074 9522
rect 7056 9522 7074 9540
rect 7056 9540 7074 9558
rect 7056 9558 7074 9576
rect 7056 9576 7074 9594
rect 7056 9594 7074 9612
rect 7056 9612 7074 9630
rect 7056 9630 7074 9648
rect 7056 9648 7074 9666
rect 7056 9666 7074 9684
rect 7056 9684 7074 9702
rect 7056 9702 7074 9720
rect 7056 9720 7074 9738
rect 7056 9738 7074 9756
rect 7056 9756 7074 9774
rect 7056 9774 7074 9792
rect 7056 9792 7074 9810
rect 7056 9810 7074 9828
rect 7056 9828 7074 9846
rect 7056 9846 7074 9864
rect 7056 9864 7074 9882
rect 7056 9882 7074 9900
rect 7056 9900 7074 9918
rect 7056 9918 7074 9936
rect 7056 9936 7074 9954
rect 7056 9954 7074 9972
rect 7056 9972 7074 9990
rect 7056 9990 7074 10008
rect 7056 10008 7074 10026
rect 7056 10026 7074 10044
rect 7056 10044 7074 10062
rect 7056 10062 7074 10080
rect 7056 10080 7074 10098
rect 7056 10098 7074 10116
rect 7056 10116 7074 10134
rect 7056 10134 7074 10152
rect 7056 10152 7074 10170
rect 7056 10170 7074 10188
rect 7056 10188 7074 10206
rect 7056 10206 7074 10224
rect 7056 10224 7074 10242
rect 7056 10242 7074 10260
rect 7056 10260 7074 10278
rect 7056 10278 7074 10296
rect 7056 10296 7074 10314
rect 7056 10314 7074 10332
rect 7056 10332 7074 10350
rect 7056 10350 7074 10368
rect 7056 10368 7074 10386
rect 7056 10386 7074 10404
rect 7056 10404 7074 10422
rect 7056 10422 7074 10440
rect 7056 10440 7074 10458
rect 7056 10458 7074 10476
rect 7056 10476 7074 10494
rect 7056 10494 7074 10512
rect 7056 10512 7074 10530
rect 7056 10530 7074 10548
rect 7074 1836 7092 1854
rect 7074 1854 7092 1872
rect 7074 1872 7092 1890
rect 7074 1890 7092 1908
rect 7074 1908 7092 1926
rect 7074 1926 7092 1944
rect 7074 1944 7092 1962
rect 7074 1962 7092 1980
rect 7074 1980 7092 1998
rect 7074 1998 7092 2016
rect 7074 2016 7092 2034
rect 7074 2034 7092 2052
rect 7074 2052 7092 2070
rect 7074 2070 7092 2088
rect 7074 2088 7092 2106
rect 7074 2106 7092 2124
rect 7074 2124 7092 2142
rect 7074 2142 7092 2160
rect 7074 2160 7092 2178
rect 7074 2178 7092 2196
rect 7074 2196 7092 2214
rect 7074 2214 7092 2232
rect 7074 2232 7092 2250
rect 7074 2250 7092 2268
rect 7074 2268 7092 2286
rect 7074 2286 7092 2304
rect 7074 2304 7092 2322
rect 7074 2322 7092 2340
rect 7074 2340 7092 2358
rect 7074 2358 7092 2376
rect 7074 2376 7092 2394
rect 7074 2394 7092 2412
rect 7074 2412 7092 2430
rect 7074 2430 7092 2448
rect 7074 2448 7092 2466
rect 7074 2466 7092 2484
rect 7074 2484 7092 2502
rect 7074 2502 7092 2520
rect 7074 2520 7092 2538
rect 7074 2538 7092 2556
rect 7074 2556 7092 2574
rect 7074 2574 7092 2592
rect 7074 2592 7092 2610
rect 7074 2610 7092 2628
rect 7074 2628 7092 2646
rect 7074 2646 7092 2664
rect 7074 2664 7092 2682
rect 7074 2682 7092 2700
rect 7074 2700 7092 2718
rect 7074 2718 7092 2736
rect 7074 2736 7092 2754
rect 7074 2754 7092 2772
rect 7074 2772 7092 2790
rect 7074 2790 7092 2808
rect 7074 2808 7092 2826
rect 7074 2826 7092 2844
rect 7074 2844 7092 2862
rect 7074 2862 7092 2880
rect 7074 2880 7092 2898
rect 7074 2898 7092 2916
rect 7074 2916 7092 2934
rect 7074 2934 7092 2952
rect 7074 2952 7092 2970
rect 7074 2970 7092 2988
rect 7074 2988 7092 3006
rect 7074 3006 7092 3024
rect 7074 3024 7092 3042
rect 7074 3042 7092 3060
rect 7074 3060 7092 3078
rect 7074 3078 7092 3096
rect 7074 3096 7092 3114
rect 7074 3294 7092 3312
rect 7074 3312 7092 3330
rect 7074 3330 7092 3348
rect 7074 3348 7092 3366
rect 7074 3366 7092 3384
rect 7074 3384 7092 3402
rect 7074 3402 7092 3420
rect 7074 3420 7092 3438
rect 7074 3438 7092 3456
rect 7074 3456 7092 3474
rect 7074 3474 7092 3492
rect 7074 3492 7092 3510
rect 7074 3510 7092 3528
rect 7074 3528 7092 3546
rect 7074 3546 7092 3564
rect 7074 3564 7092 3582
rect 7074 3582 7092 3600
rect 7074 3600 7092 3618
rect 7074 3618 7092 3636
rect 7074 3636 7092 3654
rect 7074 3654 7092 3672
rect 7074 3672 7092 3690
rect 7074 3690 7092 3708
rect 7074 3708 7092 3726
rect 7074 3726 7092 3744
rect 7074 3744 7092 3762
rect 7074 3762 7092 3780
rect 7074 3780 7092 3798
rect 7074 3798 7092 3816
rect 7074 3816 7092 3834
rect 7074 3834 7092 3852
rect 7074 3852 7092 3870
rect 7074 3870 7092 3888
rect 7074 3888 7092 3906
rect 7074 4122 7092 4140
rect 7074 4140 7092 4158
rect 7074 4158 7092 4176
rect 7074 4176 7092 4194
rect 7074 4194 7092 4212
rect 7074 4212 7092 4230
rect 7074 4230 7092 4248
rect 7074 4248 7092 4266
rect 7074 4266 7092 4284
rect 7074 4284 7092 4302
rect 7074 4302 7092 4320
rect 7074 4320 7092 4338
rect 7074 4338 7092 4356
rect 7074 4356 7092 4374
rect 7074 4374 7092 4392
rect 7074 4392 7092 4410
rect 7074 4410 7092 4428
rect 7074 4428 7092 4446
rect 7074 4446 7092 4464
rect 7074 4464 7092 4482
rect 7074 4482 7092 4500
rect 7074 4500 7092 4518
rect 7074 4518 7092 4536
rect 7074 4536 7092 4554
rect 7074 4554 7092 4572
rect 7074 4572 7092 4590
rect 7074 4590 7092 4608
rect 7074 4608 7092 4626
rect 7074 4626 7092 4644
rect 7074 4644 7092 4662
rect 7074 4662 7092 4680
rect 7074 4680 7092 4698
rect 7074 4698 7092 4716
rect 7074 4716 7092 4734
rect 7074 4734 7092 4752
rect 7074 4752 7092 4770
rect 7074 4770 7092 4788
rect 7074 4788 7092 4806
rect 7074 4806 7092 4824
rect 7074 4824 7092 4842
rect 7074 4842 7092 4860
rect 7074 4860 7092 4878
rect 7074 4878 7092 4896
rect 7074 4896 7092 4914
rect 7074 4914 7092 4932
rect 7074 4932 7092 4950
rect 7074 4950 7092 4968
rect 7074 4968 7092 4986
rect 7074 4986 7092 5004
rect 7074 5004 7092 5022
rect 7074 5022 7092 5040
rect 7074 5040 7092 5058
rect 7074 5058 7092 5076
rect 7074 5076 7092 5094
rect 7074 5094 7092 5112
rect 7074 5112 7092 5130
rect 7074 5130 7092 5148
rect 7074 5148 7092 5166
rect 7074 5166 7092 5184
rect 7074 5184 7092 5202
rect 7074 5202 7092 5220
rect 7074 5220 7092 5238
rect 7074 5238 7092 5256
rect 7074 5256 7092 5274
rect 7074 5274 7092 5292
rect 7074 5292 7092 5310
rect 7074 5310 7092 5328
rect 7074 5328 7092 5346
rect 7074 5346 7092 5364
rect 7074 5364 7092 5382
rect 7074 5382 7092 5400
rect 7074 5400 7092 5418
rect 7074 5418 7092 5436
rect 7074 5436 7092 5454
rect 7074 5454 7092 5472
rect 7074 5472 7092 5490
rect 7074 5490 7092 5508
rect 7074 5508 7092 5526
rect 7074 5526 7092 5544
rect 7074 5544 7092 5562
rect 7074 5562 7092 5580
rect 7074 5580 7092 5598
rect 7074 5598 7092 5616
rect 7074 5616 7092 5634
rect 7074 5634 7092 5652
rect 7074 5652 7092 5670
rect 7074 5670 7092 5688
rect 7074 5688 7092 5706
rect 7074 5706 7092 5724
rect 7074 5724 7092 5742
rect 7074 5742 7092 5760
rect 7074 5760 7092 5778
rect 7074 5778 7092 5796
rect 7074 5796 7092 5814
rect 7074 5814 7092 5832
rect 7074 5832 7092 5850
rect 7074 5850 7092 5868
rect 7074 5868 7092 5886
rect 7074 5886 7092 5904
rect 7074 5904 7092 5922
rect 7074 5922 7092 5940
rect 7074 5940 7092 5958
rect 7074 5958 7092 5976
rect 7074 5976 7092 5994
rect 7074 5994 7092 6012
rect 7074 6012 7092 6030
rect 7074 6030 7092 6048
rect 7074 6048 7092 6066
rect 7074 6066 7092 6084
rect 7074 6084 7092 6102
rect 7074 6102 7092 6120
rect 7074 6120 7092 6138
rect 7074 6138 7092 6156
rect 7074 6156 7092 6174
rect 7074 6174 7092 6192
rect 7074 6192 7092 6210
rect 7074 6210 7092 6228
rect 7074 6228 7092 6246
rect 7074 6246 7092 6264
rect 7074 6264 7092 6282
rect 7074 6282 7092 6300
rect 7074 6300 7092 6318
rect 7074 8082 7092 8100
rect 7074 8100 7092 8118
rect 7074 8118 7092 8136
rect 7074 8136 7092 8154
rect 7074 8154 7092 8172
rect 7074 8172 7092 8190
rect 7074 8190 7092 8208
rect 7074 8208 7092 8226
rect 7074 8226 7092 8244
rect 7074 8244 7092 8262
rect 7074 8262 7092 8280
rect 7074 8280 7092 8298
rect 7074 8298 7092 8316
rect 7074 8316 7092 8334
rect 7074 8334 7092 8352
rect 7074 8352 7092 8370
rect 7074 8370 7092 8388
rect 7074 8388 7092 8406
rect 7074 8406 7092 8424
rect 7074 8424 7092 8442
rect 7074 8442 7092 8460
rect 7074 8460 7092 8478
rect 7074 8478 7092 8496
rect 7074 8496 7092 8514
rect 7074 8514 7092 8532
rect 7074 8532 7092 8550
rect 7074 8550 7092 8568
rect 7074 8568 7092 8586
rect 7074 8586 7092 8604
rect 7074 8604 7092 8622
rect 7074 8622 7092 8640
rect 7074 8640 7092 8658
rect 7074 8658 7092 8676
rect 7074 8676 7092 8694
rect 7074 8694 7092 8712
rect 7074 8712 7092 8730
rect 7074 8730 7092 8748
rect 7074 8748 7092 8766
rect 7074 8766 7092 8784
rect 7074 8784 7092 8802
rect 7074 8802 7092 8820
rect 7074 8820 7092 8838
rect 7074 8838 7092 8856
rect 7074 8856 7092 8874
rect 7074 8874 7092 8892
rect 7074 8892 7092 8910
rect 7074 8910 7092 8928
rect 7074 8928 7092 8946
rect 7074 8946 7092 8964
rect 7074 8964 7092 8982
rect 7074 8982 7092 9000
rect 7074 9000 7092 9018
rect 7074 9018 7092 9036
rect 7074 9036 7092 9054
rect 7074 9054 7092 9072
rect 7074 9072 7092 9090
rect 7074 9090 7092 9108
rect 7074 9108 7092 9126
rect 7074 9126 7092 9144
rect 7074 9144 7092 9162
rect 7074 9162 7092 9180
rect 7074 9180 7092 9198
rect 7074 9198 7092 9216
rect 7074 9216 7092 9234
rect 7074 9234 7092 9252
rect 7074 9252 7092 9270
rect 7074 9270 7092 9288
rect 7074 9288 7092 9306
rect 7074 9306 7092 9324
rect 7074 9324 7092 9342
rect 7074 9342 7092 9360
rect 7074 9360 7092 9378
rect 7074 9378 7092 9396
rect 7074 9396 7092 9414
rect 7074 9414 7092 9432
rect 7074 9432 7092 9450
rect 7074 9450 7092 9468
rect 7074 9468 7092 9486
rect 7074 9486 7092 9504
rect 7074 9504 7092 9522
rect 7074 9522 7092 9540
rect 7074 9540 7092 9558
rect 7074 9558 7092 9576
rect 7074 9576 7092 9594
rect 7074 9594 7092 9612
rect 7074 9612 7092 9630
rect 7074 9630 7092 9648
rect 7074 9648 7092 9666
rect 7074 9666 7092 9684
rect 7074 9684 7092 9702
rect 7074 9702 7092 9720
rect 7074 9720 7092 9738
rect 7074 9738 7092 9756
rect 7074 9756 7092 9774
rect 7074 9774 7092 9792
rect 7074 9792 7092 9810
rect 7074 9810 7092 9828
rect 7074 9828 7092 9846
rect 7074 9846 7092 9864
rect 7074 9864 7092 9882
rect 7074 9882 7092 9900
rect 7074 9900 7092 9918
rect 7074 9918 7092 9936
rect 7074 9936 7092 9954
rect 7074 9954 7092 9972
rect 7074 9972 7092 9990
rect 7074 9990 7092 10008
rect 7074 10008 7092 10026
rect 7074 10026 7092 10044
rect 7074 10044 7092 10062
rect 7074 10062 7092 10080
rect 7074 10080 7092 10098
rect 7074 10098 7092 10116
rect 7074 10116 7092 10134
rect 7074 10134 7092 10152
rect 7074 10152 7092 10170
rect 7074 10170 7092 10188
rect 7074 10188 7092 10206
rect 7074 10206 7092 10224
rect 7074 10224 7092 10242
rect 7074 10242 7092 10260
rect 7074 10260 7092 10278
rect 7074 10278 7092 10296
rect 7074 10296 7092 10314
rect 7074 10314 7092 10332
rect 7074 10332 7092 10350
rect 7074 10350 7092 10368
rect 7074 10368 7092 10386
rect 7074 10386 7092 10404
rect 7074 10404 7092 10422
rect 7074 10422 7092 10440
rect 7074 10440 7092 10458
rect 7074 10458 7092 10476
rect 7074 10476 7092 10494
rect 7074 10494 7092 10512
rect 7074 10512 7092 10530
rect 7074 10530 7092 10548
rect 7092 1836 7110 1854
rect 7092 1854 7110 1872
rect 7092 1872 7110 1890
rect 7092 1890 7110 1908
rect 7092 1908 7110 1926
rect 7092 1926 7110 1944
rect 7092 1944 7110 1962
rect 7092 1962 7110 1980
rect 7092 1980 7110 1998
rect 7092 1998 7110 2016
rect 7092 2016 7110 2034
rect 7092 2034 7110 2052
rect 7092 2052 7110 2070
rect 7092 2070 7110 2088
rect 7092 2088 7110 2106
rect 7092 2106 7110 2124
rect 7092 2124 7110 2142
rect 7092 2142 7110 2160
rect 7092 2160 7110 2178
rect 7092 2178 7110 2196
rect 7092 2196 7110 2214
rect 7092 2214 7110 2232
rect 7092 2232 7110 2250
rect 7092 2250 7110 2268
rect 7092 2268 7110 2286
rect 7092 2286 7110 2304
rect 7092 2304 7110 2322
rect 7092 2322 7110 2340
rect 7092 2340 7110 2358
rect 7092 2358 7110 2376
rect 7092 2376 7110 2394
rect 7092 2394 7110 2412
rect 7092 2412 7110 2430
rect 7092 2430 7110 2448
rect 7092 2448 7110 2466
rect 7092 2466 7110 2484
rect 7092 2484 7110 2502
rect 7092 2502 7110 2520
rect 7092 2520 7110 2538
rect 7092 2538 7110 2556
rect 7092 2556 7110 2574
rect 7092 2574 7110 2592
rect 7092 2592 7110 2610
rect 7092 2610 7110 2628
rect 7092 2628 7110 2646
rect 7092 2646 7110 2664
rect 7092 2664 7110 2682
rect 7092 2682 7110 2700
rect 7092 2700 7110 2718
rect 7092 2718 7110 2736
rect 7092 2736 7110 2754
rect 7092 2754 7110 2772
rect 7092 2772 7110 2790
rect 7092 2790 7110 2808
rect 7092 2808 7110 2826
rect 7092 2826 7110 2844
rect 7092 2844 7110 2862
rect 7092 2862 7110 2880
rect 7092 2880 7110 2898
rect 7092 2898 7110 2916
rect 7092 2916 7110 2934
rect 7092 2934 7110 2952
rect 7092 2952 7110 2970
rect 7092 2970 7110 2988
rect 7092 2988 7110 3006
rect 7092 3006 7110 3024
rect 7092 3024 7110 3042
rect 7092 3042 7110 3060
rect 7092 3060 7110 3078
rect 7092 3078 7110 3096
rect 7092 3096 7110 3114
rect 7092 3312 7110 3330
rect 7092 3330 7110 3348
rect 7092 3348 7110 3366
rect 7092 3366 7110 3384
rect 7092 3384 7110 3402
rect 7092 3402 7110 3420
rect 7092 3420 7110 3438
rect 7092 3438 7110 3456
rect 7092 3456 7110 3474
rect 7092 3474 7110 3492
rect 7092 3492 7110 3510
rect 7092 3510 7110 3528
rect 7092 3528 7110 3546
rect 7092 3546 7110 3564
rect 7092 3564 7110 3582
rect 7092 3582 7110 3600
rect 7092 3600 7110 3618
rect 7092 3618 7110 3636
rect 7092 3636 7110 3654
rect 7092 3654 7110 3672
rect 7092 3672 7110 3690
rect 7092 3690 7110 3708
rect 7092 3708 7110 3726
rect 7092 3726 7110 3744
rect 7092 3744 7110 3762
rect 7092 3762 7110 3780
rect 7092 3780 7110 3798
rect 7092 3798 7110 3816
rect 7092 3816 7110 3834
rect 7092 3834 7110 3852
rect 7092 3852 7110 3870
rect 7092 3870 7110 3888
rect 7092 3888 7110 3906
rect 7092 3906 7110 3924
rect 7092 4140 7110 4158
rect 7092 4158 7110 4176
rect 7092 4176 7110 4194
rect 7092 4194 7110 4212
rect 7092 4212 7110 4230
rect 7092 4230 7110 4248
rect 7092 4248 7110 4266
rect 7092 4266 7110 4284
rect 7092 4284 7110 4302
rect 7092 4302 7110 4320
rect 7092 4320 7110 4338
rect 7092 4338 7110 4356
rect 7092 4356 7110 4374
rect 7092 4374 7110 4392
rect 7092 4392 7110 4410
rect 7092 4410 7110 4428
rect 7092 4428 7110 4446
rect 7092 4446 7110 4464
rect 7092 4464 7110 4482
rect 7092 4482 7110 4500
rect 7092 4500 7110 4518
rect 7092 4518 7110 4536
rect 7092 4536 7110 4554
rect 7092 4554 7110 4572
rect 7092 4572 7110 4590
rect 7092 4590 7110 4608
rect 7092 4608 7110 4626
rect 7092 4626 7110 4644
rect 7092 4644 7110 4662
rect 7092 4662 7110 4680
rect 7092 4680 7110 4698
rect 7092 4698 7110 4716
rect 7092 4716 7110 4734
rect 7092 4734 7110 4752
rect 7092 4752 7110 4770
rect 7092 4770 7110 4788
rect 7092 4788 7110 4806
rect 7092 4806 7110 4824
rect 7092 4824 7110 4842
rect 7092 4842 7110 4860
rect 7092 4860 7110 4878
rect 7092 4878 7110 4896
rect 7092 4896 7110 4914
rect 7092 4914 7110 4932
rect 7092 4932 7110 4950
rect 7092 4950 7110 4968
rect 7092 4968 7110 4986
rect 7092 4986 7110 5004
rect 7092 5004 7110 5022
rect 7092 5022 7110 5040
rect 7092 5040 7110 5058
rect 7092 5058 7110 5076
rect 7092 5076 7110 5094
rect 7092 5094 7110 5112
rect 7092 5112 7110 5130
rect 7092 5130 7110 5148
rect 7092 5148 7110 5166
rect 7092 5166 7110 5184
rect 7092 5184 7110 5202
rect 7092 5202 7110 5220
rect 7092 5220 7110 5238
rect 7092 5238 7110 5256
rect 7092 5256 7110 5274
rect 7092 5274 7110 5292
rect 7092 5292 7110 5310
rect 7092 5310 7110 5328
rect 7092 5328 7110 5346
rect 7092 5346 7110 5364
rect 7092 5364 7110 5382
rect 7092 5382 7110 5400
rect 7092 5400 7110 5418
rect 7092 5418 7110 5436
rect 7092 5436 7110 5454
rect 7092 5454 7110 5472
rect 7092 5472 7110 5490
rect 7092 5490 7110 5508
rect 7092 5508 7110 5526
rect 7092 5526 7110 5544
rect 7092 5544 7110 5562
rect 7092 5562 7110 5580
rect 7092 5580 7110 5598
rect 7092 5598 7110 5616
rect 7092 5616 7110 5634
rect 7092 5634 7110 5652
rect 7092 5652 7110 5670
rect 7092 5670 7110 5688
rect 7092 5688 7110 5706
rect 7092 5706 7110 5724
rect 7092 5724 7110 5742
rect 7092 5742 7110 5760
rect 7092 5760 7110 5778
rect 7092 5778 7110 5796
rect 7092 5796 7110 5814
rect 7092 5814 7110 5832
rect 7092 5832 7110 5850
rect 7092 5850 7110 5868
rect 7092 5868 7110 5886
rect 7092 5886 7110 5904
rect 7092 5904 7110 5922
rect 7092 5922 7110 5940
rect 7092 5940 7110 5958
rect 7092 5958 7110 5976
rect 7092 5976 7110 5994
rect 7092 5994 7110 6012
rect 7092 6012 7110 6030
rect 7092 6030 7110 6048
rect 7092 6048 7110 6066
rect 7092 6066 7110 6084
rect 7092 6084 7110 6102
rect 7092 6102 7110 6120
rect 7092 6120 7110 6138
rect 7092 6138 7110 6156
rect 7092 6156 7110 6174
rect 7092 6174 7110 6192
rect 7092 6192 7110 6210
rect 7092 6210 7110 6228
rect 7092 6228 7110 6246
rect 7092 6246 7110 6264
rect 7092 6264 7110 6282
rect 7092 6282 7110 6300
rect 7092 6300 7110 6318
rect 7092 6318 7110 6336
rect 7092 8136 7110 8154
rect 7092 8154 7110 8172
rect 7092 8172 7110 8190
rect 7092 8190 7110 8208
rect 7092 8208 7110 8226
rect 7092 8226 7110 8244
rect 7092 8244 7110 8262
rect 7092 8262 7110 8280
rect 7092 8280 7110 8298
rect 7092 8298 7110 8316
rect 7092 8316 7110 8334
rect 7092 8334 7110 8352
rect 7092 8352 7110 8370
rect 7092 8370 7110 8388
rect 7092 8388 7110 8406
rect 7092 8406 7110 8424
rect 7092 8424 7110 8442
rect 7092 8442 7110 8460
rect 7092 8460 7110 8478
rect 7092 8478 7110 8496
rect 7092 8496 7110 8514
rect 7092 8514 7110 8532
rect 7092 8532 7110 8550
rect 7092 8550 7110 8568
rect 7092 8568 7110 8586
rect 7092 8586 7110 8604
rect 7092 8604 7110 8622
rect 7092 8622 7110 8640
rect 7092 8640 7110 8658
rect 7092 8658 7110 8676
rect 7092 8676 7110 8694
rect 7092 8694 7110 8712
rect 7092 8712 7110 8730
rect 7092 8730 7110 8748
rect 7092 8748 7110 8766
rect 7092 8766 7110 8784
rect 7092 8784 7110 8802
rect 7092 8802 7110 8820
rect 7092 8820 7110 8838
rect 7092 8838 7110 8856
rect 7092 8856 7110 8874
rect 7092 8874 7110 8892
rect 7092 8892 7110 8910
rect 7092 8910 7110 8928
rect 7092 8928 7110 8946
rect 7092 8946 7110 8964
rect 7092 8964 7110 8982
rect 7092 8982 7110 9000
rect 7092 9000 7110 9018
rect 7092 9018 7110 9036
rect 7092 9036 7110 9054
rect 7092 9054 7110 9072
rect 7092 9072 7110 9090
rect 7092 9090 7110 9108
rect 7092 9108 7110 9126
rect 7092 9126 7110 9144
rect 7092 9144 7110 9162
rect 7092 9162 7110 9180
rect 7092 9180 7110 9198
rect 7092 9198 7110 9216
rect 7092 9216 7110 9234
rect 7092 9234 7110 9252
rect 7092 9252 7110 9270
rect 7092 9270 7110 9288
rect 7092 9288 7110 9306
rect 7092 9306 7110 9324
rect 7092 9324 7110 9342
rect 7092 9342 7110 9360
rect 7092 9360 7110 9378
rect 7092 9378 7110 9396
rect 7092 9396 7110 9414
rect 7092 9414 7110 9432
rect 7092 9432 7110 9450
rect 7092 9450 7110 9468
rect 7092 9468 7110 9486
rect 7092 9486 7110 9504
rect 7092 9504 7110 9522
rect 7092 9522 7110 9540
rect 7092 9540 7110 9558
rect 7092 9558 7110 9576
rect 7092 9576 7110 9594
rect 7092 9594 7110 9612
rect 7092 9612 7110 9630
rect 7092 9630 7110 9648
rect 7092 9648 7110 9666
rect 7092 9666 7110 9684
rect 7092 9684 7110 9702
rect 7092 9702 7110 9720
rect 7092 9720 7110 9738
rect 7092 9738 7110 9756
rect 7092 9756 7110 9774
rect 7092 9774 7110 9792
rect 7092 9792 7110 9810
rect 7092 9810 7110 9828
rect 7092 9828 7110 9846
rect 7092 9846 7110 9864
rect 7092 9864 7110 9882
rect 7092 9882 7110 9900
rect 7092 9900 7110 9918
rect 7092 9918 7110 9936
rect 7092 9936 7110 9954
rect 7092 9954 7110 9972
rect 7092 9972 7110 9990
rect 7092 9990 7110 10008
rect 7092 10008 7110 10026
rect 7092 10026 7110 10044
rect 7092 10044 7110 10062
rect 7092 10062 7110 10080
rect 7092 10080 7110 10098
rect 7092 10098 7110 10116
rect 7092 10116 7110 10134
rect 7092 10134 7110 10152
rect 7092 10152 7110 10170
rect 7092 10170 7110 10188
rect 7092 10188 7110 10206
rect 7092 10206 7110 10224
rect 7092 10224 7110 10242
rect 7092 10242 7110 10260
rect 7092 10260 7110 10278
rect 7092 10278 7110 10296
rect 7092 10296 7110 10314
rect 7092 10314 7110 10332
rect 7092 10332 7110 10350
rect 7092 10350 7110 10368
rect 7092 10368 7110 10386
rect 7092 10386 7110 10404
rect 7092 10404 7110 10422
rect 7092 10422 7110 10440
rect 7092 10440 7110 10458
rect 7092 10458 7110 10476
rect 7110 1854 7128 1872
rect 7110 1872 7128 1890
rect 7110 1890 7128 1908
rect 7110 1908 7128 1926
rect 7110 1926 7128 1944
rect 7110 1944 7128 1962
rect 7110 1962 7128 1980
rect 7110 1980 7128 1998
rect 7110 1998 7128 2016
rect 7110 2016 7128 2034
rect 7110 2034 7128 2052
rect 7110 2052 7128 2070
rect 7110 2070 7128 2088
rect 7110 2088 7128 2106
rect 7110 2106 7128 2124
rect 7110 2124 7128 2142
rect 7110 2142 7128 2160
rect 7110 2160 7128 2178
rect 7110 2178 7128 2196
rect 7110 2196 7128 2214
rect 7110 2214 7128 2232
rect 7110 2232 7128 2250
rect 7110 2250 7128 2268
rect 7110 2268 7128 2286
rect 7110 2286 7128 2304
rect 7110 2304 7128 2322
rect 7110 2322 7128 2340
rect 7110 2340 7128 2358
rect 7110 2358 7128 2376
rect 7110 2376 7128 2394
rect 7110 2394 7128 2412
rect 7110 2412 7128 2430
rect 7110 2430 7128 2448
rect 7110 2448 7128 2466
rect 7110 2466 7128 2484
rect 7110 2484 7128 2502
rect 7110 2502 7128 2520
rect 7110 2520 7128 2538
rect 7110 2538 7128 2556
rect 7110 2556 7128 2574
rect 7110 2574 7128 2592
rect 7110 2592 7128 2610
rect 7110 2610 7128 2628
rect 7110 2628 7128 2646
rect 7110 2646 7128 2664
rect 7110 2664 7128 2682
rect 7110 2682 7128 2700
rect 7110 2700 7128 2718
rect 7110 2718 7128 2736
rect 7110 2736 7128 2754
rect 7110 2754 7128 2772
rect 7110 2772 7128 2790
rect 7110 2790 7128 2808
rect 7110 2808 7128 2826
rect 7110 2826 7128 2844
rect 7110 2844 7128 2862
rect 7110 2862 7128 2880
rect 7110 2880 7128 2898
rect 7110 2898 7128 2916
rect 7110 2916 7128 2934
rect 7110 2934 7128 2952
rect 7110 2952 7128 2970
rect 7110 2970 7128 2988
rect 7110 2988 7128 3006
rect 7110 3006 7128 3024
rect 7110 3024 7128 3042
rect 7110 3042 7128 3060
rect 7110 3060 7128 3078
rect 7110 3078 7128 3096
rect 7110 3096 7128 3114
rect 7110 3114 7128 3132
rect 7110 3312 7128 3330
rect 7110 3330 7128 3348
rect 7110 3348 7128 3366
rect 7110 3366 7128 3384
rect 7110 3384 7128 3402
rect 7110 3402 7128 3420
rect 7110 3420 7128 3438
rect 7110 3438 7128 3456
rect 7110 3456 7128 3474
rect 7110 3474 7128 3492
rect 7110 3492 7128 3510
rect 7110 3510 7128 3528
rect 7110 3528 7128 3546
rect 7110 3546 7128 3564
rect 7110 3564 7128 3582
rect 7110 3582 7128 3600
rect 7110 3600 7128 3618
rect 7110 3618 7128 3636
rect 7110 3636 7128 3654
rect 7110 3654 7128 3672
rect 7110 3672 7128 3690
rect 7110 3690 7128 3708
rect 7110 3708 7128 3726
rect 7110 3726 7128 3744
rect 7110 3744 7128 3762
rect 7110 3762 7128 3780
rect 7110 3780 7128 3798
rect 7110 3798 7128 3816
rect 7110 3816 7128 3834
rect 7110 3834 7128 3852
rect 7110 3852 7128 3870
rect 7110 3870 7128 3888
rect 7110 3888 7128 3906
rect 7110 3906 7128 3924
rect 7110 3924 7128 3942
rect 7110 4158 7128 4176
rect 7110 4176 7128 4194
rect 7110 4194 7128 4212
rect 7110 4212 7128 4230
rect 7110 4230 7128 4248
rect 7110 4248 7128 4266
rect 7110 4266 7128 4284
rect 7110 4284 7128 4302
rect 7110 4302 7128 4320
rect 7110 4320 7128 4338
rect 7110 4338 7128 4356
rect 7110 4356 7128 4374
rect 7110 4374 7128 4392
rect 7110 4392 7128 4410
rect 7110 4410 7128 4428
rect 7110 4428 7128 4446
rect 7110 4446 7128 4464
rect 7110 4464 7128 4482
rect 7110 4482 7128 4500
rect 7110 4500 7128 4518
rect 7110 4518 7128 4536
rect 7110 4536 7128 4554
rect 7110 4554 7128 4572
rect 7110 4572 7128 4590
rect 7110 4590 7128 4608
rect 7110 4608 7128 4626
rect 7110 4626 7128 4644
rect 7110 4644 7128 4662
rect 7110 4662 7128 4680
rect 7110 4680 7128 4698
rect 7110 4698 7128 4716
rect 7110 4716 7128 4734
rect 7110 4734 7128 4752
rect 7110 4752 7128 4770
rect 7110 4770 7128 4788
rect 7110 4788 7128 4806
rect 7110 4806 7128 4824
rect 7110 4824 7128 4842
rect 7110 4842 7128 4860
rect 7110 4860 7128 4878
rect 7110 4878 7128 4896
rect 7110 4896 7128 4914
rect 7110 4914 7128 4932
rect 7110 4932 7128 4950
rect 7110 4950 7128 4968
rect 7110 4968 7128 4986
rect 7110 4986 7128 5004
rect 7110 5004 7128 5022
rect 7110 5022 7128 5040
rect 7110 5040 7128 5058
rect 7110 5058 7128 5076
rect 7110 5076 7128 5094
rect 7110 5094 7128 5112
rect 7110 5112 7128 5130
rect 7110 5130 7128 5148
rect 7110 5148 7128 5166
rect 7110 5166 7128 5184
rect 7110 5184 7128 5202
rect 7110 5202 7128 5220
rect 7110 5220 7128 5238
rect 7110 5238 7128 5256
rect 7110 5256 7128 5274
rect 7110 5274 7128 5292
rect 7110 5292 7128 5310
rect 7110 5310 7128 5328
rect 7110 5328 7128 5346
rect 7110 5346 7128 5364
rect 7110 5364 7128 5382
rect 7110 5382 7128 5400
rect 7110 5400 7128 5418
rect 7110 5418 7128 5436
rect 7110 5436 7128 5454
rect 7110 5454 7128 5472
rect 7110 5472 7128 5490
rect 7110 5490 7128 5508
rect 7110 5508 7128 5526
rect 7110 5526 7128 5544
rect 7110 5544 7128 5562
rect 7110 5562 7128 5580
rect 7110 5580 7128 5598
rect 7110 5598 7128 5616
rect 7110 5616 7128 5634
rect 7110 5634 7128 5652
rect 7110 5652 7128 5670
rect 7110 5670 7128 5688
rect 7110 5688 7128 5706
rect 7110 5706 7128 5724
rect 7110 5724 7128 5742
rect 7110 5742 7128 5760
rect 7110 5760 7128 5778
rect 7110 5778 7128 5796
rect 7110 5796 7128 5814
rect 7110 5814 7128 5832
rect 7110 5832 7128 5850
rect 7110 5850 7128 5868
rect 7110 5868 7128 5886
rect 7110 5886 7128 5904
rect 7110 5904 7128 5922
rect 7110 5922 7128 5940
rect 7110 5940 7128 5958
rect 7110 5958 7128 5976
rect 7110 5976 7128 5994
rect 7110 5994 7128 6012
rect 7110 6012 7128 6030
rect 7110 6030 7128 6048
rect 7110 6048 7128 6066
rect 7110 6066 7128 6084
rect 7110 6084 7128 6102
rect 7110 6102 7128 6120
rect 7110 6120 7128 6138
rect 7110 6138 7128 6156
rect 7110 6156 7128 6174
rect 7110 6174 7128 6192
rect 7110 6192 7128 6210
rect 7110 6210 7128 6228
rect 7110 6228 7128 6246
rect 7110 6246 7128 6264
rect 7110 6264 7128 6282
rect 7110 6282 7128 6300
rect 7110 6300 7128 6318
rect 7110 6318 7128 6336
rect 7110 6336 7128 6354
rect 7110 8190 7128 8208
rect 7110 8208 7128 8226
rect 7110 8226 7128 8244
rect 7110 8244 7128 8262
rect 7110 8262 7128 8280
rect 7110 8280 7128 8298
rect 7110 8298 7128 8316
rect 7110 8316 7128 8334
rect 7110 8334 7128 8352
rect 7110 8352 7128 8370
rect 7110 8370 7128 8388
rect 7110 8388 7128 8406
rect 7110 8406 7128 8424
rect 7110 8424 7128 8442
rect 7110 8442 7128 8460
rect 7110 8460 7128 8478
rect 7110 8478 7128 8496
rect 7110 8496 7128 8514
rect 7110 8514 7128 8532
rect 7110 8532 7128 8550
rect 7110 8550 7128 8568
rect 7110 8568 7128 8586
rect 7110 8586 7128 8604
rect 7110 8604 7128 8622
rect 7110 8622 7128 8640
rect 7110 8640 7128 8658
rect 7110 8658 7128 8676
rect 7110 8676 7128 8694
rect 7110 8694 7128 8712
rect 7110 8712 7128 8730
rect 7110 8730 7128 8748
rect 7110 8748 7128 8766
rect 7110 8766 7128 8784
rect 7110 8784 7128 8802
rect 7110 8802 7128 8820
rect 7110 8820 7128 8838
rect 7110 8838 7128 8856
rect 7110 8856 7128 8874
rect 7110 8874 7128 8892
rect 7110 8892 7128 8910
rect 7110 8910 7128 8928
rect 7110 8928 7128 8946
rect 7110 8946 7128 8964
rect 7110 8964 7128 8982
rect 7110 8982 7128 9000
rect 7110 9000 7128 9018
rect 7110 9018 7128 9036
rect 7110 9036 7128 9054
rect 7110 9054 7128 9072
rect 7110 9072 7128 9090
rect 7110 9090 7128 9108
rect 7110 9108 7128 9126
rect 7110 9126 7128 9144
rect 7110 9144 7128 9162
rect 7110 9162 7128 9180
rect 7110 9180 7128 9198
rect 7110 9198 7128 9216
rect 7110 9216 7128 9234
rect 7110 9234 7128 9252
rect 7110 9252 7128 9270
rect 7110 9270 7128 9288
rect 7110 9288 7128 9306
rect 7110 9306 7128 9324
rect 7110 9324 7128 9342
rect 7110 9342 7128 9360
rect 7110 9360 7128 9378
rect 7110 9378 7128 9396
rect 7110 9396 7128 9414
rect 7110 9414 7128 9432
rect 7110 9432 7128 9450
rect 7110 9450 7128 9468
rect 7110 9468 7128 9486
rect 7110 9486 7128 9504
rect 7110 9504 7128 9522
rect 7110 9522 7128 9540
rect 7110 9540 7128 9558
rect 7110 9558 7128 9576
rect 7110 9576 7128 9594
rect 7110 9594 7128 9612
rect 7110 9612 7128 9630
rect 7110 9630 7128 9648
rect 7110 9648 7128 9666
rect 7110 9666 7128 9684
rect 7110 9684 7128 9702
rect 7110 9702 7128 9720
rect 7110 9720 7128 9738
rect 7110 9738 7128 9756
rect 7110 9756 7128 9774
rect 7110 9774 7128 9792
rect 7110 9792 7128 9810
rect 7110 9810 7128 9828
rect 7110 9828 7128 9846
rect 7110 9846 7128 9864
rect 7110 9864 7128 9882
rect 7110 9882 7128 9900
rect 7110 9900 7128 9918
rect 7110 9918 7128 9936
rect 7110 9936 7128 9954
rect 7110 9954 7128 9972
rect 7110 9972 7128 9990
rect 7110 9990 7128 10008
rect 7110 10008 7128 10026
rect 7110 10026 7128 10044
rect 7110 10044 7128 10062
rect 7110 10062 7128 10080
rect 7110 10080 7128 10098
rect 7110 10098 7128 10116
rect 7110 10116 7128 10134
rect 7110 10134 7128 10152
rect 7110 10152 7128 10170
rect 7110 10170 7128 10188
rect 7110 10188 7128 10206
rect 7110 10206 7128 10224
rect 7110 10224 7128 10242
rect 7110 10242 7128 10260
rect 7110 10260 7128 10278
rect 7110 10278 7128 10296
rect 7110 10296 7128 10314
rect 7110 10314 7128 10332
rect 7110 10332 7128 10350
rect 7110 10350 7128 10368
rect 7110 10368 7128 10386
rect 7110 10386 7128 10404
rect 7128 1872 7146 1890
rect 7128 1890 7146 1908
rect 7128 1908 7146 1926
rect 7128 1926 7146 1944
rect 7128 1944 7146 1962
rect 7128 1962 7146 1980
rect 7128 1980 7146 1998
rect 7128 1998 7146 2016
rect 7128 2016 7146 2034
rect 7128 2034 7146 2052
rect 7128 2052 7146 2070
rect 7128 2070 7146 2088
rect 7128 2088 7146 2106
rect 7128 2106 7146 2124
rect 7128 2124 7146 2142
rect 7128 2142 7146 2160
rect 7128 2160 7146 2178
rect 7128 2178 7146 2196
rect 7128 2196 7146 2214
rect 7128 2214 7146 2232
rect 7128 2232 7146 2250
rect 7128 2250 7146 2268
rect 7128 2268 7146 2286
rect 7128 2286 7146 2304
rect 7128 2304 7146 2322
rect 7128 2322 7146 2340
rect 7128 2340 7146 2358
rect 7128 2358 7146 2376
rect 7128 2376 7146 2394
rect 7128 2394 7146 2412
rect 7128 2412 7146 2430
rect 7128 2430 7146 2448
rect 7128 2448 7146 2466
rect 7128 2466 7146 2484
rect 7128 2484 7146 2502
rect 7128 2502 7146 2520
rect 7128 2520 7146 2538
rect 7128 2538 7146 2556
rect 7128 2556 7146 2574
rect 7128 2574 7146 2592
rect 7128 2592 7146 2610
rect 7128 2610 7146 2628
rect 7128 2628 7146 2646
rect 7128 2646 7146 2664
rect 7128 2664 7146 2682
rect 7128 2682 7146 2700
rect 7128 2700 7146 2718
rect 7128 2718 7146 2736
rect 7128 2736 7146 2754
rect 7128 2754 7146 2772
rect 7128 2772 7146 2790
rect 7128 2790 7146 2808
rect 7128 2808 7146 2826
rect 7128 2826 7146 2844
rect 7128 2844 7146 2862
rect 7128 2862 7146 2880
rect 7128 2880 7146 2898
rect 7128 2898 7146 2916
rect 7128 2916 7146 2934
rect 7128 2934 7146 2952
rect 7128 2952 7146 2970
rect 7128 2970 7146 2988
rect 7128 2988 7146 3006
rect 7128 3006 7146 3024
rect 7128 3024 7146 3042
rect 7128 3042 7146 3060
rect 7128 3060 7146 3078
rect 7128 3078 7146 3096
rect 7128 3096 7146 3114
rect 7128 3114 7146 3132
rect 7128 3312 7146 3330
rect 7128 3330 7146 3348
rect 7128 3348 7146 3366
rect 7128 3366 7146 3384
rect 7128 3384 7146 3402
rect 7128 3402 7146 3420
rect 7128 3420 7146 3438
rect 7128 3438 7146 3456
rect 7128 3456 7146 3474
rect 7128 3474 7146 3492
rect 7128 3492 7146 3510
rect 7128 3510 7146 3528
rect 7128 3528 7146 3546
rect 7128 3546 7146 3564
rect 7128 3564 7146 3582
rect 7128 3582 7146 3600
rect 7128 3600 7146 3618
rect 7128 3618 7146 3636
rect 7128 3636 7146 3654
rect 7128 3654 7146 3672
rect 7128 3672 7146 3690
rect 7128 3690 7146 3708
rect 7128 3708 7146 3726
rect 7128 3726 7146 3744
rect 7128 3744 7146 3762
rect 7128 3762 7146 3780
rect 7128 3780 7146 3798
rect 7128 3798 7146 3816
rect 7128 3816 7146 3834
rect 7128 3834 7146 3852
rect 7128 3852 7146 3870
rect 7128 3870 7146 3888
rect 7128 3888 7146 3906
rect 7128 3906 7146 3924
rect 7128 3924 7146 3942
rect 7128 3942 7146 3960
rect 7128 4176 7146 4194
rect 7128 4194 7146 4212
rect 7128 4212 7146 4230
rect 7128 4230 7146 4248
rect 7128 4248 7146 4266
rect 7128 4266 7146 4284
rect 7128 4284 7146 4302
rect 7128 4302 7146 4320
rect 7128 4320 7146 4338
rect 7128 4338 7146 4356
rect 7128 4356 7146 4374
rect 7128 4374 7146 4392
rect 7128 4392 7146 4410
rect 7128 4410 7146 4428
rect 7128 4428 7146 4446
rect 7128 4446 7146 4464
rect 7128 4464 7146 4482
rect 7128 4482 7146 4500
rect 7128 4500 7146 4518
rect 7128 4518 7146 4536
rect 7128 4536 7146 4554
rect 7128 4554 7146 4572
rect 7128 4572 7146 4590
rect 7128 4590 7146 4608
rect 7128 4608 7146 4626
rect 7128 4626 7146 4644
rect 7128 4644 7146 4662
rect 7128 4662 7146 4680
rect 7128 4680 7146 4698
rect 7128 4698 7146 4716
rect 7128 4716 7146 4734
rect 7128 4734 7146 4752
rect 7128 4752 7146 4770
rect 7128 4770 7146 4788
rect 7128 4788 7146 4806
rect 7128 4806 7146 4824
rect 7128 4824 7146 4842
rect 7128 4842 7146 4860
rect 7128 4860 7146 4878
rect 7128 4878 7146 4896
rect 7128 4896 7146 4914
rect 7128 4914 7146 4932
rect 7128 4932 7146 4950
rect 7128 4950 7146 4968
rect 7128 4968 7146 4986
rect 7128 4986 7146 5004
rect 7128 5004 7146 5022
rect 7128 5022 7146 5040
rect 7128 5040 7146 5058
rect 7128 5058 7146 5076
rect 7128 5076 7146 5094
rect 7128 5094 7146 5112
rect 7128 5112 7146 5130
rect 7128 5130 7146 5148
rect 7128 5148 7146 5166
rect 7128 5166 7146 5184
rect 7128 5184 7146 5202
rect 7128 5202 7146 5220
rect 7128 5220 7146 5238
rect 7128 5238 7146 5256
rect 7128 5256 7146 5274
rect 7128 5274 7146 5292
rect 7128 5292 7146 5310
rect 7128 5310 7146 5328
rect 7128 5328 7146 5346
rect 7128 5346 7146 5364
rect 7128 5364 7146 5382
rect 7128 5382 7146 5400
rect 7128 5400 7146 5418
rect 7128 5418 7146 5436
rect 7128 5436 7146 5454
rect 7128 5454 7146 5472
rect 7128 5472 7146 5490
rect 7128 5490 7146 5508
rect 7128 5508 7146 5526
rect 7128 5526 7146 5544
rect 7128 5544 7146 5562
rect 7128 5562 7146 5580
rect 7128 5580 7146 5598
rect 7128 5598 7146 5616
rect 7128 5616 7146 5634
rect 7128 5634 7146 5652
rect 7128 5652 7146 5670
rect 7128 5670 7146 5688
rect 7128 5688 7146 5706
rect 7128 5706 7146 5724
rect 7128 5724 7146 5742
rect 7128 5742 7146 5760
rect 7128 5760 7146 5778
rect 7128 5778 7146 5796
rect 7128 5796 7146 5814
rect 7128 5814 7146 5832
rect 7128 5832 7146 5850
rect 7128 5850 7146 5868
rect 7128 5868 7146 5886
rect 7128 5886 7146 5904
rect 7128 5904 7146 5922
rect 7128 5922 7146 5940
rect 7128 5940 7146 5958
rect 7128 5958 7146 5976
rect 7128 5976 7146 5994
rect 7128 5994 7146 6012
rect 7128 6012 7146 6030
rect 7128 6030 7146 6048
rect 7128 6048 7146 6066
rect 7128 6066 7146 6084
rect 7128 6084 7146 6102
rect 7128 6102 7146 6120
rect 7128 6120 7146 6138
rect 7128 6138 7146 6156
rect 7128 6156 7146 6174
rect 7128 6174 7146 6192
rect 7128 6192 7146 6210
rect 7128 6210 7146 6228
rect 7128 6228 7146 6246
rect 7128 6246 7146 6264
rect 7128 6264 7146 6282
rect 7128 6282 7146 6300
rect 7128 6300 7146 6318
rect 7128 6318 7146 6336
rect 7128 6336 7146 6354
rect 7128 6354 7146 6372
rect 7128 8244 7146 8262
rect 7128 8262 7146 8280
rect 7128 8280 7146 8298
rect 7128 8298 7146 8316
rect 7128 8316 7146 8334
rect 7128 8334 7146 8352
rect 7128 8352 7146 8370
rect 7128 8370 7146 8388
rect 7128 8388 7146 8406
rect 7128 8406 7146 8424
rect 7128 8424 7146 8442
rect 7128 8442 7146 8460
rect 7128 8460 7146 8478
rect 7128 8478 7146 8496
rect 7128 8496 7146 8514
rect 7128 8514 7146 8532
rect 7128 8532 7146 8550
rect 7128 8550 7146 8568
rect 7128 8568 7146 8586
rect 7128 8586 7146 8604
rect 7128 8604 7146 8622
rect 7128 8622 7146 8640
rect 7128 8640 7146 8658
rect 7128 8658 7146 8676
rect 7128 8676 7146 8694
rect 7128 8694 7146 8712
rect 7128 8712 7146 8730
rect 7128 8730 7146 8748
rect 7128 8748 7146 8766
rect 7128 8766 7146 8784
rect 7128 8784 7146 8802
rect 7128 8802 7146 8820
rect 7128 8820 7146 8838
rect 7128 8838 7146 8856
rect 7128 8856 7146 8874
rect 7128 8874 7146 8892
rect 7128 8892 7146 8910
rect 7128 8910 7146 8928
rect 7128 8928 7146 8946
rect 7128 8946 7146 8964
rect 7128 8964 7146 8982
rect 7128 8982 7146 9000
rect 7128 9000 7146 9018
rect 7128 9018 7146 9036
rect 7128 9036 7146 9054
rect 7128 9054 7146 9072
rect 7128 9072 7146 9090
rect 7128 9090 7146 9108
rect 7128 9108 7146 9126
rect 7128 9126 7146 9144
rect 7128 9144 7146 9162
rect 7128 9162 7146 9180
rect 7128 9180 7146 9198
rect 7128 9198 7146 9216
rect 7128 9216 7146 9234
rect 7128 9234 7146 9252
rect 7128 9252 7146 9270
rect 7128 9270 7146 9288
rect 7128 9288 7146 9306
rect 7128 9306 7146 9324
rect 7128 9324 7146 9342
rect 7128 9342 7146 9360
rect 7128 9360 7146 9378
rect 7128 9378 7146 9396
rect 7128 9396 7146 9414
rect 7128 9414 7146 9432
rect 7128 9432 7146 9450
rect 7128 9450 7146 9468
rect 7128 9468 7146 9486
rect 7128 9486 7146 9504
rect 7128 9504 7146 9522
rect 7128 9522 7146 9540
rect 7128 9540 7146 9558
rect 7128 9558 7146 9576
rect 7128 9576 7146 9594
rect 7128 9594 7146 9612
rect 7128 9612 7146 9630
rect 7128 9630 7146 9648
rect 7128 9648 7146 9666
rect 7128 9666 7146 9684
rect 7128 9684 7146 9702
rect 7128 9702 7146 9720
rect 7128 9720 7146 9738
rect 7128 9738 7146 9756
rect 7128 9756 7146 9774
rect 7128 9774 7146 9792
rect 7128 9792 7146 9810
rect 7128 9810 7146 9828
rect 7128 9828 7146 9846
rect 7128 9846 7146 9864
rect 7128 9864 7146 9882
rect 7128 9882 7146 9900
rect 7128 9900 7146 9918
rect 7128 9918 7146 9936
rect 7128 9936 7146 9954
rect 7128 9954 7146 9972
rect 7128 9972 7146 9990
rect 7128 9990 7146 10008
rect 7128 10008 7146 10026
rect 7128 10026 7146 10044
rect 7128 10044 7146 10062
rect 7128 10062 7146 10080
rect 7128 10080 7146 10098
rect 7128 10098 7146 10116
rect 7128 10116 7146 10134
rect 7128 10134 7146 10152
rect 7128 10152 7146 10170
rect 7128 10170 7146 10188
rect 7128 10188 7146 10206
rect 7128 10206 7146 10224
rect 7128 10224 7146 10242
rect 7128 10242 7146 10260
rect 7128 10260 7146 10278
rect 7128 10278 7146 10296
rect 7128 10296 7146 10314
rect 7128 10314 7146 10332
rect 7128 10332 7146 10350
rect 7146 1872 7164 1890
rect 7146 1890 7164 1908
rect 7146 1908 7164 1926
rect 7146 1926 7164 1944
rect 7146 1944 7164 1962
rect 7146 1962 7164 1980
rect 7146 1980 7164 1998
rect 7146 1998 7164 2016
rect 7146 2016 7164 2034
rect 7146 2034 7164 2052
rect 7146 2052 7164 2070
rect 7146 2070 7164 2088
rect 7146 2088 7164 2106
rect 7146 2106 7164 2124
rect 7146 2124 7164 2142
rect 7146 2142 7164 2160
rect 7146 2160 7164 2178
rect 7146 2178 7164 2196
rect 7146 2196 7164 2214
rect 7146 2214 7164 2232
rect 7146 2232 7164 2250
rect 7146 2250 7164 2268
rect 7146 2268 7164 2286
rect 7146 2286 7164 2304
rect 7146 2304 7164 2322
rect 7146 2322 7164 2340
rect 7146 2340 7164 2358
rect 7146 2358 7164 2376
rect 7146 2376 7164 2394
rect 7146 2394 7164 2412
rect 7146 2412 7164 2430
rect 7146 2430 7164 2448
rect 7146 2448 7164 2466
rect 7146 2466 7164 2484
rect 7146 2484 7164 2502
rect 7146 2502 7164 2520
rect 7146 2520 7164 2538
rect 7146 2538 7164 2556
rect 7146 2556 7164 2574
rect 7146 2574 7164 2592
rect 7146 2592 7164 2610
rect 7146 2610 7164 2628
rect 7146 2628 7164 2646
rect 7146 2646 7164 2664
rect 7146 2664 7164 2682
rect 7146 2682 7164 2700
rect 7146 2700 7164 2718
rect 7146 2718 7164 2736
rect 7146 2736 7164 2754
rect 7146 2754 7164 2772
rect 7146 2772 7164 2790
rect 7146 2790 7164 2808
rect 7146 2808 7164 2826
rect 7146 2826 7164 2844
rect 7146 2844 7164 2862
rect 7146 2862 7164 2880
rect 7146 2880 7164 2898
rect 7146 2898 7164 2916
rect 7146 2916 7164 2934
rect 7146 2934 7164 2952
rect 7146 2952 7164 2970
rect 7146 2970 7164 2988
rect 7146 2988 7164 3006
rect 7146 3006 7164 3024
rect 7146 3024 7164 3042
rect 7146 3042 7164 3060
rect 7146 3060 7164 3078
rect 7146 3078 7164 3096
rect 7146 3096 7164 3114
rect 7146 3114 7164 3132
rect 7146 3330 7164 3348
rect 7146 3348 7164 3366
rect 7146 3366 7164 3384
rect 7146 3384 7164 3402
rect 7146 3402 7164 3420
rect 7146 3420 7164 3438
rect 7146 3438 7164 3456
rect 7146 3456 7164 3474
rect 7146 3474 7164 3492
rect 7146 3492 7164 3510
rect 7146 3510 7164 3528
rect 7146 3528 7164 3546
rect 7146 3546 7164 3564
rect 7146 3564 7164 3582
rect 7146 3582 7164 3600
rect 7146 3600 7164 3618
rect 7146 3618 7164 3636
rect 7146 3636 7164 3654
rect 7146 3654 7164 3672
rect 7146 3672 7164 3690
rect 7146 3690 7164 3708
rect 7146 3708 7164 3726
rect 7146 3726 7164 3744
rect 7146 3744 7164 3762
rect 7146 3762 7164 3780
rect 7146 3780 7164 3798
rect 7146 3798 7164 3816
rect 7146 3816 7164 3834
rect 7146 3834 7164 3852
rect 7146 3852 7164 3870
rect 7146 3870 7164 3888
rect 7146 3888 7164 3906
rect 7146 3906 7164 3924
rect 7146 3924 7164 3942
rect 7146 3942 7164 3960
rect 7146 3960 7164 3978
rect 7146 3978 7164 3996
rect 7146 4212 7164 4230
rect 7146 4230 7164 4248
rect 7146 4248 7164 4266
rect 7146 4266 7164 4284
rect 7146 4284 7164 4302
rect 7146 4302 7164 4320
rect 7146 4320 7164 4338
rect 7146 4338 7164 4356
rect 7146 4356 7164 4374
rect 7146 4374 7164 4392
rect 7146 4392 7164 4410
rect 7146 4410 7164 4428
rect 7146 4428 7164 4446
rect 7146 4446 7164 4464
rect 7146 4464 7164 4482
rect 7146 4482 7164 4500
rect 7146 4500 7164 4518
rect 7146 4518 7164 4536
rect 7146 4536 7164 4554
rect 7146 4554 7164 4572
rect 7146 4572 7164 4590
rect 7146 4590 7164 4608
rect 7146 4608 7164 4626
rect 7146 4626 7164 4644
rect 7146 4644 7164 4662
rect 7146 4662 7164 4680
rect 7146 4680 7164 4698
rect 7146 4698 7164 4716
rect 7146 4716 7164 4734
rect 7146 4734 7164 4752
rect 7146 4752 7164 4770
rect 7146 4770 7164 4788
rect 7146 4788 7164 4806
rect 7146 4806 7164 4824
rect 7146 4824 7164 4842
rect 7146 4842 7164 4860
rect 7146 4860 7164 4878
rect 7146 4878 7164 4896
rect 7146 4896 7164 4914
rect 7146 4914 7164 4932
rect 7146 4932 7164 4950
rect 7146 4950 7164 4968
rect 7146 4968 7164 4986
rect 7146 4986 7164 5004
rect 7146 5004 7164 5022
rect 7146 5022 7164 5040
rect 7146 5040 7164 5058
rect 7146 5058 7164 5076
rect 7146 5076 7164 5094
rect 7146 5094 7164 5112
rect 7146 5112 7164 5130
rect 7146 5130 7164 5148
rect 7146 5148 7164 5166
rect 7146 5166 7164 5184
rect 7146 5184 7164 5202
rect 7146 5202 7164 5220
rect 7146 5220 7164 5238
rect 7146 5238 7164 5256
rect 7146 5256 7164 5274
rect 7146 5274 7164 5292
rect 7146 5292 7164 5310
rect 7146 5310 7164 5328
rect 7146 5328 7164 5346
rect 7146 5346 7164 5364
rect 7146 5364 7164 5382
rect 7146 5382 7164 5400
rect 7146 5400 7164 5418
rect 7146 5418 7164 5436
rect 7146 5436 7164 5454
rect 7146 5454 7164 5472
rect 7146 5472 7164 5490
rect 7146 5490 7164 5508
rect 7146 5508 7164 5526
rect 7146 5526 7164 5544
rect 7146 5544 7164 5562
rect 7146 5562 7164 5580
rect 7146 5580 7164 5598
rect 7146 5598 7164 5616
rect 7146 5616 7164 5634
rect 7146 5634 7164 5652
rect 7146 5652 7164 5670
rect 7146 5670 7164 5688
rect 7146 5688 7164 5706
rect 7146 5706 7164 5724
rect 7146 5724 7164 5742
rect 7146 5742 7164 5760
rect 7146 5760 7164 5778
rect 7146 5778 7164 5796
rect 7146 5796 7164 5814
rect 7146 5814 7164 5832
rect 7146 5832 7164 5850
rect 7146 5850 7164 5868
rect 7146 5868 7164 5886
rect 7146 5886 7164 5904
rect 7146 5904 7164 5922
rect 7146 5922 7164 5940
rect 7146 5940 7164 5958
rect 7146 5958 7164 5976
rect 7146 5976 7164 5994
rect 7146 5994 7164 6012
rect 7146 6012 7164 6030
rect 7146 6030 7164 6048
rect 7146 6048 7164 6066
rect 7146 6066 7164 6084
rect 7146 6084 7164 6102
rect 7146 6102 7164 6120
rect 7146 6120 7164 6138
rect 7146 6138 7164 6156
rect 7146 6156 7164 6174
rect 7146 6174 7164 6192
rect 7146 6192 7164 6210
rect 7146 6210 7164 6228
rect 7146 6228 7164 6246
rect 7146 6246 7164 6264
rect 7146 6264 7164 6282
rect 7146 6282 7164 6300
rect 7146 6300 7164 6318
rect 7146 6318 7164 6336
rect 7146 6336 7164 6354
rect 7146 6354 7164 6372
rect 7146 8298 7164 8316
rect 7146 8316 7164 8334
rect 7146 8334 7164 8352
rect 7146 8352 7164 8370
rect 7146 8370 7164 8388
rect 7146 8388 7164 8406
rect 7146 8406 7164 8424
rect 7146 8424 7164 8442
rect 7146 8442 7164 8460
rect 7146 8460 7164 8478
rect 7146 8478 7164 8496
rect 7146 8496 7164 8514
rect 7146 8514 7164 8532
rect 7146 8532 7164 8550
rect 7146 8550 7164 8568
rect 7146 8568 7164 8586
rect 7146 8586 7164 8604
rect 7146 8604 7164 8622
rect 7146 8622 7164 8640
rect 7146 8640 7164 8658
rect 7146 8658 7164 8676
rect 7146 8676 7164 8694
rect 7146 8694 7164 8712
rect 7146 8712 7164 8730
rect 7146 8730 7164 8748
rect 7146 8748 7164 8766
rect 7146 8766 7164 8784
rect 7146 8784 7164 8802
rect 7146 8802 7164 8820
rect 7146 8820 7164 8838
rect 7146 8838 7164 8856
rect 7146 8856 7164 8874
rect 7146 8874 7164 8892
rect 7146 8892 7164 8910
rect 7146 8910 7164 8928
rect 7146 8928 7164 8946
rect 7146 8946 7164 8964
rect 7146 8964 7164 8982
rect 7146 8982 7164 9000
rect 7146 9000 7164 9018
rect 7146 9018 7164 9036
rect 7146 9036 7164 9054
rect 7146 9054 7164 9072
rect 7146 9072 7164 9090
rect 7146 9090 7164 9108
rect 7146 9108 7164 9126
rect 7146 9126 7164 9144
rect 7146 9144 7164 9162
rect 7146 9162 7164 9180
rect 7146 9180 7164 9198
rect 7146 9198 7164 9216
rect 7146 9216 7164 9234
rect 7146 9234 7164 9252
rect 7146 9252 7164 9270
rect 7146 9270 7164 9288
rect 7146 9288 7164 9306
rect 7146 9306 7164 9324
rect 7146 9324 7164 9342
rect 7146 9342 7164 9360
rect 7146 9360 7164 9378
rect 7146 9378 7164 9396
rect 7146 9396 7164 9414
rect 7146 9414 7164 9432
rect 7146 9432 7164 9450
rect 7146 9450 7164 9468
rect 7146 9468 7164 9486
rect 7146 9486 7164 9504
rect 7146 9504 7164 9522
rect 7146 9522 7164 9540
rect 7146 9540 7164 9558
rect 7146 9558 7164 9576
rect 7146 9576 7164 9594
rect 7146 9594 7164 9612
rect 7146 9612 7164 9630
rect 7146 9630 7164 9648
rect 7146 9648 7164 9666
rect 7146 9666 7164 9684
rect 7146 9684 7164 9702
rect 7146 9702 7164 9720
rect 7146 9720 7164 9738
rect 7146 9738 7164 9756
rect 7146 9756 7164 9774
rect 7146 9774 7164 9792
rect 7146 9792 7164 9810
rect 7146 9810 7164 9828
rect 7146 9828 7164 9846
rect 7146 9846 7164 9864
rect 7146 9864 7164 9882
rect 7146 9882 7164 9900
rect 7146 9900 7164 9918
rect 7146 9918 7164 9936
rect 7146 9936 7164 9954
rect 7146 9954 7164 9972
rect 7146 9972 7164 9990
rect 7146 9990 7164 10008
rect 7146 10008 7164 10026
rect 7146 10026 7164 10044
rect 7146 10044 7164 10062
rect 7146 10062 7164 10080
rect 7146 10080 7164 10098
rect 7146 10098 7164 10116
rect 7146 10116 7164 10134
rect 7146 10134 7164 10152
rect 7146 10152 7164 10170
rect 7146 10170 7164 10188
rect 7146 10188 7164 10206
rect 7146 10206 7164 10224
rect 7146 10224 7164 10242
rect 7146 10242 7164 10260
rect 7146 10260 7164 10278
rect 7164 1890 7182 1908
rect 7164 1908 7182 1926
rect 7164 1926 7182 1944
rect 7164 1944 7182 1962
rect 7164 1962 7182 1980
rect 7164 1980 7182 1998
rect 7164 1998 7182 2016
rect 7164 2016 7182 2034
rect 7164 2034 7182 2052
rect 7164 2052 7182 2070
rect 7164 2070 7182 2088
rect 7164 2088 7182 2106
rect 7164 2106 7182 2124
rect 7164 2124 7182 2142
rect 7164 2142 7182 2160
rect 7164 2160 7182 2178
rect 7164 2178 7182 2196
rect 7164 2196 7182 2214
rect 7164 2214 7182 2232
rect 7164 2232 7182 2250
rect 7164 2250 7182 2268
rect 7164 2268 7182 2286
rect 7164 2286 7182 2304
rect 7164 2304 7182 2322
rect 7164 2322 7182 2340
rect 7164 2340 7182 2358
rect 7164 2358 7182 2376
rect 7164 2376 7182 2394
rect 7164 2394 7182 2412
rect 7164 2412 7182 2430
rect 7164 2430 7182 2448
rect 7164 2448 7182 2466
rect 7164 2466 7182 2484
rect 7164 2484 7182 2502
rect 7164 2502 7182 2520
rect 7164 2520 7182 2538
rect 7164 2538 7182 2556
rect 7164 2556 7182 2574
rect 7164 2574 7182 2592
rect 7164 2592 7182 2610
rect 7164 2610 7182 2628
rect 7164 2628 7182 2646
rect 7164 2646 7182 2664
rect 7164 2664 7182 2682
rect 7164 2682 7182 2700
rect 7164 2700 7182 2718
rect 7164 2718 7182 2736
rect 7164 2736 7182 2754
rect 7164 2754 7182 2772
rect 7164 2772 7182 2790
rect 7164 2790 7182 2808
rect 7164 2808 7182 2826
rect 7164 2826 7182 2844
rect 7164 2844 7182 2862
rect 7164 2862 7182 2880
rect 7164 2880 7182 2898
rect 7164 2898 7182 2916
rect 7164 2916 7182 2934
rect 7164 2934 7182 2952
rect 7164 2952 7182 2970
rect 7164 2970 7182 2988
rect 7164 2988 7182 3006
rect 7164 3006 7182 3024
rect 7164 3024 7182 3042
rect 7164 3042 7182 3060
rect 7164 3060 7182 3078
rect 7164 3078 7182 3096
rect 7164 3096 7182 3114
rect 7164 3114 7182 3132
rect 7164 3330 7182 3348
rect 7164 3348 7182 3366
rect 7164 3366 7182 3384
rect 7164 3384 7182 3402
rect 7164 3402 7182 3420
rect 7164 3420 7182 3438
rect 7164 3438 7182 3456
rect 7164 3456 7182 3474
rect 7164 3474 7182 3492
rect 7164 3492 7182 3510
rect 7164 3510 7182 3528
rect 7164 3528 7182 3546
rect 7164 3546 7182 3564
rect 7164 3564 7182 3582
rect 7164 3582 7182 3600
rect 7164 3600 7182 3618
rect 7164 3618 7182 3636
rect 7164 3636 7182 3654
rect 7164 3654 7182 3672
rect 7164 3672 7182 3690
rect 7164 3690 7182 3708
rect 7164 3708 7182 3726
rect 7164 3726 7182 3744
rect 7164 3744 7182 3762
rect 7164 3762 7182 3780
rect 7164 3780 7182 3798
rect 7164 3798 7182 3816
rect 7164 3816 7182 3834
rect 7164 3834 7182 3852
rect 7164 3852 7182 3870
rect 7164 3870 7182 3888
rect 7164 3888 7182 3906
rect 7164 3906 7182 3924
rect 7164 3924 7182 3942
rect 7164 3942 7182 3960
rect 7164 3960 7182 3978
rect 7164 3978 7182 3996
rect 7164 3996 7182 4014
rect 7164 4230 7182 4248
rect 7164 4248 7182 4266
rect 7164 4266 7182 4284
rect 7164 4284 7182 4302
rect 7164 4302 7182 4320
rect 7164 4320 7182 4338
rect 7164 4338 7182 4356
rect 7164 4356 7182 4374
rect 7164 4374 7182 4392
rect 7164 4392 7182 4410
rect 7164 4410 7182 4428
rect 7164 4428 7182 4446
rect 7164 4446 7182 4464
rect 7164 4464 7182 4482
rect 7164 4482 7182 4500
rect 7164 4500 7182 4518
rect 7164 4518 7182 4536
rect 7164 4536 7182 4554
rect 7164 4554 7182 4572
rect 7164 4572 7182 4590
rect 7164 4590 7182 4608
rect 7164 4608 7182 4626
rect 7164 4626 7182 4644
rect 7164 4644 7182 4662
rect 7164 4662 7182 4680
rect 7164 4680 7182 4698
rect 7164 4698 7182 4716
rect 7164 4716 7182 4734
rect 7164 4734 7182 4752
rect 7164 4752 7182 4770
rect 7164 4770 7182 4788
rect 7164 4788 7182 4806
rect 7164 4806 7182 4824
rect 7164 4824 7182 4842
rect 7164 4842 7182 4860
rect 7164 4860 7182 4878
rect 7164 4878 7182 4896
rect 7164 4896 7182 4914
rect 7164 4914 7182 4932
rect 7164 4932 7182 4950
rect 7164 4950 7182 4968
rect 7164 4968 7182 4986
rect 7164 4986 7182 5004
rect 7164 5004 7182 5022
rect 7164 5022 7182 5040
rect 7164 5040 7182 5058
rect 7164 5058 7182 5076
rect 7164 5076 7182 5094
rect 7164 5094 7182 5112
rect 7164 5112 7182 5130
rect 7164 5130 7182 5148
rect 7164 5148 7182 5166
rect 7164 5166 7182 5184
rect 7164 5184 7182 5202
rect 7164 5202 7182 5220
rect 7164 5220 7182 5238
rect 7164 5238 7182 5256
rect 7164 5256 7182 5274
rect 7164 5274 7182 5292
rect 7164 5292 7182 5310
rect 7164 5310 7182 5328
rect 7164 5328 7182 5346
rect 7164 5346 7182 5364
rect 7164 5364 7182 5382
rect 7164 5382 7182 5400
rect 7164 5400 7182 5418
rect 7164 5418 7182 5436
rect 7164 5436 7182 5454
rect 7164 5454 7182 5472
rect 7164 5472 7182 5490
rect 7164 5490 7182 5508
rect 7164 5508 7182 5526
rect 7164 5526 7182 5544
rect 7164 5544 7182 5562
rect 7164 5562 7182 5580
rect 7164 5580 7182 5598
rect 7164 5598 7182 5616
rect 7164 5616 7182 5634
rect 7164 5634 7182 5652
rect 7164 5652 7182 5670
rect 7164 5670 7182 5688
rect 7164 5688 7182 5706
rect 7164 5706 7182 5724
rect 7164 5724 7182 5742
rect 7164 5742 7182 5760
rect 7164 5760 7182 5778
rect 7164 5778 7182 5796
rect 7164 5796 7182 5814
rect 7164 5814 7182 5832
rect 7164 5832 7182 5850
rect 7164 5850 7182 5868
rect 7164 5868 7182 5886
rect 7164 5886 7182 5904
rect 7164 5904 7182 5922
rect 7164 5922 7182 5940
rect 7164 5940 7182 5958
rect 7164 5958 7182 5976
rect 7164 5976 7182 5994
rect 7164 5994 7182 6012
rect 7164 6012 7182 6030
rect 7164 6030 7182 6048
rect 7164 6048 7182 6066
rect 7164 6066 7182 6084
rect 7164 6084 7182 6102
rect 7164 6102 7182 6120
rect 7164 6120 7182 6138
rect 7164 6138 7182 6156
rect 7164 6156 7182 6174
rect 7164 6174 7182 6192
rect 7164 6192 7182 6210
rect 7164 6210 7182 6228
rect 7164 6228 7182 6246
rect 7164 6246 7182 6264
rect 7164 6264 7182 6282
rect 7164 6282 7182 6300
rect 7164 6300 7182 6318
rect 7164 6318 7182 6336
rect 7164 6336 7182 6354
rect 7164 6354 7182 6372
rect 7164 6372 7182 6390
rect 7164 8370 7182 8388
rect 7164 8388 7182 8406
rect 7164 8406 7182 8424
rect 7164 8424 7182 8442
rect 7164 8442 7182 8460
rect 7164 8460 7182 8478
rect 7164 8478 7182 8496
rect 7164 8496 7182 8514
rect 7164 8514 7182 8532
rect 7164 8532 7182 8550
rect 7164 8550 7182 8568
rect 7164 8568 7182 8586
rect 7164 8586 7182 8604
rect 7164 8604 7182 8622
rect 7164 8622 7182 8640
rect 7164 8640 7182 8658
rect 7164 8658 7182 8676
rect 7164 8676 7182 8694
rect 7164 8694 7182 8712
rect 7164 8712 7182 8730
rect 7164 8730 7182 8748
rect 7164 8748 7182 8766
rect 7164 8766 7182 8784
rect 7164 8784 7182 8802
rect 7164 8802 7182 8820
rect 7164 8820 7182 8838
rect 7164 8838 7182 8856
rect 7164 8856 7182 8874
rect 7164 8874 7182 8892
rect 7164 8892 7182 8910
rect 7164 8910 7182 8928
rect 7164 8928 7182 8946
rect 7164 8946 7182 8964
rect 7164 8964 7182 8982
rect 7164 8982 7182 9000
rect 7164 9000 7182 9018
rect 7164 9018 7182 9036
rect 7164 9036 7182 9054
rect 7164 9054 7182 9072
rect 7164 9072 7182 9090
rect 7164 9090 7182 9108
rect 7164 9108 7182 9126
rect 7164 9126 7182 9144
rect 7164 9144 7182 9162
rect 7164 9162 7182 9180
rect 7164 9180 7182 9198
rect 7164 9198 7182 9216
rect 7164 9216 7182 9234
rect 7164 9234 7182 9252
rect 7164 9252 7182 9270
rect 7164 9270 7182 9288
rect 7164 9288 7182 9306
rect 7164 9306 7182 9324
rect 7164 9324 7182 9342
rect 7164 9342 7182 9360
rect 7164 9360 7182 9378
rect 7164 9378 7182 9396
rect 7164 9396 7182 9414
rect 7164 9414 7182 9432
rect 7164 9432 7182 9450
rect 7164 9450 7182 9468
rect 7164 9468 7182 9486
rect 7164 9486 7182 9504
rect 7164 9504 7182 9522
rect 7164 9522 7182 9540
rect 7164 9540 7182 9558
rect 7164 9558 7182 9576
rect 7164 9576 7182 9594
rect 7164 9594 7182 9612
rect 7164 9612 7182 9630
rect 7164 9630 7182 9648
rect 7164 9648 7182 9666
rect 7164 9666 7182 9684
rect 7164 9684 7182 9702
rect 7164 9702 7182 9720
rect 7164 9720 7182 9738
rect 7164 9738 7182 9756
rect 7164 9756 7182 9774
rect 7164 9774 7182 9792
rect 7164 9792 7182 9810
rect 7164 9810 7182 9828
rect 7164 9828 7182 9846
rect 7164 9846 7182 9864
rect 7164 9864 7182 9882
rect 7164 9882 7182 9900
rect 7164 9900 7182 9918
rect 7164 9918 7182 9936
rect 7164 9936 7182 9954
rect 7164 9954 7182 9972
rect 7164 9972 7182 9990
rect 7164 9990 7182 10008
rect 7164 10008 7182 10026
rect 7164 10026 7182 10044
rect 7164 10044 7182 10062
rect 7164 10062 7182 10080
rect 7164 10080 7182 10098
rect 7164 10098 7182 10116
rect 7164 10116 7182 10134
rect 7164 10134 7182 10152
rect 7164 10152 7182 10170
rect 7164 10170 7182 10188
rect 7164 10188 7182 10206
rect 7182 1890 7200 1908
rect 7182 1908 7200 1926
rect 7182 1926 7200 1944
rect 7182 1944 7200 1962
rect 7182 1962 7200 1980
rect 7182 1980 7200 1998
rect 7182 1998 7200 2016
rect 7182 2016 7200 2034
rect 7182 2034 7200 2052
rect 7182 2052 7200 2070
rect 7182 2070 7200 2088
rect 7182 2088 7200 2106
rect 7182 2106 7200 2124
rect 7182 2124 7200 2142
rect 7182 2142 7200 2160
rect 7182 2160 7200 2178
rect 7182 2178 7200 2196
rect 7182 2196 7200 2214
rect 7182 2214 7200 2232
rect 7182 2232 7200 2250
rect 7182 2250 7200 2268
rect 7182 2268 7200 2286
rect 7182 2286 7200 2304
rect 7182 2304 7200 2322
rect 7182 2322 7200 2340
rect 7182 2340 7200 2358
rect 7182 2358 7200 2376
rect 7182 2376 7200 2394
rect 7182 2394 7200 2412
rect 7182 2412 7200 2430
rect 7182 2430 7200 2448
rect 7182 2448 7200 2466
rect 7182 2466 7200 2484
rect 7182 2484 7200 2502
rect 7182 2502 7200 2520
rect 7182 2520 7200 2538
rect 7182 2538 7200 2556
rect 7182 2556 7200 2574
rect 7182 2574 7200 2592
rect 7182 2592 7200 2610
rect 7182 2610 7200 2628
rect 7182 2628 7200 2646
rect 7182 2646 7200 2664
rect 7182 2664 7200 2682
rect 7182 2682 7200 2700
rect 7182 2700 7200 2718
rect 7182 2718 7200 2736
rect 7182 2736 7200 2754
rect 7182 2754 7200 2772
rect 7182 2772 7200 2790
rect 7182 2790 7200 2808
rect 7182 2808 7200 2826
rect 7182 2826 7200 2844
rect 7182 2844 7200 2862
rect 7182 2862 7200 2880
rect 7182 2880 7200 2898
rect 7182 2898 7200 2916
rect 7182 2916 7200 2934
rect 7182 2934 7200 2952
rect 7182 2952 7200 2970
rect 7182 2970 7200 2988
rect 7182 2988 7200 3006
rect 7182 3006 7200 3024
rect 7182 3024 7200 3042
rect 7182 3042 7200 3060
rect 7182 3060 7200 3078
rect 7182 3078 7200 3096
rect 7182 3096 7200 3114
rect 7182 3114 7200 3132
rect 7182 3132 7200 3150
rect 7182 3348 7200 3366
rect 7182 3366 7200 3384
rect 7182 3384 7200 3402
rect 7182 3402 7200 3420
rect 7182 3420 7200 3438
rect 7182 3438 7200 3456
rect 7182 3456 7200 3474
rect 7182 3474 7200 3492
rect 7182 3492 7200 3510
rect 7182 3510 7200 3528
rect 7182 3528 7200 3546
rect 7182 3546 7200 3564
rect 7182 3564 7200 3582
rect 7182 3582 7200 3600
rect 7182 3600 7200 3618
rect 7182 3618 7200 3636
rect 7182 3636 7200 3654
rect 7182 3654 7200 3672
rect 7182 3672 7200 3690
rect 7182 3690 7200 3708
rect 7182 3708 7200 3726
rect 7182 3726 7200 3744
rect 7182 3744 7200 3762
rect 7182 3762 7200 3780
rect 7182 3780 7200 3798
rect 7182 3798 7200 3816
rect 7182 3816 7200 3834
rect 7182 3834 7200 3852
rect 7182 3852 7200 3870
rect 7182 3870 7200 3888
rect 7182 3888 7200 3906
rect 7182 3906 7200 3924
rect 7182 3924 7200 3942
rect 7182 3942 7200 3960
rect 7182 3960 7200 3978
rect 7182 3978 7200 3996
rect 7182 3996 7200 4014
rect 7182 4014 7200 4032
rect 7182 4248 7200 4266
rect 7182 4266 7200 4284
rect 7182 4284 7200 4302
rect 7182 4302 7200 4320
rect 7182 4320 7200 4338
rect 7182 4338 7200 4356
rect 7182 4356 7200 4374
rect 7182 4374 7200 4392
rect 7182 4392 7200 4410
rect 7182 4410 7200 4428
rect 7182 4428 7200 4446
rect 7182 4446 7200 4464
rect 7182 4464 7200 4482
rect 7182 4482 7200 4500
rect 7182 4500 7200 4518
rect 7182 4518 7200 4536
rect 7182 4536 7200 4554
rect 7182 4554 7200 4572
rect 7182 4572 7200 4590
rect 7182 4590 7200 4608
rect 7182 4608 7200 4626
rect 7182 4626 7200 4644
rect 7182 4644 7200 4662
rect 7182 4662 7200 4680
rect 7182 4680 7200 4698
rect 7182 4698 7200 4716
rect 7182 4716 7200 4734
rect 7182 4734 7200 4752
rect 7182 4752 7200 4770
rect 7182 4770 7200 4788
rect 7182 4788 7200 4806
rect 7182 4806 7200 4824
rect 7182 4824 7200 4842
rect 7182 4842 7200 4860
rect 7182 4860 7200 4878
rect 7182 4878 7200 4896
rect 7182 4896 7200 4914
rect 7182 4914 7200 4932
rect 7182 4932 7200 4950
rect 7182 4950 7200 4968
rect 7182 4968 7200 4986
rect 7182 4986 7200 5004
rect 7182 5004 7200 5022
rect 7182 5022 7200 5040
rect 7182 5040 7200 5058
rect 7182 5058 7200 5076
rect 7182 5076 7200 5094
rect 7182 5094 7200 5112
rect 7182 5112 7200 5130
rect 7182 5130 7200 5148
rect 7182 5148 7200 5166
rect 7182 5166 7200 5184
rect 7182 5184 7200 5202
rect 7182 5202 7200 5220
rect 7182 5220 7200 5238
rect 7182 5238 7200 5256
rect 7182 5256 7200 5274
rect 7182 5274 7200 5292
rect 7182 5292 7200 5310
rect 7182 5310 7200 5328
rect 7182 5328 7200 5346
rect 7182 5346 7200 5364
rect 7182 5364 7200 5382
rect 7182 5382 7200 5400
rect 7182 5400 7200 5418
rect 7182 5418 7200 5436
rect 7182 5436 7200 5454
rect 7182 5454 7200 5472
rect 7182 5472 7200 5490
rect 7182 5490 7200 5508
rect 7182 5508 7200 5526
rect 7182 5526 7200 5544
rect 7182 5544 7200 5562
rect 7182 5562 7200 5580
rect 7182 5580 7200 5598
rect 7182 5598 7200 5616
rect 7182 5616 7200 5634
rect 7182 5634 7200 5652
rect 7182 5652 7200 5670
rect 7182 5670 7200 5688
rect 7182 5688 7200 5706
rect 7182 5706 7200 5724
rect 7182 5724 7200 5742
rect 7182 5742 7200 5760
rect 7182 5760 7200 5778
rect 7182 5778 7200 5796
rect 7182 5796 7200 5814
rect 7182 5814 7200 5832
rect 7182 5832 7200 5850
rect 7182 5850 7200 5868
rect 7182 5868 7200 5886
rect 7182 5886 7200 5904
rect 7182 5904 7200 5922
rect 7182 5922 7200 5940
rect 7182 5940 7200 5958
rect 7182 5958 7200 5976
rect 7182 5976 7200 5994
rect 7182 5994 7200 6012
rect 7182 6012 7200 6030
rect 7182 6030 7200 6048
rect 7182 6048 7200 6066
rect 7182 6066 7200 6084
rect 7182 6084 7200 6102
rect 7182 6102 7200 6120
rect 7182 6120 7200 6138
rect 7182 6138 7200 6156
rect 7182 6156 7200 6174
rect 7182 6174 7200 6192
rect 7182 6192 7200 6210
rect 7182 6210 7200 6228
rect 7182 6228 7200 6246
rect 7182 6246 7200 6264
rect 7182 6264 7200 6282
rect 7182 6282 7200 6300
rect 7182 6300 7200 6318
rect 7182 6318 7200 6336
rect 7182 6336 7200 6354
rect 7182 6354 7200 6372
rect 7182 6372 7200 6390
rect 7182 6390 7200 6408
rect 7182 8424 7200 8442
rect 7182 8442 7200 8460
rect 7182 8460 7200 8478
rect 7182 8478 7200 8496
rect 7182 8496 7200 8514
rect 7182 8514 7200 8532
rect 7182 8532 7200 8550
rect 7182 8550 7200 8568
rect 7182 8568 7200 8586
rect 7182 8586 7200 8604
rect 7182 8604 7200 8622
rect 7182 8622 7200 8640
rect 7182 8640 7200 8658
rect 7182 8658 7200 8676
rect 7182 8676 7200 8694
rect 7182 8694 7200 8712
rect 7182 8712 7200 8730
rect 7182 8730 7200 8748
rect 7182 8748 7200 8766
rect 7182 8766 7200 8784
rect 7182 8784 7200 8802
rect 7182 8802 7200 8820
rect 7182 8820 7200 8838
rect 7182 8838 7200 8856
rect 7182 8856 7200 8874
rect 7182 8874 7200 8892
rect 7182 8892 7200 8910
rect 7182 8910 7200 8928
rect 7182 8928 7200 8946
rect 7182 8946 7200 8964
rect 7182 8964 7200 8982
rect 7182 8982 7200 9000
rect 7182 9000 7200 9018
rect 7182 9018 7200 9036
rect 7182 9036 7200 9054
rect 7182 9054 7200 9072
rect 7182 9072 7200 9090
rect 7182 9090 7200 9108
rect 7182 9108 7200 9126
rect 7182 9126 7200 9144
rect 7182 9144 7200 9162
rect 7182 9162 7200 9180
rect 7182 9180 7200 9198
rect 7182 9198 7200 9216
rect 7182 9216 7200 9234
rect 7182 9234 7200 9252
rect 7182 9252 7200 9270
rect 7182 9270 7200 9288
rect 7182 9288 7200 9306
rect 7182 9306 7200 9324
rect 7182 9324 7200 9342
rect 7182 9342 7200 9360
rect 7182 9360 7200 9378
rect 7182 9378 7200 9396
rect 7182 9396 7200 9414
rect 7182 9414 7200 9432
rect 7182 9432 7200 9450
rect 7182 9450 7200 9468
rect 7182 9468 7200 9486
rect 7182 9486 7200 9504
rect 7182 9504 7200 9522
rect 7182 9522 7200 9540
rect 7182 9540 7200 9558
rect 7182 9558 7200 9576
rect 7182 9576 7200 9594
rect 7182 9594 7200 9612
rect 7182 9612 7200 9630
rect 7182 9630 7200 9648
rect 7182 9648 7200 9666
rect 7182 9666 7200 9684
rect 7182 9684 7200 9702
rect 7182 9702 7200 9720
rect 7182 9720 7200 9738
rect 7182 9738 7200 9756
rect 7182 9756 7200 9774
rect 7182 9774 7200 9792
rect 7182 9792 7200 9810
rect 7182 9810 7200 9828
rect 7182 9828 7200 9846
rect 7182 9846 7200 9864
rect 7182 9864 7200 9882
rect 7182 9882 7200 9900
rect 7182 9900 7200 9918
rect 7182 9918 7200 9936
rect 7182 9936 7200 9954
rect 7182 9954 7200 9972
rect 7182 9972 7200 9990
rect 7182 9990 7200 10008
rect 7182 10008 7200 10026
rect 7182 10026 7200 10044
rect 7182 10044 7200 10062
rect 7182 10062 7200 10080
rect 7182 10080 7200 10098
rect 7182 10098 7200 10116
rect 7182 10116 7200 10134
rect 7200 1908 7218 1926
rect 7200 1926 7218 1944
rect 7200 1944 7218 1962
rect 7200 1962 7218 1980
rect 7200 1980 7218 1998
rect 7200 1998 7218 2016
rect 7200 2016 7218 2034
rect 7200 2034 7218 2052
rect 7200 2052 7218 2070
rect 7200 2070 7218 2088
rect 7200 2088 7218 2106
rect 7200 2106 7218 2124
rect 7200 2124 7218 2142
rect 7200 2142 7218 2160
rect 7200 2160 7218 2178
rect 7200 2178 7218 2196
rect 7200 2196 7218 2214
rect 7200 2214 7218 2232
rect 7200 2232 7218 2250
rect 7200 2250 7218 2268
rect 7200 2268 7218 2286
rect 7200 2286 7218 2304
rect 7200 2304 7218 2322
rect 7200 2322 7218 2340
rect 7200 2340 7218 2358
rect 7200 2358 7218 2376
rect 7200 2376 7218 2394
rect 7200 2394 7218 2412
rect 7200 2412 7218 2430
rect 7200 2430 7218 2448
rect 7200 2448 7218 2466
rect 7200 2466 7218 2484
rect 7200 2484 7218 2502
rect 7200 2502 7218 2520
rect 7200 2520 7218 2538
rect 7200 2538 7218 2556
rect 7200 2556 7218 2574
rect 7200 2574 7218 2592
rect 7200 2592 7218 2610
rect 7200 2610 7218 2628
rect 7200 2628 7218 2646
rect 7200 2646 7218 2664
rect 7200 2664 7218 2682
rect 7200 2682 7218 2700
rect 7200 2700 7218 2718
rect 7200 2718 7218 2736
rect 7200 2736 7218 2754
rect 7200 2754 7218 2772
rect 7200 2772 7218 2790
rect 7200 2790 7218 2808
rect 7200 2808 7218 2826
rect 7200 2826 7218 2844
rect 7200 2844 7218 2862
rect 7200 2862 7218 2880
rect 7200 2880 7218 2898
rect 7200 2898 7218 2916
rect 7200 2916 7218 2934
rect 7200 2934 7218 2952
rect 7200 2952 7218 2970
rect 7200 2970 7218 2988
rect 7200 2988 7218 3006
rect 7200 3006 7218 3024
rect 7200 3024 7218 3042
rect 7200 3042 7218 3060
rect 7200 3060 7218 3078
rect 7200 3078 7218 3096
rect 7200 3096 7218 3114
rect 7200 3114 7218 3132
rect 7200 3132 7218 3150
rect 7200 3348 7218 3366
rect 7200 3366 7218 3384
rect 7200 3384 7218 3402
rect 7200 3402 7218 3420
rect 7200 3420 7218 3438
rect 7200 3438 7218 3456
rect 7200 3456 7218 3474
rect 7200 3474 7218 3492
rect 7200 3492 7218 3510
rect 7200 3510 7218 3528
rect 7200 3528 7218 3546
rect 7200 3546 7218 3564
rect 7200 3564 7218 3582
rect 7200 3582 7218 3600
rect 7200 3600 7218 3618
rect 7200 3618 7218 3636
rect 7200 3636 7218 3654
rect 7200 3654 7218 3672
rect 7200 3672 7218 3690
rect 7200 3690 7218 3708
rect 7200 3708 7218 3726
rect 7200 3726 7218 3744
rect 7200 3744 7218 3762
rect 7200 3762 7218 3780
rect 7200 3780 7218 3798
rect 7200 3798 7218 3816
rect 7200 3816 7218 3834
rect 7200 3834 7218 3852
rect 7200 3852 7218 3870
rect 7200 3870 7218 3888
rect 7200 3888 7218 3906
rect 7200 3906 7218 3924
rect 7200 3924 7218 3942
rect 7200 3942 7218 3960
rect 7200 3960 7218 3978
rect 7200 3978 7218 3996
rect 7200 3996 7218 4014
rect 7200 4014 7218 4032
rect 7200 4032 7218 4050
rect 7200 4266 7218 4284
rect 7200 4284 7218 4302
rect 7200 4302 7218 4320
rect 7200 4320 7218 4338
rect 7200 4338 7218 4356
rect 7200 4356 7218 4374
rect 7200 4374 7218 4392
rect 7200 4392 7218 4410
rect 7200 4410 7218 4428
rect 7200 4428 7218 4446
rect 7200 4446 7218 4464
rect 7200 4464 7218 4482
rect 7200 4482 7218 4500
rect 7200 4500 7218 4518
rect 7200 4518 7218 4536
rect 7200 4536 7218 4554
rect 7200 4554 7218 4572
rect 7200 4572 7218 4590
rect 7200 4590 7218 4608
rect 7200 4608 7218 4626
rect 7200 4626 7218 4644
rect 7200 4644 7218 4662
rect 7200 4662 7218 4680
rect 7200 4680 7218 4698
rect 7200 4698 7218 4716
rect 7200 4716 7218 4734
rect 7200 4734 7218 4752
rect 7200 4752 7218 4770
rect 7200 4770 7218 4788
rect 7200 4788 7218 4806
rect 7200 4806 7218 4824
rect 7200 4824 7218 4842
rect 7200 4842 7218 4860
rect 7200 4860 7218 4878
rect 7200 4878 7218 4896
rect 7200 4896 7218 4914
rect 7200 4914 7218 4932
rect 7200 4932 7218 4950
rect 7200 4950 7218 4968
rect 7200 4968 7218 4986
rect 7200 4986 7218 5004
rect 7200 5004 7218 5022
rect 7200 5022 7218 5040
rect 7200 5040 7218 5058
rect 7200 5058 7218 5076
rect 7200 5076 7218 5094
rect 7200 5094 7218 5112
rect 7200 5112 7218 5130
rect 7200 5130 7218 5148
rect 7200 5148 7218 5166
rect 7200 5166 7218 5184
rect 7200 5184 7218 5202
rect 7200 5202 7218 5220
rect 7200 5220 7218 5238
rect 7200 5238 7218 5256
rect 7200 5256 7218 5274
rect 7200 5274 7218 5292
rect 7200 5292 7218 5310
rect 7200 5310 7218 5328
rect 7200 5328 7218 5346
rect 7200 5346 7218 5364
rect 7200 5364 7218 5382
rect 7200 5382 7218 5400
rect 7200 5400 7218 5418
rect 7200 5418 7218 5436
rect 7200 5436 7218 5454
rect 7200 5454 7218 5472
rect 7200 5472 7218 5490
rect 7200 5490 7218 5508
rect 7200 5508 7218 5526
rect 7200 5526 7218 5544
rect 7200 5544 7218 5562
rect 7200 5562 7218 5580
rect 7200 5580 7218 5598
rect 7200 5598 7218 5616
rect 7200 5616 7218 5634
rect 7200 5634 7218 5652
rect 7200 5652 7218 5670
rect 7200 5670 7218 5688
rect 7200 5688 7218 5706
rect 7200 5706 7218 5724
rect 7200 5724 7218 5742
rect 7200 5742 7218 5760
rect 7200 5760 7218 5778
rect 7200 5778 7218 5796
rect 7200 5796 7218 5814
rect 7200 5814 7218 5832
rect 7200 5832 7218 5850
rect 7200 5850 7218 5868
rect 7200 5868 7218 5886
rect 7200 5886 7218 5904
rect 7200 5904 7218 5922
rect 7200 5922 7218 5940
rect 7200 5940 7218 5958
rect 7200 5958 7218 5976
rect 7200 5976 7218 5994
rect 7200 5994 7218 6012
rect 7200 6012 7218 6030
rect 7200 6030 7218 6048
rect 7200 6048 7218 6066
rect 7200 6066 7218 6084
rect 7200 6084 7218 6102
rect 7200 6102 7218 6120
rect 7200 6120 7218 6138
rect 7200 6138 7218 6156
rect 7200 6156 7218 6174
rect 7200 6174 7218 6192
rect 7200 6192 7218 6210
rect 7200 6210 7218 6228
rect 7200 6228 7218 6246
rect 7200 6246 7218 6264
rect 7200 6264 7218 6282
rect 7200 6282 7218 6300
rect 7200 6300 7218 6318
rect 7200 6318 7218 6336
rect 7200 6336 7218 6354
rect 7200 6354 7218 6372
rect 7200 6372 7218 6390
rect 7200 6390 7218 6408
rect 7200 6408 7218 6426
rect 7200 8478 7218 8496
rect 7200 8496 7218 8514
rect 7200 8514 7218 8532
rect 7200 8532 7218 8550
rect 7200 8550 7218 8568
rect 7200 8568 7218 8586
rect 7200 8586 7218 8604
rect 7200 8604 7218 8622
rect 7200 8622 7218 8640
rect 7200 8640 7218 8658
rect 7200 8658 7218 8676
rect 7200 8676 7218 8694
rect 7200 8694 7218 8712
rect 7200 8712 7218 8730
rect 7200 8730 7218 8748
rect 7200 8748 7218 8766
rect 7200 8766 7218 8784
rect 7200 8784 7218 8802
rect 7200 8802 7218 8820
rect 7200 8820 7218 8838
rect 7200 8838 7218 8856
rect 7200 8856 7218 8874
rect 7200 8874 7218 8892
rect 7200 8892 7218 8910
rect 7200 8910 7218 8928
rect 7200 8928 7218 8946
rect 7200 8946 7218 8964
rect 7200 8964 7218 8982
rect 7200 8982 7218 9000
rect 7200 9000 7218 9018
rect 7200 9018 7218 9036
rect 7200 9036 7218 9054
rect 7200 9054 7218 9072
rect 7200 9072 7218 9090
rect 7200 9090 7218 9108
rect 7200 9108 7218 9126
rect 7200 9126 7218 9144
rect 7200 9144 7218 9162
rect 7200 9162 7218 9180
rect 7200 9180 7218 9198
rect 7200 9198 7218 9216
rect 7200 9216 7218 9234
rect 7200 9234 7218 9252
rect 7200 9252 7218 9270
rect 7200 9270 7218 9288
rect 7200 9288 7218 9306
rect 7200 9306 7218 9324
rect 7200 9324 7218 9342
rect 7200 9342 7218 9360
rect 7200 9360 7218 9378
rect 7200 9378 7218 9396
rect 7200 9396 7218 9414
rect 7200 9414 7218 9432
rect 7200 9432 7218 9450
rect 7200 9450 7218 9468
rect 7200 9468 7218 9486
rect 7200 9486 7218 9504
rect 7200 9504 7218 9522
rect 7200 9522 7218 9540
rect 7200 9540 7218 9558
rect 7200 9558 7218 9576
rect 7200 9576 7218 9594
rect 7200 9594 7218 9612
rect 7200 9612 7218 9630
rect 7200 9630 7218 9648
rect 7200 9648 7218 9666
rect 7200 9666 7218 9684
rect 7200 9684 7218 9702
rect 7200 9702 7218 9720
rect 7200 9720 7218 9738
rect 7200 9738 7218 9756
rect 7200 9756 7218 9774
rect 7200 9774 7218 9792
rect 7200 9792 7218 9810
rect 7200 9810 7218 9828
rect 7200 9828 7218 9846
rect 7200 9846 7218 9864
rect 7200 9864 7218 9882
rect 7200 9882 7218 9900
rect 7200 9900 7218 9918
rect 7200 9918 7218 9936
rect 7200 9936 7218 9954
rect 7200 9954 7218 9972
rect 7200 9972 7218 9990
rect 7200 9990 7218 10008
rect 7200 10008 7218 10026
rect 7200 10026 7218 10044
rect 7200 10044 7218 10062
rect 7218 1926 7236 1944
rect 7218 1944 7236 1962
rect 7218 1962 7236 1980
rect 7218 1980 7236 1998
rect 7218 1998 7236 2016
rect 7218 2016 7236 2034
rect 7218 2034 7236 2052
rect 7218 2052 7236 2070
rect 7218 2070 7236 2088
rect 7218 2088 7236 2106
rect 7218 2106 7236 2124
rect 7218 2124 7236 2142
rect 7218 2142 7236 2160
rect 7218 2160 7236 2178
rect 7218 2178 7236 2196
rect 7218 2196 7236 2214
rect 7218 2214 7236 2232
rect 7218 2232 7236 2250
rect 7218 2250 7236 2268
rect 7218 2268 7236 2286
rect 7218 2286 7236 2304
rect 7218 2304 7236 2322
rect 7218 2322 7236 2340
rect 7218 2340 7236 2358
rect 7218 2358 7236 2376
rect 7218 2376 7236 2394
rect 7218 2394 7236 2412
rect 7218 2412 7236 2430
rect 7218 2430 7236 2448
rect 7218 2448 7236 2466
rect 7218 2466 7236 2484
rect 7218 2484 7236 2502
rect 7218 2502 7236 2520
rect 7218 2520 7236 2538
rect 7218 2538 7236 2556
rect 7218 2556 7236 2574
rect 7218 2574 7236 2592
rect 7218 2592 7236 2610
rect 7218 2610 7236 2628
rect 7218 2628 7236 2646
rect 7218 2646 7236 2664
rect 7218 2664 7236 2682
rect 7218 2682 7236 2700
rect 7218 2700 7236 2718
rect 7218 2718 7236 2736
rect 7218 2736 7236 2754
rect 7218 2754 7236 2772
rect 7218 2772 7236 2790
rect 7218 2790 7236 2808
rect 7218 2808 7236 2826
rect 7218 2826 7236 2844
rect 7218 2844 7236 2862
rect 7218 2862 7236 2880
rect 7218 2880 7236 2898
rect 7218 2898 7236 2916
rect 7218 2916 7236 2934
rect 7218 2934 7236 2952
rect 7218 2952 7236 2970
rect 7218 2970 7236 2988
rect 7218 2988 7236 3006
rect 7218 3006 7236 3024
rect 7218 3024 7236 3042
rect 7218 3042 7236 3060
rect 7218 3060 7236 3078
rect 7218 3078 7236 3096
rect 7218 3096 7236 3114
rect 7218 3114 7236 3132
rect 7218 3132 7236 3150
rect 7218 3348 7236 3366
rect 7218 3366 7236 3384
rect 7218 3384 7236 3402
rect 7218 3402 7236 3420
rect 7218 3420 7236 3438
rect 7218 3438 7236 3456
rect 7218 3456 7236 3474
rect 7218 3474 7236 3492
rect 7218 3492 7236 3510
rect 7218 3510 7236 3528
rect 7218 3528 7236 3546
rect 7218 3546 7236 3564
rect 7218 3564 7236 3582
rect 7218 3582 7236 3600
rect 7218 3600 7236 3618
rect 7218 3618 7236 3636
rect 7218 3636 7236 3654
rect 7218 3654 7236 3672
rect 7218 3672 7236 3690
rect 7218 3690 7236 3708
rect 7218 3708 7236 3726
rect 7218 3726 7236 3744
rect 7218 3744 7236 3762
rect 7218 3762 7236 3780
rect 7218 3780 7236 3798
rect 7218 3798 7236 3816
rect 7218 3816 7236 3834
rect 7218 3834 7236 3852
rect 7218 3852 7236 3870
rect 7218 3870 7236 3888
rect 7218 3888 7236 3906
rect 7218 3906 7236 3924
rect 7218 3924 7236 3942
rect 7218 3942 7236 3960
rect 7218 3960 7236 3978
rect 7218 3978 7236 3996
rect 7218 3996 7236 4014
rect 7218 4014 7236 4032
rect 7218 4032 7236 4050
rect 7218 4050 7236 4068
rect 7218 4302 7236 4320
rect 7218 4320 7236 4338
rect 7218 4338 7236 4356
rect 7218 4356 7236 4374
rect 7218 4374 7236 4392
rect 7218 4392 7236 4410
rect 7218 4410 7236 4428
rect 7218 4428 7236 4446
rect 7218 4446 7236 4464
rect 7218 4464 7236 4482
rect 7218 4482 7236 4500
rect 7218 4500 7236 4518
rect 7218 4518 7236 4536
rect 7218 4536 7236 4554
rect 7218 4554 7236 4572
rect 7218 4572 7236 4590
rect 7218 4590 7236 4608
rect 7218 4608 7236 4626
rect 7218 4626 7236 4644
rect 7218 4644 7236 4662
rect 7218 4662 7236 4680
rect 7218 4680 7236 4698
rect 7218 4698 7236 4716
rect 7218 4716 7236 4734
rect 7218 4734 7236 4752
rect 7218 4752 7236 4770
rect 7218 4770 7236 4788
rect 7218 4788 7236 4806
rect 7218 4806 7236 4824
rect 7218 4824 7236 4842
rect 7218 4842 7236 4860
rect 7218 4860 7236 4878
rect 7218 4878 7236 4896
rect 7218 4896 7236 4914
rect 7218 4914 7236 4932
rect 7218 4932 7236 4950
rect 7218 4950 7236 4968
rect 7218 4968 7236 4986
rect 7218 4986 7236 5004
rect 7218 5004 7236 5022
rect 7218 5022 7236 5040
rect 7218 5040 7236 5058
rect 7218 5058 7236 5076
rect 7218 5076 7236 5094
rect 7218 5094 7236 5112
rect 7218 5112 7236 5130
rect 7218 5130 7236 5148
rect 7218 5148 7236 5166
rect 7218 5166 7236 5184
rect 7218 5184 7236 5202
rect 7218 5202 7236 5220
rect 7218 5220 7236 5238
rect 7218 5238 7236 5256
rect 7218 5256 7236 5274
rect 7218 5274 7236 5292
rect 7218 5292 7236 5310
rect 7218 5310 7236 5328
rect 7218 5328 7236 5346
rect 7218 5346 7236 5364
rect 7218 5364 7236 5382
rect 7218 5382 7236 5400
rect 7218 5400 7236 5418
rect 7218 5418 7236 5436
rect 7218 5436 7236 5454
rect 7218 5454 7236 5472
rect 7218 5472 7236 5490
rect 7218 5490 7236 5508
rect 7218 5508 7236 5526
rect 7218 5526 7236 5544
rect 7218 5544 7236 5562
rect 7218 5562 7236 5580
rect 7218 5580 7236 5598
rect 7218 5598 7236 5616
rect 7218 5616 7236 5634
rect 7218 5634 7236 5652
rect 7218 5652 7236 5670
rect 7218 5670 7236 5688
rect 7218 5688 7236 5706
rect 7218 5706 7236 5724
rect 7218 5724 7236 5742
rect 7218 5742 7236 5760
rect 7218 5760 7236 5778
rect 7218 5778 7236 5796
rect 7218 5796 7236 5814
rect 7218 5814 7236 5832
rect 7218 5832 7236 5850
rect 7218 5850 7236 5868
rect 7218 5868 7236 5886
rect 7218 5886 7236 5904
rect 7218 5904 7236 5922
rect 7218 5922 7236 5940
rect 7218 5940 7236 5958
rect 7218 5958 7236 5976
rect 7218 5976 7236 5994
rect 7218 5994 7236 6012
rect 7218 6012 7236 6030
rect 7218 6030 7236 6048
rect 7218 6048 7236 6066
rect 7218 6066 7236 6084
rect 7218 6084 7236 6102
rect 7218 6102 7236 6120
rect 7218 6120 7236 6138
rect 7218 6138 7236 6156
rect 7218 6156 7236 6174
rect 7218 6174 7236 6192
rect 7218 6192 7236 6210
rect 7218 6210 7236 6228
rect 7218 6228 7236 6246
rect 7218 6246 7236 6264
rect 7218 6264 7236 6282
rect 7218 6282 7236 6300
rect 7218 6300 7236 6318
rect 7218 6318 7236 6336
rect 7218 6336 7236 6354
rect 7218 6354 7236 6372
rect 7218 6372 7236 6390
rect 7218 6390 7236 6408
rect 7218 6408 7236 6426
rect 7218 6426 7236 6444
rect 7218 8550 7236 8568
rect 7218 8568 7236 8586
rect 7218 8586 7236 8604
rect 7218 8604 7236 8622
rect 7218 8622 7236 8640
rect 7218 8640 7236 8658
rect 7218 8658 7236 8676
rect 7218 8676 7236 8694
rect 7218 8694 7236 8712
rect 7218 8712 7236 8730
rect 7218 8730 7236 8748
rect 7218 8748 7236 8766
rect 7218 8766 7236 8784
rect 7218 8784 7236 8802
rect 7218 8802 7236 8820
rect 7218 8820 7236 8838
rect 7218 8838 7236 8856
rect 7218 8856 7236 8874
rect 7218 8874 7236 8892
rect 7218 8892 7236 8910
rect 7218 8910 7236 8928
rect 7218 8928 7236 8946
rect 7218 8946 7236 8964
rect 7218 8964 7236 8982
rect 7218 8982 7236 9000
rect 7218 9000 7236 9018
rect 7218 9018 7236 9036
rect 7218 9036 7236 9054
rect 7218 9054 7236 9072
rect 7218 9072 7236 9090
rect 7218 9090 7236 9108
rect 7218 9108 7236 9126
rect 7218 9126 7236 9144
rect 7218 9144 7236 9162
rect 7218 9162 7236 9180
rect 7218 9180 7236 9198
rect 7218 9198 7236 9216
rect 7218 9216 7236 9234
rect 7218 9234 7236 9252
rect 7218 9252 7236 9270
rect 7218 9270 7236 9288
rect 7218 9288 7236 9306
rect 7218 9306 7236 9324
rect 7218 9324 7236 9342
rect 7218 9342 7236 9360
rect 7218 9360 7236 9378
rect 7218 9378 7236 9396
rect 7218 9396 7236 9414
rect 7218 9414 7236 9432
rect 7218 9432 7236 9450
rect 7218 9450 7236 9468
rect 7218 9468 7236 9486
rect 7218 9486 7236 9504
rect 7218 9504 7236 9522
rect 7218 9522 7236 9540
rect 7218 9540 7236 9558
rect 7218 9558 7236 9576
rect 7218 9576 7236 9594
rect 7218 9594 7236 9612
rect 7218 9612 7236 9630
rect 7218 9630 7236 9648
rect 7218 9648 7236 9666
rect 7218 9666 7236 9684
rect 7218 9684 7236 9702
rect 7218 9702 7236 9720
rect 7218 9720 7236 9738
rect 7218 9738 7236 9756
rect 7218 9756 7236 9774
rect 7218 9774 7236 9792
rect 7218 9792 7236 9810
rect 7218 9810 7236 9828
rect 7218 9828 7236 9846
rect 7218 9846 7236 9864
rect 7218 9864 7236 9882
rect 7218 9882 7236 9900
rect 7218 9900 7236 9918
rect 7218 9918 7236 9936
rect 7218 9936 7236 9954
rect 7218 9954 7236 9972
rect 7218 9972 7236 9990
rect 7236 1926 7254 1944
rect 7236 1944 7254 1962
rect 7236 1962 7254 1980
rect 7236 1980 7254 1998
rect 7236 1998 7254 2016
rect 7236 2016 7254 2034
rect 7236 2034 7254 2052
rect 7236 2052 7254 2070
rect 7236 2070 7254 2088
rect 7236 2088 7254 2106
rect 7236 2106 7254 2124
rect 7236 2124 7254 2142
rect 7236 2142 7254 2160
rect 7236 2160 7254 2178
rect 7236 2178 7254 2196
rect 7236 2196 7254 2214
rect 7236 2214 7254 2232
rect 7236 2232 7254 2250
rect 7236 2250 7254 2268
rect 7236 2268 7254 2286
rect 7236 2286 7254 2304
rect 7236 2304 7254 2322
rect 7236 2322 7254 2340
rect 7236 2340 7254 2358
rect 7236 2358 7254 2376
rect 7236 2376 7254 2394
rect 7236 2394 7254 2412
rect 7236 2412 7254 2430
rect 7236 2430 7254 2448
rect 7236 2448 7254 2466
rect 7236 2466 7254 2484
rect 7236 2484 7254 2502
rect 7236 2502 7254 2520
rect 7236 2520 7254 2538
rect 7236 2538 7254 2556
rect 7236 2556 7254 2574
rect 7236 2574 7254 2592
rect 7236 2592 7254 2610
rect 7236 2610 7254 2628
rect 7236 2628 7254 2646
rect 7236 2646 7254 2664
rect 7236 2664 7254 2682
rect 7236 2682 7254 2700
rect 7236 2700 7254 2718
rect 7236 2718 7254 2736
rect 7236 2736 7254 2754
rect 7236 2754 7254 2772
rect 7236 2772 7254 2790
rect 7236 2790 7254 2808
rect 7236 2808 7254 2826
rect 7236 2826 7254 2844
rect 7236 2844 7254 2862
rect 7236 2862 7254 2880
rect 7236 2880 7254 2898
rect 7236 2898 7254 2916
rect 7236 2916 7254 2934
rect 7236 2934 7254 2952
rect 7236 2952 7254 2970
rect 7236 2970 7254 2988
rect 7236 2988 7254 3006
rect 7236 3006 7254 3024
rect 7236 3024 7254 3042
rect 7236 3042 7254 3060
rect 7236 3060 7254 3078
rect 7236 3078 7254 3096
rect 7236 3096 7254 3114
rect 7236 3114 7254 3132
rect 7236 3132 7254 3150
rect 7236 3150 7254 3168
rect 7236 3366 7254 3384
rect 7236 3384 7254 3402
rect 7236 3402 7254 3420
rect 7236 3420 7254 3438
rect 7236 3438 7254 3456
rect 7236 3456 7254 3474
rect 7236 3474 7254 3492
rect 7236 3492 7254 3510
rect 7236 3510 7254 3528
rect 7236 3528 7254 3546
rect 7236 3546 7254 3564
rect 7236 3564 7254 3582
rect 7236 3582 7254 3600
rect 7236 3600 7254 3618
rect 7236 3618 7254 3636
rect 7236 3636 7254 3654
rect 7236 3654 7254 3672
rect 7236 3672 7254 3690
rect 7236 3690 7254 3708
rect 7236 3708 7254 3726
rect 7236 3726 7254 3744
rect 7236 3744 7254 3762
rect 7236 3762 7254 3780
rect 7236 3780 7254 3798
rect 7236 3798 7254 3816
rect 7236 3816 7254 3834
rect 7236 3834 7254 3852
rect 7236 3852 7254 3870
rect 7236 3870 7254 3888
rect 7236 3888 7254 3906
rect 7236 3906 7254 3924
rect 7236 3924 7254 3942
rect 7236 3942 7254 3960
rect 7236 3960 7254 3978
rect 7236 3978 7254 3996
rect 7236 3996 7254 4014
rect 7236 4014 7254 4032
rect 7236 4032 7254 4050
rect 7236 4050 7254 4068
rect 7236 4068 7254 4086
rect 7236 4320 7254 4338
rect 7236 4338 7254 4356
rect 7236 4356 7254 4374
rect 7236 4374 7254 4392
rect 7236 4392 7254 4410
rect 7236 4410 7254 4428
rect 7236 4428 7254 4446
rect 7236 4446 7254 4464
rect 7236 4464 7254 4482
rect 7236 4482 7254 4500
rect 7236 4500 7254 4518
rect 7236 4518 7254 4536
rect 7236 4536 7254 4554
rect 7236 4554 7254 4572
rect 7236 4572 7254 4590
rect 7236 4590 7254 4608
rect 7236 4608 7254 4626
rect 7236 4626 7254 4644
rect 7236 4644 7254 4662
rect 7236 4662 7254 4680
rect 7236 4680 7254 4698
rect 7236 4698 7254 4716
rect 7236 4716 7254 4734
rect 7236 4734 7254 4752
rect 7236 4752 7254 4770
rect 7236 4770 7254 4788
rect 7236 4788 7254 4806
rect 7236 4806 7254 4824
rect 7236 4824 7254 4842
rect 7236 4842 7254 4860
rect 7236 4860 7254 4878
rect 7236 4878 7254 4896
rect 7236 4896 7254 4914
rect 7236 4914 7254 4932
rect 7236 4932 7254 4950
rect 7236 4950 7254 4968
rect 7236 4968 7254 4986
rect 7236 4986 7254 5004
rect 7236 5004 7254 5022
rect 7236 5022 7254 5040
rect 7236 5040 7254 5058
rect 7236 5058 7254 5076
rect 7236 5076 7254 5094
rect 7236 5094 7254 5112
rect 7236 5112 7254 5130
rect 7236 5130 7254 5148
rect 7236 5148 7254 5166
rect 7236 5166 7254 5184
rect 7236 5184 7254 5202
rect 7236 5202 7254 5220
rect 7236 5220 7254 5238
rect 7236 5238 7254 5256
rect 7236 5256 7254 5274
rect 7236 5274 7254 5292
rect 7236 5292 7254 5310
rect 7236 5310 7254 5328
rect 7236 5328 7254 5346
rect 7236 5346 7254 5364
rect 7236 5364 7254 5382
rect 7236 5382 7254 5400
rect 7236 5400 7254 5418
rect 7236 5418 7254 5436
rect 7236 5436 7254 5454
rect 7236 5454 7254 5472
rect 7236 5472 7254 5490
rect 7236 5490 7254 5508
rect 7236 5508 7254 5526
rect 7236 5526 7254 5544
rect 7236 5544 7254 5562
rect 7236 5562 7254 5580
rect 7236 5580 7254 5598
rect 7236 5598 7254 5616
rect 7236 5616 7254 5634
rect 7236 5634 7254 5652
rect 7236 5652 7254 5670
rect 7236 5670 7254 5688
rect 7236 5688 7254 5706
rect 7236 5706 7254 5724
rect 7236 5724 7254 5742
rect 7236 5742 7254 5760
rect 7236 5760 7254 5778
rect 7236 5778 7254 5796
rect 7236 5796 7254 5814
rect 7236 5814 7254 5832
rect 7236 5832 7254 5850
rect 7236 5850 7254 5868
rect 7236 5868 7254 5886
rect 7236 5886 7254 5904
rect 7236 5904 7254 5922
rect 7236 5922 7254 5940
rect 7236 5940 7254 5958
rect 7236 5958 7254 5976
rect 7236 5976 7254 5994
rect 7236 5994 7254 6012
rect 7236 6012 7254 6030
rect 7236 6030 7254 6048
rect 7236 6048 7254 6066
rect 7236 6066 7254 6084
rect 7236 6084 7254 6102
rect 7236 6102 7254 6120
rect 7236 6120 7254 6138
rect 7236 6138 7254 6156
rect 7236 6156 7254 6174
rect 7236 6174 7254 6192
rect 7236 6192 7254 6210
rect 7236 6210 7254 6228
rect 7236 6228 7254 6246
rect 7236 6246 7254 6264
rect 7236 6264 7254 6282
rect 7236 6282 7254 6300
rect 7236 6300 7254 6318
rect 7236 6318 7254 6336
rect 7236 6336 7254 6354
rect 7236 6354 7254 6372
rect 7236 6372 7254 6390
rect 7236 6390 7254 6408
rect 7236 6408 7254 6426
rect 7236 6426 7254 6444
rect 7236 6444 7254 6462
rect 7236 8622 7254 8640
rect 7236 8640 7254 8658
rect 7236 8658 7254 8676
rect 7236 8676 7254 8694
rect 7236 8694 7254 8712
rect 7236 8712 7254 8730
rect 7236 8730 7254 8748
rect 7236 8748 7254 8766
rect 7236 8766 7254 8784
rect 7236 8784 7254 8802
rect 7236 8802 7254 8820
rect 7236 8820 7254 8838
rect 7236 8838 7254 8856
rect 7236 8856 7254 8874
rect 7236 8874 7254 8892
rect 7236 8892 7254 8910
rect 7236 8910 7254 8928
rect 7236 8928 7254 8946
rect 7236 8946 7254 8964
rect 7236 8964 7254 8982
rect 7236 8982 7254 9000
rect 7236 9000 7254 9018
rect 7236 9018 7254 9036
rect 7236 9036 7254 9054
rect 7236 9054 7254 9072
rect 7236 9072 7254 9090
rect 7236 9090 7254 9108
rect 7236 9108 7254 9126
rect 7236 9126 7254 9144
rect 7236 9144 7254 9162
rect 7236 9162 7254 9180
rect 7236 9180 7254 9198
rect 7236 9198 7254 9216
rect 7236 9216 7254 9234
rect 7236 9234 7254 9252
rect 7236 9252 7254 9270
rect 7236 9270 7254 9288
rect 7236 9288 7254 9306
rect 7236 9306 7254 9324
rect 7236 9324 7254 9342
rect 7236 9342 7254 9360
rect 7236 9360 7254 9378
rect 7236 9378 7254 9396
rect 7236 9396 7254 9414
rect 7236 9414 7254 9432
rect 7236 9432 7254 9450
rect 7236 9450 7254 9468
rect 7236 9468 7254 9486
rect 7236 9486 7254 9504
rect 7236 9504 7254 9522
rect 7236 9522 7254 9540
rect 7236 9540 7254 9558
rect 7236 9558 7254 9576
rect 7236 9576 7254 9594
rect 7236 9594 7254 9612
rect 7236 9612 7254 9630
rect 7236 9630 7254 9648
rect 7236 9648 7254 9666
rect 7236 9666 7254 9684
rect 7236 9684 7254 9702
rect 7236 9702 7254 9720
rect 7236 9720 7254 9738
rect 7236 9738 7254 9756
rect 7236 9756 7254 9774
rect 7236 9774 7254 9792
rect 7236 9792 7254 9810
rect 7236 9810 7254 9828
rect 7236 9828 7254 9846
rect 7236 9846 7254 9864
rect 7236 9864 7254 9882
rect 7236 9882 7254 9900
rect 7236 9900 7254 9918
rect 7254 1944 7272 1962
rect 7254 1962 7272 1980
rect 7254 1980 7272 1998
rect 7254 1998 7272 2016
rect 7254 2016 7272 2034
rect 7254 2034 7272 2052
rect 7254 2052 7272 2070
rect 7254 2070 7272 2088
rect 7254 2088 7272 2106
rect 7254 2106 7272 2124
rect 7254 2124 7272 2142
rect 7254 2142 7272 2160
rect 7254 2160 7272 2178
rect 7254 2178 7272 2196
rect 7254 2196 7272 2214
rect 7254 2214 7272 2232
rect 7254 2232 7272 2250
rect 7254 2250 7272 2268
rect 7254 2268 7272 2286
rect 7254 2286 7272 2304
rect 7254 2304 7272 2322
rect 7254 2322 7272 2340
rect 7254 2340 7272 2358
rect 7254 2358 7272 2376
rect 7254 2376 7272 2394
rect 7254 2394 7272 2412
rect 7254 2412 7272 2430
rect 7254 2430 7272 2448
rect 7254 2448 7272 2466
rect 7254 2466 7272 2484
rect 7254 2484 7272 2502
rect 7254 2502 7272 2520
rect 7254 2520 7272 2538
rect 7254 2538 7272 2556
rect 7254 2556 7272 2574
rect 7254 2574 7272 2592
rect 7254 2592 7272 2610
rect 7254 2610 7272 2628
rect 7254 2628 7272 2646
rect 7254 2646 7272 2664
rect 7254 2664 7272 2682
rect 7254 2682 7272 2700
rect 7254 2700 7272 2718
rect 7254 2718 7272 2736
rect 7254 2736 7272 2754
rect 7254 2754 7272 2772
rect 7254 2772 7272 2790
rect 7254 2790 7272 2808
rect 7254 2808 7272 2826
rect 7254 2826 7272 2844
rect 7254 2844 7272 2862
rect 7254 2862 7272 2880
rect 7254 2880 7272 2898
rect 7254 2898 7272 2916
rect 7254 2916 7272 2934
rect 7254 2934 7272 2952
rect 7254 2952 7272 2970
rect 7254 2970 7272 2988
rect 7254 2988 7272 3006
rect 7254 3006 7272 3024
rect 7254 3024 7272 3042
rect 7254 3042 7272 3060
rect 7254 3060 7272 3078
rect 7254 3078 7272 3096
rect 7254 3096 7272 3114
rect 7254 3114 7272 3132
rect 7254 3132 7272 3150
rect 7254 3150 7272 3168
rect 7254 3366 7272 3384
rect 7254 3384 7272 3402
rect 7254 3402 7272 3420
rect 7254 3420 7272 3438
rect 7254 3438 7272 3456
rect 7254 3456 7272 3474
rect 7254 3474 7272 3492
rect 7254 3492 7272 3510
rect 7254 3510 7272 3528
rect 7254 3528 7272 3546
rect 7254 3546 7272 3564
rect 7254 3564 7272 3582
rect 7254 3582 7272 3600
rect 7254 3600 7272 3618
rect 7254 3618 7272 3636
rect 7254 3636 7272 3654
rect 7254 3654 7272 3672
rect 7254 3672 7272 3690
rect 7254 3690 7272 3708
rect 7254 3708 7272 3726
rect 7254 3726 7272 3744
rect 7254 3744 7272 3762
rect 7254 3762 7272 3780
rect 7254 3780 7272 3798
rect 7254 3798 7272 3816
rect 7254 3816 7272 3834
rect 7254 3834 7272 3852
rect 7254 3852 7272 3870
rect 7254 3870 7272 3888
rect 7254 3888 7272 3906
rect 7254 3906 7272 3924
rect 7254 3924 7272 3942
rect 7254 3942 7272 3960
rect 7254 3960 7272 3978
rect 7254 3978 7272 3996
rect 7254 3996 7272 4014
rect 7254 4014 7272 4032
rect 7254 4032 7272 4050
rect 7254 4338 7272 4356
rect 7254 4356 7272 4374
rect 7254 4374 7272 4392
rect 7254 4392 7272 4410
rect 7254 4410 7272 4428
rect 7254 4428 7272 4446
rect 7254 4446 7272 4464
rect 7254 4464 7272 4482
rect 7254 4482 7272 4500
rect 7254 4500 7272 4518
rect 7254 4518 7272 4536
rect 7254 4536 7272 4554
rect 7254 4554 7272 4572
rect 7254 4572 7272 4590
rect 7254 4590 7272 4608
rect 7254 4608 7272 4626
rect 7254 4626 7272 4644
rect 7254 4644 7272 4662
rect 7254 4662 7272 4680
rect 7254 4680 7272 4698
rect 7254 4698 7272 4716
rect 7254 4716 7272 4734
rect 7254 4734 7272 4752
rect 7254 4752 7272 4770
rect 7254 4770 7272 4788
rect 7254 4788 7272 4806
rect 7254 4806 7272 4824
rect 7254 4824 7272 4842
rect 7254 4842 7272 4860
rect 7254 4860 7272 4878
rect 7254 4878 7272 4896
rect 7254 4896 7272 4914
rect 7254 4914 7272 4932
rect 7254 4932 7272 4950
rect 7254 4950 7272 4968
rect 7254 4968 7272 4986
rect 7254 4986 7272 5004
rect 7254 5004 7272 5022
rect 7254 5022 7272 5040
rect 7254 5040 7272 5058
rect 7254 5058 7272 5076
rect 7254 5076 7272 5094
rect 7254 5094 7272 5112
rect 7254 5112 7272 5130
rect 7254 5130 7272 5148
rect 7254 5148 7272 5166
rect 7254 5166 7272 5184
rect 7254 5184 7272 5202
rect 7254 5202 7272 5220
rect 7254 5220 7272 5238
rect 7254 5238 7272 5256
rect 7254 5256 7272 5274
rect 7254 5274 7272 5292
rect 7254 5292 7272 5310
rect 7254 5310 7272 5328
rect 7254 5328 7272 5346
rect 7254 5346 7272 5364
rect 7254 5364 7272 5382
rect 7254 5382 7272 5400
rect 7254 5400 7272 5418
rect 7254 5418 7272 5436
rect 7254 5436 7272 5454
rect 7254 5454 7272 5472
rect 7254 5472 7272 5490
rect 7254 5490 7272 5508
rect 7254 5508 7272 5526
rect 7254 5526 7272 5544
rect 7254 5544 7272 5562
rect 7254 5562 7272 5580
rect 7254 5580 7272 5598
rect 7254 5598 7272 5616
rect 7254 5616 7272 5634
rect 7254 5634 7272 5652
rect 7254 5652 7272 5670
rect 7254 5670 7272 5688
rect 7254 5688 7272 5706
rect 7254 5706 7272 5724
rect 7254 5724 7272 5742
rect 7254 5742 7272 5760
rect 7254 5760 7272 5778
rect 7254 5778 7272 5796
rect 7254 5796 7272 5814
rect 7254 5814 7272 5832
rect 7254 5832 7272 5850
rect 7254 5850 7272 5868
rect 7254 5868 7272 5886
rect 7254 5886 7272 5904
rect 7254 5904 7272 5922
rect 7254 5922 7272 5940
rect 7254 5940 7272 5958
rect 7254 5958 7272 5976
rect 7254 5976 7272 5994
rect 7254 5994 7272 6012
rect 7254 6012 7272 6030
rect 7254 6030 7272 6048
rect 7254 6048 7272 6066
rect 7254 6066 7272 6084
rect 7254 6084 7272 6102
rect 7254 6102 7272 6120
rect 7254 6120 7272 6138
rect 7254 6138 7272 6156
rect 7254 6156 7272 6174
rect 7254 6174 7272 6192
rect 7254 6192 7272 6210
rect 7254 6210 7272 6228
rect 7254 6228 7272 6246
rect 7254 6246 7272 6264
rect 7254 6264 7272 6282
rect 7254 6282 7272 6300
rect 7254 6300 7272 6318
rect 7254 6318 7272 6336
rect 7254 6336 7272 6354
rect 7254 6354 7272 6372
rect 7254 6372 7272 6390
rect 7254 6390 7272 6408
rect 7254 6408 7272 6426
rect 7254 6426 7272 6444
rect 7254 6444 7272 6462
rect 7254 8694 7272 8712
rect 7254 8712 7272 8730
rect 7254 8730 7272 8748
rect 7254 8748 7272 8766
rect 7254 8766 7272 8784
rect 7254 8784 7272 8802
rect 7254 8802 7272 8820
rect 7254 8820 7272 8838
rect 7254 8838 7272 8856
rect 7254 8856 7272 8874
rect 7254 8874 7272 8892
rect 7254 8892 7272 8910
rect 7254 8910 7272 8928
rect 7254 8928 7272 8946
rect 7254 8946 7272 8964
rect 7254 8964 7272 8982
rect 7254 8982 7272 9000
rect 7254 9000 7272 9018
rect 7254 9018 7272 9036
rect 7254 9036 7272 9054
rect 7254 9054 7272 9072
rect 7254 9072 7272 9090
rect 7254 9090 7272 9108
rect 7254 9108 7272 9126
rect 7254 9126 7272 9144
rect 7254 9144 7272 9162
rect 7254 9162 7272 9180
rect 7254 9180 7272 9198
rect 7254 9198 7272 9216
rect 7254 9216 7272 9234
rect 7254 9234 7272 9252
rect 7254 9252 7272 9270
rect 7254 9270 7272 9288
rect 7254 9288 7272 9306
rect 7254 9306 7272 9324
rect 7254 9324 7272 9342
rect 7254 9342 7272 9360
rect 7254 9360 7272 9378
rect 7254 9378 7272 9396
rect 7254 9396 7272 9414
rect 7254 9414 7272 9432
rect 7254 9432 7272 9450
rect 7254 9450 7272 9468
rect 7254 9468 7272 9486
rect 7254 9486 7272 9504
rect 7254 9504 7272 9522
rect 7254 9522 7272 9540
rect 7254 9540 7272 9558
rect 7254 9558 7272 9576
rect 7254 9576 7272 9594
rect 7254 9594 7272 9612
rect 7254 9612 7272 9630
rect 7254 9630 7272 9648
rect 7254 9648 7272 9666
rect 7254 9666 7272 9684
rect 7254 9684 7272 9702
rect 7254 9702 7272 9720
rect 7254 9720 7272 9738
rect 7254 9738 7272 9756
rect 7254 9756 7272 9774
rect 7254 9774 7272 9792
rect 7254 9792 7272 9810
rect 7254 9810 7272 9828
rect 7272 1944 7290 1962
rect 7272 1962 7290 1980
rect 7272 1980 7290 1998
rect 7272 1998 7290 2016
rect 7272 2016 7290 2034
rect 7272 2034 7290 2052
rect 7272 2052 7290 2070
rect 7272 2070 7290 2088
rect 7272 2088 7290 2106
rect 7272 2106 7290 2124
rect 7272 2124 7290 2142
rect 7272 2142 7290 2160
rect 7272 2160 7290 2178
rect 7272 2178 7290 2196
rect 7272 2196 7290 2214
rect 7272 2214 7290 2232
rect 7272 2232 7290 2250
rect 7272 2250 7290 2268
rect 7272 2268 7290 2286
rect 7272 2286 7290 2304
rect 7272 2304 7290 2322
rect 7272 2322 7290 2340
rect 7272 2340 7290 2358
rect 7272 2358 7290 2376
rect 7272 2376 7290 2394
rect 7272 2394 7290 2412
rect 7272 2412 7290 2430
rect 7272 2430 7290 2448
rect 7272 2448 7290 2466
rect 7272 2466 7290 2484
rect 7272 2484 7290 2502
rect 7272 2502 7290 2520
rect 7272 2520 7290 2538
rect 7272 2538 7290 2556
rect 7272 2556 7290 2574
rect 7272 2574 7290 2592
rect 7272 2592 7290 2610
rect 7272 2610 7290 2628
rect 7272 2628 7290 2646
rect 7272 2646 7290 2664
rect 7272 2664 7290 2682
rect 7272 2682 7290 2700
rect 7272 2700 7290 2718
rect 7272 2718 7290 2736
rect 7272 2736 7290 2754
rect 7272 2754 7290 2772
rect 7272 2772 7290 2790
rect 7272 2790 7290 2808
rect 7272 2808 7290 2826
rect 7272 2826 7290 2844
rect 7272 2844 7290 2862
rect 7272 2862 7290 2880
rect 7272 2880 7290 2898
rect 7272 2898 7290 2916
rect 7272 2916 7290 2934
rect 7272 2934 7290 2952
rect 7272 2952 7290 2970
rect 7272 2970 7290 2988
rect 7272 2988 7290 3006
rect 7272 3006 7290 3024
rect 7272 3024 7290 3042
rect 7272 3042 7290 3060
rect 7272 3060 7290 3078
rect 7272 3078 7290 3096
rect 7272 3096 7290 3114
rect 7272 3114 7290 3132
rect 7272 3132 7290 3150
rect 7272 3150 7290 3168
rect 7272 3438 7290 3456
rect 7272 3456 7290 3474
rect 7272 3474 7290 3492
rect 7272 3492 7290 3510
rect 7272 3510 7290 3528
rect 7272 3528 7290 3546
rect 7272 3546 7290 3564
rect 7272 3564 7290 3582
rect 7272 3582 7290 3600
rect 7272 3600 7290 3618
rect 7272 3618 7290 3636
rect 7272 3636 7290 3654
rect 7272 3654 7290 3672
rect 7272 3672 7290 3690
rect 7272 3690 7290 3708
rect 7272 3708 7290 3726
rect 7272 3726 7290 3744
rect 7272 3744 7290 3762
rect 7272 3762 7290 3780
rect 7272 3780 7290 3798
rect 7272 3798 7290 3816
rect 7272 3816 7290 3834
rect 7272 3834 7290 3852
rect 7272 3852 7290 3870
rect 7272 3870 7290 3888
rect 7272 3888 7290 3906
rect 7272 3906 7290 3924
rect 7272 3924 7290 3942
rect 7272 4356 7290 4374
rect 7272 4374 7290 4392
rect 7272 4392 7290 4410
rect 7272 4410 7290 4428
rect 7272 4428 7290 4446
rect 7272 4446 7290 4464
rect 7272 4464 7290 4482
rect 7272 4482 7290 4500
rect 7272 4500 7290 4518
rect 7272 4518 7290 4536
rect 7272 4536 7290 4554
rect 7272 4554 7290 4572
rect 7272 4572 7290 4590
rect 7272 4590 7290 4608
rect 7272 4608 7290 4626
rect 7272 4626 7290 4644
rect 7272 4644 7290 4662
rect 7272 4662 7290 4680
rect 7272 4680 7290 4698
rect 7272 4698 7290 4716
rect 7272 4716 7290 4734
rect 7272 4734 7290 4752
rect 7272 4752 7290 4770
rect 7272 4770 7290 4788
rect 7272 4788 7290 4806
rect 7272 4806 7290 4824
rect 7272 4824 7290 4842
rect 7272 4842 7290 4860
rect 7272 4860 7290 4878
rect 7272 4878 7290 4896
rect 7272 4896 7290 4914
rect 7272 4914 7290 4932
rect 7272 4932 7290 4950
rect 7272 4950 7290 4968
rect 7272 4968 7290 4986
rect 7272 4986 7290 5004
rect 7272 5004 7290 5022
rect 7272 5022 7290 5040
rect 7272 5040 7290 5058
rect 7272 5058 7290 5076
rect 7272 5076 7290 5094
rect 7272 5094 7290 5112
rect 7272 5112 7290 5130
rect 7272 5130 7290 5148
rect 7272 5148 7290 5166
rect 7272 5166 7290 5184
rect 7272 5184 7290 5202
rect 7272 5202 7290 5220
rect 7272 5220 7290 5238
rect 7272 5238 7290 5256
rect 7272 5256 7290 5274
rect 7272 5274 7290 5292
rect 7272 5292 7290 5310
rect 7272 5310 7290 5328
rect 7272 5328 7290 5346
rect 7272 5346 7290 5364
rect 7272 5364 7290 5382
rect 7272 5382 7290 5400
rect 7272 5400 7290 5418
rect 7272 5418 7290 5436
rect 7272 5436 7290 5454
rect 7272 5454 7290 5472
rect 7272 5472 7290 5490
rect 7272 5490 7290 5508
rect 7272 5508 7290 5526
rect 7272 5526 7290 5544
rect 7272 5544 7290 5562
rect 7272 5562 7290 5580
rect 7272 5580 7290 5598
rect 7272 5598 7290 5616
rect 7272 5616 7290 5634
rect 7272 5634 7290 5652
rect 7272 5652 7290 5670
rect 7272 5670 7290 5688
rect 7272 5688 7290 5706
rect 7272 5706 7290 5724
rect 7272 5724 7290 5742
rect 7272 5742 7290 5760
rect 7272 5760 7290 5778
rect 7272 5778 7290 5796
rect 7272 5796 7290 5814
rect 7272 5814 7290 5832
rect 7272 5832 7290 5850
rect 7272 5850 7290 5868
rect 7272 5868 7290 5886
rect 7272 5886 7290 5904
rect 7272 5904 7290 5922
rect 7272 5922 7290 5940
rect 7272 5940 7290 5958
rect 7272 5958 7290 5976
rect 7272 5976 7290 5994
rect 7272 5994 7290 6012
rect 7272 6012 7290 6030
rect 7272 6030 7290 6048
rect 7272 6048 7290 6066
rect 7272 6066 7290 6084
rect 7272 6084 7290 6102
rect 7272 6102 7290 6120
rect 7272 6120 7290 6138
rect 7272 6138 7290 6156
rect 7272 6156 7290 6174
rect 7272 6174 7290 6192
rect 7272 6192 7290 6210
rect 7272 6210 7290 6228
rect 7272 6228 7290 6246
rect 7272 6246 7290 6264
rect 7272 6264 7290 6282
rect 7272 6282 7290 6300
rect 7272 6300 7290 6318
rect 7272 6318 7290 6336
rect 7272 6336 7290 6354
rect 7272 6354 7290 6372
rect 7272 6372 7290 6390
rect 7272 6390 7290 6408
rect 7272 6408 7290 6426
rect 7272 6426 7290 6444
rect 7272 6444 7290 6462
rect 7272 6462 7290 6480
rect 7272 8766 7290 8784
rect 7272 8784 7290 8802
rect 7272 8802 7290 8820
rect 7272 8820 7290 8838
rect 7272 8838 7290 8856
rect 7272 8856 7290 8874
rect 7272 8874 7290 8892
rect 7272 8892 7290 8910
rect 7272 8910 7290 8928
rect 7272 8928 7290 8946
rect 7272 8946 7290 8964
rect 7272 8964 7290 8982
rect 7272 8982 7290 9000
rect 7272 9000 7290 9018
rect 7272 9018 7290 9036
rect 7272 9036 7290 9054
rect 7272 9054 7290 9072
rect 7272 9072 7290 9090
rect 7272 9090 7290 9108
rect 7272 9108 7290 9126
rect 7272 9126 7290 9144
rect 7272 9144 7290 9162
rect 7272 9162 7290 9180
rect 7272 9180 7290 9198
rect 7272 9198 7290 9216
rect 7272 9216 7290 9234
rect 7272 9234 7290 9252
rect 7272 9252 7290 9270
rect 7272 9270 7290 9288
rect 7272 9288 7290 9306
rect 7272 9306 7290 9324
rect 7272 9324 7290 9342
rect 7272 9342 7290 9360
rect 7272 9360 7290 9378
rect 7272 9378 7290 9396
rect 7272 9396 7290 9414
rect 7272 9414 7290 9432
rect 7272 9432 7290 9450
rect 7272 9450 7290 9468
rect 7272 9468 7290 9486
rect 7272 9486 7290 9504
rect 7272 9504 7290 9522
rect 7272 9522 7290 9540
rect 7272 9540 7290 9558
rect 7272 9558 7290 9576
rect 7272 9576 7290 9594
rect 7272 9594 7290 9612
rect 7272 9612 7290 9630
rect 7272 9630 7290 9648
rect 7272 9648 7290 9666
rect 7272 9666 7290 9684
rect 7272 9684 7290 9702
rect 7272 9702 7290 9720
rect 7272 9720 7290 9738
rect 7290 1962 7308 1980
rect 7290 1980 7308 1998
rect 7290 1998 7308 2016
rect 7290 2016 7308 2034
rect 7290 2034 7308 2052
rect 7290 2052 7308 2070
rect 7290 2070 7308 2088
rect 7290 2088 7308 2106
rect 7290 2106 7308 2124
rect 7290 2124 7308 2142
rect 7290 2142 7308 2160
rect 7290 2160 7308 2178
rect 7290 2178 7308 2196
rect 7290 2196 7308 2214
rect 7290 2214 7308 2232
rect 7290 2232 7308 2250
rect 7290 2250 7308 2268
rect 7290 2268 7308 2286
rect 7290 2286 7308 2304
rect 7290 2304 7308 2322
rect 7290 2322 7308 2340
rect 7290 2340 7308 2358
rect 7290 2358 7308 2376
rect 7290 2376 7308 2394
rect 7290 2394 7308 2412
rect 7290 2412 7308 2430
rect 7290 2430 7308 2448
rect 7290 2448 7308 2466
rect 7290 2466 7308 2484
rect 7290 2484 7308 2502
rect 7290 2502 7308 2520
rect 7290 2520 7308 2538
rect 7290 2538 7308 2556
rect 7290 2556 7308 2574
rect 7290 2574 7308 2592
rect 7290 2592 7308 2610
rect 7290 2610 7308 2628
rect 7290 2628 7308 2646
rect 7290 2646 7308 2664
rect 7290 2664 7308 2682
rect 7290 2682 7308 2700
rect 7290 2700 7308 2718
rect 7290 2718 7308 2736
rect 7290 2736 7308 2754
rect 7290 2754 7308 2772
rect 7290 2772 7308 2790
rect 7290 2790 7308 2808
rect 7290 2808 7308 2826
rect 7290 2826 7308 2844
rect 7290 2844 7308 2862
rect 7290 2862 7308 2880
rect 7290 2880 7308 2898
rect 7290 2898 7308 2916
rect 7290 2916 7308 2934
rect 7290 2934 7308 2952
rect 7290 2952 7308 2970
rect 7290 2970 7308 2988
rect 7290 2988 7308 3006
rect 7290 3006 7308 3024
rect 7290 3024 7308 3042
rect 7290 3042 7308 3060
rect 7290 3060 7308 3078
rect 7290 3078 7308 3096
rect 7290 3096 7308 3114
rect 7290 3114 7308 3132
rect 7290 3132 7308 3150
rect 7290 3150 7308 3168
rect 7290 4392 7308 4410
rect 7290 4410 7308 4428
rect 7290 4428 7308 4446
rect 7290 4446 7308 4464
rect 7290 4464 7308 4482
rect 7290 4482 7308 4500
rect 7290 4500 7308 4518
rect 7290 4518 7308 4536
rect 7290 4536 7308 4554
rect 7290 4554 7308 4572
rect 7290 4572 7308 4590
rect 7290 4590 7308 4608
rect 7290 4608 7308 4626
rect 7290 4626 7308 4644
rect 7290 4644 7308 4662
rect 7290 4662 7308 4680
rect 7290 4680 7308 4698
rect 7290 4698 7308 4716
rect 7290 4716 7308 4734
rect 7290 4734 7308 4752
rect 7290 4752 7308 4770
rect 7290 4770 7308 4788
rect 7290 4788 7308 4806
rect 7290 4806 7308 4824
rect 7290 4824 7308 4842
rect 7290 4842 7308 4860
rect 7290 4860 7308 4878
rect 7290 4878 7308 4896
rect 7290 4896 7308 4914
rect 7290 4914 7308 4932
rect 7290 4932 7308 4950
rect 7290 4950 7308 4968
rect 7290 4968 7308 4986
rect 7290 4986 7308 5004
rect 7290 5004 7308 5022
rect 7290 5022 7308 5040
rect 7290 5040 7308 5058
rect 7290 5058 7308 5076
rect 7290 5076 7308 5094
rect 7290 5094 7308 5112
rect 7290 5112 7308 5130
rect 7290 5130 7308 5148
rect 7290 5148 7308 5166
rect 7290 5166 7308 5184
rect 7290 5184 7308 5202
rect 7290 5202 7308 5220
rect 7290 5220 7308 5238
rect 7290 5238 7308 5256
rect 7290 5256 7308 5274
rect 7290 5274 7308 5292
rect 7290 5292 7308 5310
rect 7290 5310 7308 5328
rect 7290 5328 7308 5346
rect 7290 5346 7308 5364
rect 7290 5364 7308 5382
rect 7290 5382 7308 5400
rect 7290 5400 7308 5418
rect 7290 5418 7308 5436
rect 7290 5436 7308 5454
rect 7290 5454 7308 5472
rect 7290 5472 7308 5490
rect 7290 5490 7308 5508
rect 7290 5508 7308 5526
rect 7290 5526 7308 5544
rect 7290 5544 7308 5562
rect 7290 5562 7308 5580
rect 7290 5580 7308 5598
rect 7290 5598 7308 5616
rect 7290 5616 7308 5634
rect 7290 5634 7308 5652
rect 7290 5652 7308 5670
rect 7290 5670 7308 5688
rect 7290 5688 7308 5706
rect 7290 5706 7308 5724
rect 7290 5724 7308 5742
rect 7290 5742 7308 5760
rect 7290 5760 7308 5778
rect 7290 5778 7308 5796
rect 7290 5796 7308 5814
rect 7290 5814 7308 5832
rect 7290 5832 7308 5850
rect 7290 5850 7308 5868
rect 7290 5868 7308 5886
rect 7290 5886 7308 5904
rect 7290 5904 7308 5922
rect 7290 5922 7308 5940
rect 7290 5940 7308 5958
rect 7290 5958 7308 5976
rect 7290 5976 7308 5994
rect 7290 5994 7308 6012
rect 7290 6012 7308 6030
rect 7290 6030 7308 6048
rect 7290 6048 7308 6066
rect 7290 6066 7308 6084
rect 7290 6084 7308 6102
rect 7290 6102 7308 6120
rect 7290 6120 7308 6138
rect 7290 6138 7308 6156
rect 7290 6156 7308 6174
rect 7290 6174 7308 6192
rect 7290 6192 7308 6210
rect 7290 6210 7308 6228
rect 7290 6228 7308 6246
rect 7290 6246 7308 6264
rect 7290 6264 7308 6282
rect 7290 6282 7308 6300
rect 7290 6300 7308 6318
rect 7290 6318 7308 6336
rect 7290 6336 7308 6354
rect 7290 6354 7308 6372
rect 7290 6372 7308 6390
rect 7290 6390 7308 6408
rect 7290 6408 7308 6426
rect 7290 6426 7308 6444
rect 7290 6444 7308 6462
rect 7290 6462 7308 6480
rect 7290 6480 7308 6498
rect 7290 8874 7308 8892
rect 7290 8892 7308 8910
rect 7290 8910 7308 8928
rect 7290 8928 7308 8946
rect 7290 8946 7308 8964
rect 7290 8964 7308 8982
rect 7290 8982 7308 9000
rect 7290 9000 7308 9018
rect 7290 9018 7308 9036
rect 7290 9036 7308 9054
rect 7290 9054 7308 9072
rect 7290 9072 7308 9090
rect 7290 9090 7308 9108
rect 7290 9108 7308 9126
rect 7290 9126 7308 9144
rect 7290 9144 7308 9162
rect 7290 9162 7308 9180
rect 7290 9180 7308 9198
rect 7290 9198 7308 9216
rect 7290 9216 7308 9234
rect 7290 9234 7308 9252
rect 7290 9252 7308 9270
rect 7290 9270 7308 9288
rect 7290 9288 7308 9306
rect 7290 9306 7308 9324
rect 7290 9324 7308 9342
rect 7290 9342 7308 9360
rect 7290 9360 7308 9378
rect 7290 9378 7308 9396
rect 7290 9396 7308 9414
rect 7290 9414 7308 9432
rect 7290 9432 7308 9450
rect 7290 9450 7308 9468
rect 7290 9468 7308 9486
rect 7290 9486 7308 9504
rect 7290 9504 7308 9522
rect 7290 9522 7308 9540
rect 7290 9540 7308 9558
rect 7290 9558 7308 9576
rect 7290 9576 7308 9594
rect 7290 9594 7308 9612
rect 7290 9612 7308 9630
rect 7290 9630 7308 9648
rect 7308 1980 7326 1998
rect 7308 1998 7326 2016
rect 7308 2016 7326 2034
rect 7308 2034 7326 2052
rect 7308 2052 7326 2070
rect 7308 2070 7326 2088
rect 7308 2088 7326 2106
rect 7308 2106 7326 2124
rect 7308 2124 7326 2142
rect 7308 2142 7326 2160
rect 7308 2160 7326 2178
rect 7308 2178 7326 2196
rect 7308 2196 7326 2214
rect 7308 2214 7326 2232
rect 7308 2232 7326 2250
rect 7308 2250 7326 2268
rect 7308 2268 7326 2286
rect 7308 2286 7326 2304
rect 7308 2304 7326 2322
rect 7308 2322 7326 2340
rect 7308 2340 7326 2358
rect 7308 2358 7326 2376
rect 7308 2376 7326 2394
rect 7308 2394 7326 2412
rect 7308 2412 7326 2430
rect 7308 2430 7326 2448
rect 7308 2448 7326 2466
rect 7308 2466 7326 2484
rect 7308 2484 7326 2502
rect 7308 2502 7326 2520
rect 7308 2520 7326 2538
rect 7308 2538 7326 2556
rect 7308 2556 7326 2574
rect 7308 2574 7326 2592
rect 7308 2592 7326 2610
rect 7308 2610 7326 2628
rect 7308 2628 7326 2646
rect 7308 2646 7326 2664
rect 7308 2664 7326 2682
rect 7308 2682 7326 2700
rect 7308 2700 7326 2718
rect 7308 2718 7326 2736
rect 7308 2736 7326 2754
rect 7308 2754 7326 2772
rect 7308 2772 7326 2790
rect 7308 2790 7326 2808
rect 7308 2808 7326 2826
rect 7308 2826 7326 2844
rect 7308 2844 7326 2862
rect 7308 2862 7326 2880
rect 7308 2880 7326 2898
rect 7308 2898 7326 2916
rect 7308 2916 7326 2934
rect 7308 2934 7326 2952
rect 7308 2952 7326 2970
rect 7308 2970 7326 2988
rect 7308 2988 7326 3006
rect 7308 3006 7326 3024
rect 7308 3024 7326 3042
rect 7308 3042 7326 3060
rect 7308 3060 7326 3078
rect 7308 3078 7326 3096
rect 7308 3096 7326 3114
rect 7308 3114 7326 3132
rect 7308 3132 7326 3150
rect 7308 3150 7326 3168
rect 7308 3168 7326 3186
rect 7308 4410 7326 4428
rect 7308 4428 7326 4446
rect 7308 4446 7326 4464
rect 7308 4464 7326 4482
rect 7308 4482 7326 4500
rect 7308 4500 7326 4518
rect 7308 4518 7326 4536
rect 7308 4536 7326 4554
rect 7308 4554 7326 4572
rect 7308 4572 7326 4590
rect 7308 4590 7326 4608
rect 7308 4608 7326 4626
rect 7308 4626 7326 4644
rect 7308 4644 7326 4662
rect 7308 4662 7326 4680
rect 7308 4680 7326 4698
rect 7308 4698 7326 4716
rect 7308 4716 7326 4734
rect 7308 4734 7326 4752
rect 7308 4752 7326 4770
rect 7308 4770 7326 4788
rect 7308 4788 7326 4806
rect 7308 4806 7326 4824
rect 7308 4824 7326 4842
rect 7308 4842 7326 4860
rect 7308 4860 7326 4878
rect 7308 4878 7326 4896
rect 7308 4896 7326 4914
rect 7308 4914 7326 4932
rect 7308 4932 7326 4950
rect 7308 4950 7326 4968
rect 7308 4968 7326 4986
rect 7308 4986 7326 5004
rect 7308 5004 7326 5022
rect 7308 5022 7326 5040
rect 7308 5040 7326 5058
rect 7308 5058 7326 5076
rect 7308 5076 7326 5094
rect 7308 5094 7326 5112
rect 7308 5112 7326 5130
rect 7308 5130 7326 5148
rect 7308 5148 7326 5166
rect 7308 5166 7326 5184
rect 7308 5184 7326 5202
rect 7308 5202 7326 5220
rect 7308 5220 7326 5238
rect 7308 5238 7326 5256
rect 7308 5256 7326 5274
rect 7308 5274 7326 5292
rect 7308 5292 7326 5310
rect 7308 5310 7326 5328
rect 7308 5328 7326 5346
rect 7308 5346 7326 5364
rect 7308 5364 7326 5382
rect 7308 5382 7326 5400
rect 7308 5400 7326 5418
rect 7308 5418 7326 5436
rect 7308 5436 7326 5454
rect 7308 5454 7326 5472
rect 7308 5472 7326 5490
rect 7308 5490 7326 5508
rect 7308 5508 7326 5526
rect 7308 5526 7326 5544
rect 7308 5544 7326 5562
rect 7308 5562 7326 5580
rect 7308 5580 7326 5598
rect 7308 5598 7326 5616
rect 7308 5616 7326 5634
rect 7308 5634 7326 5652
rect 7308 5652 7326 5670
rect 7308 5670 7326 5688
rect 7308 5688 7326 5706
rect 7308 5706 7326 5724
rect 7308 5724 7326 5742
rect 7308 5742 7326 5760
rect 7308 5760 7326 5778
rect 7308 5778 7326 5796
rect 7308 5796 7326 5814
rect 7308 5814 7326 5832
rect 7308 5832 7326 5850
rect 7308 5850 7326 5868
rect 7308 5868 7326 5886
rect 7308 5886 7326 5904
rect 7308 5904 7326 5922
rect 7308 5922 7326 5940
rect 7308 5940 7326 5958
rect 7308 5958 7326 5976
rect 7308 5976 7326 5994
rect 7308 5994 7326 6012
rect 7308 6012 7326 6030
rect 7308 6030 7326 6048
rect 7308 6048 7326 6066
rect 7308 6066 7326 6084
rect 7308 6084 7326 6102
rect 7308 6102 7326 6120
rect 7308 6120 7326 6138
rect 7308 6138 7326 6156
rect 7308 6156 7326 6174
rect 7308 6174 7326 6192
rect 7308 6192 7326 6210
rect 7308 6210 7326 6228
rect 7308 6228 7326 6246
rect 7308 6246 7326 6264
rect 7308 6264 7326 6282
rect 7308 6282 7326 6300
rect 7308 6300 7326 6318
rect 7308 6318 7326 6336
rect 7308 6336 7326 6354
rect 7308 6354 7326 6372
rect 7308 6372 7326 6390
rect 7308 6390 7326 6408
rect 7308 6408 7326 6426
rect 7308 6426 7326 6444
rect 7308 6444 7326 6462
rect 7308 6462 7326 6480
rect 7308 6480 7326 6498
rect 7308 6498 7326 6516
rect 7308 8982 7326 9000
rect 7308 9000 7326 9018
rect 7308 9018 7326 9036
rect 7308 9036 7326 9054
rect 7308 9054 7326 9072
rect 7308 9072 7326 9090
rect 7308 9090 7326 9108
rect 7308 9108 7326 9126
rect 7308 9126 7326 9144
rect 7308 9144 7326 9162
rect 7308 9162 7326 9180
rect 7308 9180 7326 9198
rect 7308 9198 7326 9216
rect 7308 9216 7326 9234
rect 7308 9234 7326 9252
rect 7308 9252 7326 9270
rect 7308 9270 7326 9288
rect 7308 9288 7326 9306
rect 7308 9306 7326 9324
rect 7308 9324 7326 9342
rect 7308 9342 7326 9360
rect 7308 9360 7326 9378
rect 7308 9378 7326 9396
rect 7308 9396 7326 9414
rect 7308 9414 7326 9432
rect 7308 9432 7326 9450
rect 7308 9450 7326 9468
rect 7308 9468 7326 9486
rect 7308 9486 7326 9504
rect 7308 9504 7326 9522
rect 7326 1980 7344 1998
rect 7326 1998 7344 2016
rect 7326 2016 7344 2034
rect 7326 2034 7344 2052
rect 7326 2052 7344 2070
rect 7326 2070 7344 2088
rect 7326 2088 7344 2106
rect 7326 2106 7344 2124
rect 7326 2124 7344 2142
rect 7326 2142 7344 2160
rect 7326 2160 7344 2178
rect 7326 2178 7344 2196
rect 7326 2196 7344 2214
rect 7326 2214 7344 2232
rect 7326 2232 7344 2250
rect 7326 2250 7344 2268
rect 7326 2268 7344 2286
rect 7326 2286 7344 2304
rect 7326 2304 7344 2322
rect 7326 2322 7344 2340
rect 7326 2340 7344 2358
rect 7326 2358 7344 2376
rect 7326 2376 7344 2394
rect 7326 2394 7344 2412
rect 7326 2412 7344 2430
rect 7326 2430 7344 2448
rect 7326 2448 7344 2466
rect 7326 2466 7344 2484
rect 7326 2484 7344 2502
rect 7326 2502 7344 2520
rect 7326 2520 7344 2538
rect 7326 2538 7344 2556
rect 7326 2556 7344 2574
rect 7326 2574 7344 2592
rect 7326 2592 7344 2610
rect 7326 2610 7344 2628
rect 7326 2628 7344 2646
rect 7326 2646 7344 2664
rect 7326 2664 7344 2682
rect 7326 2682 7344 2700
rect 7326 2700 7344 2718
rect 7326 2718 7344 2736
rect 7326 2736 7344 2754
rect 7326 2754 7344 2772
rect 7326 2772 7344 2790
rect 7326 2790 7344 2808
rect 7326 2808 7344 2826
rect 7326 2826 7344 2844
rect 7326 2844 7344 2862
rect 7326 2862 7344 2880
rect 7326 2880 7344 2898
rect 7326 2898 7344 2916
rect 7326 2916 7344 2934
rect 7326 2934 7344 2952
rect 7326 2952 7344 2970
rect 7326 2970 7344 2988
rect 7326 2988 7344 3006
rect 7326 3006 7344 3024
rect 7326 3024 7344 3042
rect 7326 3042 7344 3060
rect 7326 3060 7344 3078
rect 7326 3078 7344 3096
rect 7326 3096 7344 3114
rect 7326 3114 7344 3132
rect 7326 3132 7344 3150
rect 7326 3150 7344 3168
rect 7326 3168 7344 3186
rect 7326 4428 7344 4446
rect 7326 4446 7344 4464
rect 7326 4464 7344 4482
rect 7326 4482 7344 4500
rect 7326 4500 7344 4518
rect 7326 4518 7344 4536
rect 7326 4536 7344 4554
rect 7326 4554 7344 4572
rect 7326 4572 7344 4590
rect 7326 4590 7344 4608
rect 7326 4608 7344 4626
rect 7326 4626 7344 4644
rect 7326 4644 7344 4662
rect 7326 4662 7344 4680
rect 7326 4680 7344 4698
rect 7326 4698 7344 4716
rect 7326 4716 7344 4734
rect 7326 4734 7344 4752
rect 7326 4752 7344 4770
rect 7326 4770 7344 4788
rect 7326 4788 7344 4806
rect 7326 4806 7344 4824
rect 7326 4824 7344 4842
rect 7326 4842 7344 4860
rect 7326 4860 7344 4878
rect 7326 4878 7344 4896
rect 7326 4896 7344 4914
rect 7326 4914 7344 4932
rect 7326 4932 7344 4950
rect 7326 4950 7344 4968
rect 7326 4968 7344 4986
rect 7326 4986 7344 5004
rect 7326 5004 7344 5022
rect 7326 5022 7344 5040
rect 7326 5040 7344 5058
rect 7326 5058 7344 5076
rect 7326 5076 7344 5094
rect 7326 5094 7344 5112
rect 7326 5112 7344 5130
rect 7326 5130 7344 5148
rect 7326 5148 7344 5166
rect 7326 5166 7344 5184
rect 7326 5184 7344 5202
rect 7326 5202 7344 5220
rect 7326 5220 7344 5238
rect 7326 5238 7344 5256
rect 7326 5256 7344 5274
rect 7326 5274 7344 5292
rect 7326 5292 7344 5310
rect 7326 5310 7344 5328
rect 7326 5328 7344 5346
rect 7326 5346 7344 5364
rect 7326 5364 7344 5382
rect 7326 5382 7344 5400
rect 7326 5400 7344 5418
rect 7326 5418 7344 5436
rect 7326 5436 7344 5454
rect 7326 5454 7344 5472
rect 7326 5472 7344 5490
rect 7326 5490 7344 5508
rect 7326 5508 7344 5526
rect 7326 5526 7344 5544
rect 7326 5544 7344 5562
rect 7326 5562 7344 5580
rect 7326 5580 7344 5598
rect 7326 5598 7344 5616
rect 7326 5616 7344 5634
rect 7326 5634 7344 5652
rect 7326 5652 7344 5670
rect 7326 5670 7344 5688
rect 7326 5688 7344 5706
rect 7326 5706 7344 5724
rect 7326 5724 7344 5742
rect 7326 5742 7344 5760
rect 7326 5760 7344 5778
rect 7326 5778 7344 5796
rect 7326 5796 7344 5814
rect 7326 5814 7344 5832
rect 7326 5832 7344 5850
rect 7326 5850 7344 5868
rect 7326 5868 7344 5886
rect 7326 5886 7344 5904
rect 7326 5904 7344 5922
rect 7326 5922 7344 5940
rect 7326 5940 7344 5958
rect 7326 5958 7344 5976
rect 7326 5976 7344 5994
rect 7326 5994 7344 6012
rect 7326 6012 7344 6030
rect 7326 6030 7344 6048
rect 7326 6048 7344 6066
rect 7326 6066 7344 6084
rect 7326 6084 7344 6102
rect 7326 6102 7344 6120
rect 7326 6120 7344 6138
rect 7326 6138 7344 6156
rect 7326 6156 7344 6174
rect 7326 6174 7344 6192
rect 7326 6192 7344 6210
rect 7326 6210 7344 6228
rect 7326 6228 7344 6246
rect 7326 6246 7344 6264
rect 7326 6264 7344 6282
rect 7326 6282 7344 6300
rect 7326 6300 7344 6318
rect 7326 6318 7344 6336
rect 7326 6336 7344 6354
rect 7326 6354 7344 6372
rect 7326 6372 7344 6390
rect 7326 6390 7344 6408
rect 7326 6408 7344 6426
rect 7326 6426 7344 6444
rect 7326 6444 7344 6462
rect 7326 6462 7344 6480
rect 7326 6480 7344 6498
rect 7326 6498 7344 6516
rect 7326 9198 7344 9216
rect 7326 9216 7344 9234
rect 7326 9234 7344 9252
rect 7326 9252 7344 9270
rect 7326 9270 7344 9288
rect 7344 1998 7362 2016
rect 7344 2016 7362 2034
rect 7344 2034 7362 2052
rect 7344 2052 7362 2070
rect 7344 2070 7362 2088
rect 7344 2088 7362 2106
rect 7344 2106 7362 2124
rect 7344 2124 7362 2142
rect 7344 2142 7362 2160
rect 7344 2160 7362 2178
rect 7344 2178 7362 2196
rect 7344 2196 7362 2214
rect 7344 2214 7362 2232
rect 7344 2232 7362 2250
rect 7344 2250 7362 2268
rect 7344 2268 7362 2286
rect 7344 2286 7362 2304
rect 7344 2304 7362 2322
rect 7344 2322 7362 2340
rect 7344 2340 7362 2358
rect 7344 2358 7362 2376
rect 7344 2376 7362 2394
rect 7344 2394 7362 2412
rect 7344 2412 7362 2430
rect 7344 2430 7362 2448
rect 7344 2448 7362 2466
rect 7344 2466 7362 2484
rect 7344 2484 7362 2502
rect 7344 2502 7362 2520
rect 7344 2520 7362 2538
rect 7344 2538 7362 2556
rect 7344 2556 7362 2574
rect 7344 2574 7362 2592
rect 7344 2592 7362 2610
rect 7344 2610 7362 2628
rect 7344 2628 7362 2646
rect 7344 2646 7362 2664
rect 7344 2664 7362 2682
rect 7344 2682 7362 2700
rect 7344 2700 7362 2718
rect 7344 2718 7362 2736
rect 7344 2736 7362 2754
rect 7344 2754 7362 2772
rect 7344 2772 7362 2790
rect 7344 2790 7362 2808
rect 7344 2808 7362 2826
rect 7344 2826 7362 2844
rect 7344 2844 7362 2862
rect 7344 2862 7362 2880
rect 7344 2880 7362 2898
rect 7344 2898 7362 2916
rect 7344 2916 7362 2934
rect 7344 2934 7362 2952
rect 7344 2952 7362 2970
rect 7344 2970 7362 2988
rect 7344 2988 7362 3006
rect 7344 3006 7362 3024
rect 7344 3024 7362 3042
rect 7344 3042 7362 3060
rect 7344 3060 7362 3078
rect 7344 3078 7362 3096
rect 7344 3096 7362 3114
rect 7344 3114 7362 3132
rect 7344 3132 7362 3150
rect 7344 3150 7362 3168
rect 7344 3168 7362 3186
rect 7344 4446 7362 4464
rect 7344 4464 7362 4482
rect 7344 4482 7362 4500
rect 7344 4500 7362 4518
rect 7344 4518 7362 4536
rect 7344 4536 7362 4554
rect 7344 4554 7362 4572
rect 7344 4572 7362 4590
rect 7344 4590 7362 4608
rect 7344 4608 7362 4626
rect 7344 4626 7362 4644
rect 7344 4644 7362 4662
rect 7344 4662 7362 4680
rect 7344 4680 7362 4698
rect 7344 4698 7362 4716
rect 7344 4716 7362 4734
rect 7344 4734 7362 4752
rect 7344 4752 7362 4770
rect 7344 4770 7362 4788
rect 7344 4788 7362 4806
rect 7344 4806 7362 4824
rect 7344 4824 7362 4842
rect 7344 4842 7362 4860
rect 7344 4860 7362 4878
rect 7344 4878 7362 4896
rect 7344 4896 7362 4914
rect 7344 4914 7362 4932
rect 7344 4932 7362 4950
rect 7344 4950 7362 4968
rect 7344 4968 7362 4986
rect 7344 4986 7362 5004
rect 7344 5004 7362 5022
rect 7344 5022 7362 5040
rect 7344 5040 7362 5058
rect 7344 5058 7362 5076
rect 7344 5076 7362 5094
rect 7344 5094 7362 5112
rect 7344 5112 7362 5130
rect 7344 5130 7362 5148
rect 7344 5148 7362 5166
rect 7344 5166 7362 5184
rect 7344 5184 7362 5202
rect 7344 5202 7362 5220
rect 7344 5220 7362 5238
rect 7344 5238 7362 5256
rect 7344 5256 7362 5274
rect 7344 5274 7362 5292
rect 7344 5292 7362 5310
rect 7344 5310 7362 5328
rect 7344 5328 7362 5346
rect 7344 5346 7362 5364
rect 7344 5364 7362 5382
rect 7344 5382 7362 5400
rect 7344 5400 7362 5418
rect 7344 5418 7362 5436
rect 7344 5436 7362 5454
rect 7344 5454 7362 5472
rect 7344 5472 7362 5490
rect 7344 5490 7362 5508
rect 7344 5508 7362 5526
rect 7344 5526 7362 5544
rect 7344 5544 7362 5562
rect 7344 5562 7362 5580
rect 7344 5580 7362 5598
rect 7344 5598 7362 5616
rect 7344 5616 7362 5634
rect 7344 5634 7362 5652
rect 7344 5652 7362 5670
rect 7344 5670 7362 5688
rect 7344 5688 7362 5706
rect 7344 5706 7362 5724
rect 7344 5724 7362 5742
rect 7344 5742 7362 5760
rect 7344 5760 7362 5778
rect 7344 5778 7362 5796
rect 7344 5796 7362 5814
rect 7344 5814 7362 5832
rect 7344 5832 7362 5850
rect 7344 5850 7362 5868
rect 7344 5868 7362 5886
rect 7344 5886 7362 5904
rect 7344 5904 7362 5922
rect 7344 5922 7362 5940
rect 7344 5940 7362 5958
rect 7344 5958 7362 5976
rect 7344 5976 7362 5994
rect 7344 5994 7362 6012
rect 7344 6012 7362 6030
rect 7344 6030 7362 6048
rect 7344 6048 7362 6066
rect 7344 6066 7362 6084
rect 7344 6084 7362 6102
rect 7344 6102 7362 6120
rect 7344 6120 7362 6138
rect 7344 6138 7362 6156
rect 7344 6156 7362 6174
rect 7344 6174 7362 6192
rect 7344 6192 7362 6210
rect 7344 6210 7362 6228
rect 7344 6228 7362 6246
rect 7344 6246 7362 6264
rect 7344 6264 7362 6282
rect 7344 6282 7362 6300
rect 7344 6300 7362 6318
rect 7344 6318 7362 6336
rect 7344 6336 7362 6354
rect 7344 6354 7362 6372
rect 7344 6372 7362 6390
rect 7344 6390 7362 6408
rect 7344 6408 7362 6426
rect 7344 6426 7362 6444
rect 7344 6444 7362 6462
rect 7344 6462 7362 6480
rect 7344 6480 7362 6498
rect 7344 6498 7362 6516
rect 7344 6516 7362 6534
rect 7362 1998 7380 2016
rect 7362 2016 7380 2034
rect 7362 2034 7380 2052
rect 7362 2052 7380 2070
rect 7362 2070 7380 2088
rect 7362 2088 7380 2106
rect 7362 2106 7380 2124
rect 7362 2124 7380 2142
rect 7362 2142 7380 2160
rect 7362 2160 7380 2178
rect 7362 2178 7380 2196
rect 7362 2196 7380 2214
rect 7362 2214 7380 2232
rect 7362 2232 7380 2250
rect 7362 2250 7380 2268
rect 7362 2268 7380 2286
rect 7362 2286 7380 2304
rect 7362 2304 7380 2322
rect 7362 2322 7380 2340
rect 7362 2340 7380 2358
rect 7362 2358 7380 2376
rect 7362 2376 7380 2394
rect 7362 2394 7380 2412
rect 7362 2412 7380 2430
rect 7362 2430 7380 2448
rect 7362 2448 7380 2466
rect 7362 2466 7380 2484
rect 7362 2484 7380 2502
rect 7362 2502 7380 2520
rect 7362 2520 7380 2538
rect 7362 2538 7380 2556
rect 7362 2556 7380 2574
rect 7362 2574 7380 2592
rect 7362 2592 7380 2610
rect 7362 2610 7380 2628
rect 7362 2628 7380 2646
rect 7362 2646 7380 2664
rect 7362 2664 7380 2682
rect 7362 2682 7380 2700
rect 7362 2700 7380 2718
rect 7362 2718 7380 2736
rect 7362 2736 7380 2754
rect 7362 2754 7380 2772
rect 7362 2772 7380 2790
rect 7362 2790 7380 2808
rect 7362 2808 7380 2826
rect 7362 2826 7380 2844
rect 7362 2844 7380 2862
rect 7362 2862 7380 2880
rect 7362 2880 7380 2898
rect 7362 2898 7380 2916
rect 7362 2916 7380 2934
rect 7362 2934 7380 2952
rect 7362 2952 7380 2970
rect 7362 2970 7380 2988
rect 7362 2988 7380 3006
rect 7362 3006 7380 3024
rect 7362 3024 7380 3042
rect 7362 3042 7380 3060
rect 7362 3060 7380 3078
rect 7362 3078 7380 3096
rect 7362 3096 7380 3114
rect 7362 3114 7380 3132
rect 7362 3132 7380 3150
rect 7362 3150 7380 3168
rect 7362 3168 7380 3186
rect 7362 3186 7380 3204
rect 7362 4464 7380 4482
rect 7362 4482 7380 4500
rect 7362 4500 7380 4518
rect 7362 4518 7380 4536
rect 7362 4536 7380 4554
rect 7362 4554 7380 4572
rect 7362 4572 7380 4590
rect 7362 4590 7380 4608
rect 7362 4608 7380 4626
rect 7362 4626 7380 4644
rect 7362 4644 7380 4662
rect 7362 4662 7380 4680
rect 7362 4680 7380 4698
rect 7362 4698 7380 4716
rect 7362 4716 7380 4734
rect 7362 4734 7380 4752
rect 7362 4752 7380 4770
rect 7362 4770 7380 4788
rect 7362 4788 7380 4806
rect 7362 4806 7380 4824
rect 7362 4824 7380 4842
rect 7362 4842 7380 4860
rect 7362 4860 7380 4878
rect 7362 4878 7380 4896
rect 7362 4896 7380 4914
rect 7362 4914 7380 4932
rect 7362 4932 7380 4950
rect 7362 4950 7380 4968
rect 7362 4968 7380 4986
rect 7362 4986 7380 5004
rect 7362 5004 7380 5022
rect 7362 5022 7380 5040
rect 7362 5040 7380 5058
rect 7362 5058 7380 5076
rect 7362 5076 7380 5094
rect 7362 5094 7380 5112
rect 7362 5112 7380 5130
rect 7362 5130 7380 5148
rect 7362 5148 7380 5166
rect 7362 5166 7380 5184
rect 7362 5184 7380 5202
rect 7362 5202 7380 5220
rect 7362 5220 7380 5238
rect 7362 5238 7380 5256
rect 7362 5256 7380 5274
rect 7362 5274 7380 5292
rect 7362 5292 7380 5310
rect 7362 5310 7380 5328
rect 7362 5328 7380 5346
rect 7362 5346 7380 5364
rect 7362 5364 7380 5382
rect 7362 5382 7380 5400
rect 7362 5400 7380 5418
rect 7362 5418 7380 5436
rect 7362 5436 7380 5454
rect 7362 5454 7380 5472
rect 7362 5472 7380 5490
rect 7362 5490 7380 5508
rect 7362 5508 7380 5526
rect 7362 5526 7380 5544
rect 7362 5544 7380 5562
rect 7362 5562 7380 5580
rect 7362 5580 7380 5598
rect 7362 5598 7380 5616
rect 7362 5616 7380 5634
rect 7362 5634 7380 5652
rect 7362 5652 7380 5670
rect 7362 5670 7380 5688
rect 7362 5688 7380 5706
rect 7362 5706 7380 5724
rect 7362 5724 7380 5742
rect 7362 5742 7380 5760
rect 7362 5760 7380 5778
rect 7362 5778 7380 5796
rect 7362 5796 7380 5814
rect 7362 5814 7380 5832
rect 7362 5832 7380 5850
rect 7362 5850 7380 5868
rect 7362 5868 7380 5886
rect 7362 5886 7380 5904
rect 7362 5904 7380 5922
rect 7362 5922 7380 5940
rect 7362 5940 7380 5958
rect 7362 5958 7380 5976
rect 7362 5976 7380 5994
rect 7362 5994 7380 6012
rect 7362 6012 7380 6030
rect 7362 6030 7380 6048
rect 7362 6048 7380 6066
rect 7362 6066 7380 6084
rect 7362 6084 7380 6102
rect 7362 6102 7380 6120
rect 7362 6120 7380 6138
rect 7362 6138 7380 6156
rect 7362 6156 7380 6174
rect 7362 6174 7380 6192
rect 7362 6192 7380 6210
rect 7362 6210 7380 6228
rect 7362 6228 7380 6246
rect 7362 6246 7380 6264
rect 7362 6264 7380 6282
rect 7362 6282 7380 6300
rect 7362 6300 7380 6318
rect 7362 6318 7380 6336
rect 7362 6336 7380 6354
rect 7362 6354 7380 6372
rect 7362 6372 7380 6390
rect 7362 6390 7380 6408
rect 7362 6408 7380 6426
rect 7362 6426 7380 6444
rect 7362 6444 7380 6462
rect 7362 6462 7380 6480
rect 7362 6480 7380 6498
rect 7362 6498 7380 6516
rect 7362 6516 7380 6534
rect 7362 6534 7380 6552
rect 7380 2016 7398 2034
rect 7380 2034 7398 2052
rect 7380 2052 7398 2070
rect 7380 2070 7398 2088
rect 7380 2088 7398 2106
rect 7380 2106 7398 2124
rect 7380 2124 7398 2142
rect 7380 2142 7398 2160
rect 7380 2160 7398 2178
rect 7380 2178 7398 2196
rect 7380 2196 7398 2214
rect 7380 2214 7398 2232
rect 7380 2232 7398 2250
rect 7380 2250 7398 2268
rect 7380 2268 7398 2286
rect 7380 2286 7398 2304
rect 7380 2304 7398 2322
rect 7380 2322 7398 2340
rect 7380 2340 7398 2358
rect 7380 2358 7398 2376
rect 7380 2376 7398 2394
rect 7380 2394 7398 2412
rect 7380 2412 7398 2430
rect 7380 2430 7398 2448
rect 7380 2448 7398 2466
rect 7380 2466 7398 2484
rect 7380 2484 7398 2502
rect 7380 2502 7398 2520
rect 7380 2520 7398 2538
rect 7380 2538 7398 2556
rect 7380 2556 7398 2574
rect 7380 2574 7398 2592
rect 7380 2592 7398 2610
rect 7380 2610 7398 2628
rect 7380 2628 7398 2646
rect 7380 2646 7398 2664
rect 7380 2664 7398 2682
rect 7380 2682 7398 2700
rect 7380 2700 7398 2718
rect 7380 2718 7398 2736
rect 7380 2736 7398 2754
rect 7380 2754 7398 2772
rect 7380 2772 7398 2790
rect 7380 2790 7398 2808
rect 7380 2808 7398 2826
rect 7380 2826 7398 2844
rect 7380 2844 7398 2862
rect 7380 2862 7398 2880
rect 7380 2880 7398 2898
rect 7380 2898 7398 2916
rect 7380 2916 7398 2934
rect 7380 2934 7398 2952
rect 7380 2952 7398 2970
rect 7380 2970 7398 2988
rect 7380 2988 7398 3006
rect 7380 3006 7398 3024
rect 7380 3024 7398 3042
rect 7380 3042 7398 3060
rect 7380 3060 7398 3078
rect 7380 3078 7398 3096
rect 7380 3096 7398 3114
rect 7380 3114 7398 3132
rect 7380 3132 7398 3150
rect 7380 3150 7398 3168
rect 7380 3168 7398 3186
rect 7380 3186 7398 3204
rect 7380 4500 7398 4518
rect 7380 4518 7398 4536
rect 7380 4536 7398 4554
rect 7380 4554 7398 4572
rect 7380 4572 7398 4590
rect 7380 4590 7398 4608
rect 7380 4608 7398 4626
rect 7380 4626 7398 4644
rect 7380 4644 7398 4662
rect 7380 4662 7398 4680
rect 7380 4680 7398 4698
rect 7380 4698 7398 4716
rect 7380 4716 7398 4734
rect 7380 4734 7398 4752
rect 7380 4752 7398 4770
rect 7380 4770 7398 4788
rect 7380 4788 7398 4806
rect 7380 4806 7398 4824
rect 7380 4824 7398 4842
rect 7380 4842 7398 4860
rect 7380 4860 7398 4878
rect 7380 4878 7398 4896
rect 7380 4896 7398 4914
rect 7380 4914 7398 4932
rect 7380 4932 7398 4950
rect 7380 4950 7398 4968
rect 7380 4968 7398 4986
rect 7380 4986 7398 5004
rect 7380 5004 7398 5022
rect 7380 5022 7398 5040
rect 7380 5040 7398 5058
rect 7380 5058 7398 5076
rect 7380 5076 7398 5094
rect 7380 5094 7398 5112
rect 7380 5112 7398 5130
rect 7380 5130 7398 5148
rect 7380 5148 7398 5166
rect 7380 5166 7398 5184
rect 7380 5184 7398 5202
rect 7380 5202 7398 5220
rect 7380 5220 7398 5238
rect 7380 5238 7398 5256
rect 7380 5256 7398 5274
rect 7380 5274 7398 5292
rect 7380 5292 7398 5310
rect 7380 5310 7398 5328
rect 7380 5328 7398 5346
rect 7380 5346 7398 5364
rect 7380 5364 7398 5382
rect 7380 5382 7398 5400
rect 7380 5400 7398 5418
rect 7380 5418 7398 5436
rect 7380 5436 7398 5454
rect 7380 5454 7398 5472
rect 7380 5472 7398 5490
rect 7380 5490 7398 5508
rect 7380 5508 7398 5526
rect 7380 5526 7398 5544
rect 7380 5544 7398 5562
rect 7380 5562 7398 5580
rect 7380 5580 7398 5598
rect 7380 5598 7398 5616
rect 7380 5616 7398 5634
rect 7380 5634 7398 5652
rect 7380 5652 7398 5670
rect 7380 5670 7398 5688
rect 7380 5688 7398 5706
rect 7380 5706 7398 5724
rect 7380 5724 7398 5742
rect 7380 5742 7398 5760
rect 7380 5760 7398 5778
rect 7380 5778 7398 5796
rect 7380 5796 7398 5814
rect 7380 5814 7398 5832
rect 7380 5832 7398 5850
rect 7380 5850 7398 5868
rect 7380 5868 7398 5886
rect 7380 5886 7398 5904
rect 7380 5904 7398 5922
rect 7380 5922 7398 5940
rect 7380 5940 7398 5958
rect 7380 5958 7398 5976
rect 7380 5976 7398 5994
rect 7380 5994 7398 6012
rect 7380 6012 7398 6030
rect 7380 6030 7398 6048
rect 7380 6048 7398 6066
rect 7380 6066 7398 6084
rect 7380 6084 7398 6102
rect 7380 6102 7398 6120
rect 7380 6120 7398 6138
rect 7380 6138 7398 6156
rect 7380 6156 7398 6174
rect 7380 6174 7398 6192
rect 7380 6192 7398 6210
rect 7380 6210 7398 6228
rect 7380 6228 7398 6246
rect 7380 6246 7398 6264
rect 7380 6264 7398 6282
rect 7380 6282 7398 6300
rect 7380 6300 7398 6318
rect 7380 6318 7398 6336
rect 7380 6336 7398 6354
rect 7380 6354 7398 6372
rect 7380 6372 7398 6390
rect 7380 6390 7398 6408
rect 7380 6408 7398 6426
rect 7380 6426 7398 6444
rect 7380 6444 7398 6462
rect 7380 6462 7398 6480
rect 7380 6480 7398 6498
rect 7380 6498 7398 6516
rect 7380 6516 7398 6534
rect 7380 6534 7398 6552
rect 7380 6552 7398 6570
rect 7398 2034 7416 2052
rect 7398 2052 7416 2070
rect 7398 2070 7416 2088
rect 7398 2088 7416 2106
rect 7398 2106 7416 2124
rect 7398 2124 7416 2142
rect 7398 2142 7416 2160
rect 7398 2160 7416 2178
rect 7398 2178 7416 2196
rect 7398 2196 7416 2214
rect 7398 2214 7416 2232
rect 7398 2232 7416 2250
rect 7398 2250 7416 2268
rect 7398 2268 7416 2286
rect 7398 2286 7416 2304
rect 7398 2304 7416 2322
rect 7398 2322 7416 2340
rect 7398 2340 7416 2358
rect 7398 2358 7416 2376
rect 7398 2376 7416 2394
rect 7398 2394 7416 2412
rect 7398 2412 7416 2430
rect 7398 2430 7416 2448
rect 7398 2448 7416 2466
rect 7398 2466 7416 2484
rect 7398 2484 7416 2502
rect 7398 2502 7416 2520
rect 7398 2520 7416 2538
rect 7398 2538 7416 2556
rect 7398 2556 7416 2574
rect 7398 2574 7416 2592
rect 7398 2592 7416 2610
rect 7398 2610 7416 2628
rect 7398 2628 7416 2646
rect 7398 2646 7416 2664
rect 7398 2664 7416 2682
rect 7398 2682 7416 2700
rect 7398 2700 7416 2718
rect 7398 2718 7416 2736
rect 7398 2736 7416 2754
rect 7398 2754 7416 2772
rect 7398 2772 7416 2790
rect 7398 2790 7416 2808
rect 7398 2808 7416 2826
rect 7398 2826 7416 2844
rect 7398 2844 7416 2862
rect 7398 2862 7416 2880
rect 7398 2880 7416 2898
rect 7398 2898 7416 2916
rect 7398 2916 7416 2934
rect 7398 2934 7416 2952
rect 7398 2952 7416 2970
rect 7398 2970 7416 2988
rect 7398 2988 7416 3006
rect 7398 3006 7416 3024
rect 7398 3024 7416 3042
rect 7398 3042 7416 3060
rect 7398 3060 7416 3078
rect 7398 3078 7416 3096
rect 7398 3096 7416 3114
rect 7398 3114 7416 3132
rect 7398 3132 7416 3150
rect 7398 3150 7416 3168
rect 7398 3168 7416 3186
rect 7398 3186 7416 3204
rect 7398 4518 7416 4536
rect 7398 4536 7416 4554
rect 7398 4554 7416 4572
rect 7398 4572 7416 4590
rect 7398 4590 7416 4608
rect 7398 4608 7416 4626
rect 7398 4626 7416 4644
rect 7398 4644 7416 4662
rect 7398 4662 7416 4680
rect 7398 4680 7416 4698
rect 7398 4698 7416 4716
rect 7398 4716 7416 4734
rect 7398 4734 7416 4752
rect 7398 4752 7416 4770
rect 7398 4770 7416 4788
rect 7398 4788 7416 4806
rect 7398 4806 7416 4824
rect 7398 4824 7416 4842
rect 7398 4842 7416 4860
rect 7398 4860 7416 4878
rect 7398 4878 7416 4896
rect 7398 4896 7416 4914
rect 7398 4914 7416 4932
rect 7398 4932 7416 4950
rect 7398 4950 7416 4968
rect 7398 4968 7416 4986
rect 7398 4986 7416 5004
rect 7398 5004 7416 5022
rect 7398 5022 7416 5040
rect 7398 5040 7416 5058
rect 7398 5058 7416 5076
rect 7398 5076 7416 5094
rect 7398 5094 7416 5112
rect 7398 5112 7416 5130
rect 7398 5130 7416 5148
rect 7398 5148 7416 5166
rect 7398 5166 7416 5184
rect 7398 5184 7416 5202
rect 7398 5202 7416 5220
rect 7398 5220 7416 5238
rect 7398 5238 7416 5256
rect 7398 5256 7416 5274
rect 7398 5274 7416 5292
rect 7398 5292 7416 5310
rect 7398 5310 7416 5328
rect 7398 5328 7416 5346
rect 7398 5346 7416 5364
rect 7398 5364 7416 5382
rect 7398 5382 7416 5400
rect 7398 5400 7416 5418
rect 7398 5418 7416 5436
rect 7398 5436 7416 5454
rect 7398 5454 7416 5472
rect 7398 5472 7416 5490
rect 7398 5490 7416 5508
rect 7398 5508 7416 5526
rect 7398 5526 7416 5544
rect 7398 5544 7416 5562
rect 7398 5562 7416 5580
rect 7398 5580 7416 5598
rect 7398 5598 7416 5616
rect 7398 5616 7416 5634
rect 7398 5634 7416 5652
rect 7398 5652 7416 5670
rect 7398 5670 7416 5688
rect 7398 5688 7416 5706
rect 7398 5706 7416 5724
rect 7398 5724 7416 5742
rect 7398 5742 7416 5760
rect 7398 5760 7416 5778
rect 7398 5778 7416 5796
rect 7398 5796 7416 5814
rect 7398 5814 7416 5832
rect 7398 5832 7416 5850
rect 7398 5850 7416 5868
rect 7398 5868 7416 5886
rect 7398 5886 7416 5904
rect 7398 5904 7416 5922
rect 7398 5922 7416 5940
rect 7398 5940 7416 5958
rect 7398 5958 7416 5976
rect 7398 5976 7416 5994
rect 7398 5994 7416 6012
rect 7398 6012 7416 6030
rect 7398 6030 7416 6048
rect 7398 6048 7416 6066
rect 7398 6066 7416 6084
rect 7398 6084 7416 6102
rect 7398 6102 7416 6120
rect 7398 6120 7416 6138
rect 7398 6138 7416 6156
rect 7398 6156 7416 6174
rect 7398 6174 7416 6192
rect 7398 6192 7416 6210
rect 7398 6210 7416 6228
rect 7398 6228 7416 6246
rect 7398 6246 7416 6264
rect 7398 6264 7416 6282
rect 7398 6282 7416 6300
rect 7398 6300 7416 6318
rect 7398 6318 7416 6336
rect 7398 6336 7416 6354
rect 7398 6354 7416 6372
rect 7398 6372 7416 6390
rect 7398 6390 7416 6408
rect 7398 6408 7416 6426
rect 7398 6426 7416 6444
rect 7398 6444 7416 6462
rect 7398 6462 7416 6480
rect 7398 6480 7416 6498
rect 7398 6498 7416 6516
rect 7398 6516 7416 6534
rect 7398 6534 7416 6552
rect 7398 6552 7416 6570
rect 7398 6570 7416 6588
rect 7416 2034 7434 2052
rect 7416 2052 7434 2070
rect 7416 2070 7434 2088
rect 7416 2088 7434 2106
rect 7416 2106 7434 2124
rect 7416 2124 7434 2142
rect 7416 2142 7434 2160
rect 7416 2160 7434 2178
rect 7416 2178 7434 2196
rect 7416 2196 7434 2214
rect 7416 2214 7434 2232
rect 7416 2232 7434 2250
rect 7416 2250 7434 2268
rect 7416 2268 7434 2286
rect 7416 2286 7434 2304
rect 7416 2304 7434 2322
rect 7416 2322 7434 2340
rect 7416 2340 7434 2358
rect 7416 2358 7434 2376
rect 7416 2376 7434 2394
rect 7416 2394 7434 2412
rect 7416 2412 7434 2430
rect 7416 2430 7434 2448
rect 7416 2448 7434 2466
rect 7416 2466 7434 2484
rect 7416 2484 7434 2502
rect 7416 2502 7434 2520
rect 7416 2520 7434 2538
rect 7416 2538 7434 2556
rect 7416 2556 7434 2574
rect 7416 2574 7434 2592
rect 7416 2592 7434 2610
rect 7416 2610 7434 2628
rect 7416 2628 7434 2646
rect 7416 2646 7434 2664
rect 7416 2664 7434 2682
rect 7416 2682 7434 2700
rect 7416 2700 7434 2718
rect 7416 2718 7434 2736
rect 7416 2736 7434 2754
rect 7416 2754 7434 2772
rect 7416 2772 7434 2790
rect 7416 2790 7434 2808
rect 7416 2808 7434 2826
rect 7416 2826 7434 2844
rect 7416 2844 7434 2862
rect 7416 2862 7434 2880
rect 7416 2880 7434 2898
rect 7416 2898 7434 2916
rect 7416 2916 7434 2934
rect 7416 2934 7434 2952
rect 7416 2952 7434 2970
rect 7416 2970 7434 2988
rect 7416 2988 7434 3006
rect 7416 3006 7434 3024
rect 7416 3024 7434 3042
rect 7416 3042 7434 3060
rect 7416 3060 7434 3078
rect 7416 3078 7434 3096
rect 7416 3096 7434 3114
rect 7416 3114 7434 3132
rect 7416 3132 7434 3150
rect 7416 3150 7434 3168
rect 7416 3168 7434 3186
rect 7416 3186 7434 3204
rect 7416 4536 7434 4554
rect 7416 4554 7434 4572
rect 7416 4572 7434 4590
rect 7416 4590 7434 4608
rect 7416 4608 7434 4626
rect 7416 4626 7434 4644
rect 7416 4644 7434 4662
rect 7416 4662 7434 4680
rect 7416 4680 7434 4698
rect 7416 4698 7434 4716
rect 7416 4716 7434 4734
rect 7416 4734 7434 4752
rect 7416 4752 7434 4770
rect 7416 4770 7434 4788
rect 7416 4788 7434 4806
rect 7416 4806 7434 4824
rect 7416 4824 7434 4842
rect 7416 4842 7434 4860
rect 7416 4860 7434 4878
rect 7416 4878 7434 4896
rect 7416 4896 7434 4914
rect 7416 4914 7434 4932
rect 7416 4932 7434 4950
rect 7416 4950 7434 4968
rect 7416 4968 7434 4986
rect 7416 4986 7434 5004
rect 7416 5004 7434 5022
rect 7416 5022 7434 5040
rect 7416 5040 7434 5058
rect 7416 5058 7434 5076
rect 7416 5076 7434 5094
rect 7416 5094 7434 5112
rect 7416 5112 7434 5130
rect 7416 5130 7434 5148
rect 7416 5148 7434 5166
rect 7416 5166 7434 5184
rect 7416 5184 7434 5202
rect 7416 5202 7434 5220
rect 7416 5220 7434 5238
rect 7416 5238 7434 5256
rect 7416 5256 7434 5274
rect 7416 5274 7434 5292
rect 7416 5292 7434 5310
rect 7416 5310 7434 5328
rect 7416 5328 7434 5346
rect 7416 5346 7434 5364
rect 7416 5364 7434 5382
rect 7416 5382 7434 5400
rect 7416 5400 7434 5418
rect 7416 5418 7434 5436
rect 7416 5436 7434 5454
rect 7416 5454 7434 5472
rect 7416 5472 7434 5490
rect 7416 5490 7434 5508
rect 7416 5508 7434 5526
rect 7416 5526 7434 5544
rect 7416 5544 7434 5562
rect 7416 5562 7434 5580
rect 7416 5580 7434 5598
rect 7416 5598 7434 5616
rect 7416 5616 7434 5634
rect 7416 5634 7434 5652
rect 7416 5652 7434 5670
rect 7416 5670 7434 5688
rect 7416 5688 7434 5706
rect 7416 5706 7434 5724
rect 7416 5724 7434 5742
rect 7416 5742 7434 5760
rect 7416 5760 7434 5778
rect 7416 5778 7434 5796
rect 7416 5796 7434 5814
rect 7416 5814 7434 5832
rect 7416 5832 7434 5850
rect 7416 5850 7434 5868
rect 7416 5868 7434 5886
rect 7416 5886 7434 5904
rect 7416 5904 7434 5922
rect 7416 5922 7434 5940
rect 7416 5940 7434 5958
rect 7416 5958 7434 5976
rect 7416 5976 7434 5994
rect 7416 5994 7434 6012
rect 7416 6012 7434 6030
rect 7416 6030 7434 6048
rect 7416 6048 7434 6066
rect 7416 6066 7434 6084
rect 7416 6084 7434 6102
rect 7416 6102 7434 6120
rect 7416 6120 7434 6138
rect 7416 6138 7434 6156
rect 7416 6156 7434 6174
rect 7416 6174 7434 6192
rect 7416 6192 7434 6210
rect 7416 6210 7434 6228
rect 7416 6228 7434 6246
rect 7416 6246 7434 6264
rect 7416 6264 7434 6282
rect 7416 6282 7434 6300
rect 7416 6300 7434 6318
rect 7416 6318 7434 6336
rect 7416 6336 7434 6354
rect 7416 6354 7434 6372
rect 7416 6372 7434 6390
rect 7416 6390 7434 6408
rect 7416 6408 7434 6426
rect 7416 6426 7434 6444
rect 7416 6444 7434 6462
rect 7416 6462 7434 6480
rect 7416 6480 7434 6498
rect 7416 6498 7434 6516
rect 7416 6516 7434 6534
rect 7416 6534 7434 6552
rect 7416 6552 7434 6570
rect 7416 6570 7434 6588
rect 7434 2052 7452 2070
rect 7434 2070 7452 2088
rect 7434 2088 7452 2106
rect 7434 2106 7452 2124
rect 7434 2124 7452 2142
rect 7434 2142 7452 2160
rect 7434 2160 7452 2178
rect 7434 2178 7452 2196
rect 7434 2196 7452 2214
rect 7434 2214 7452 2232
rect 7434 2232 7452 2250
rect 7434 2250 7452 2268
rect 7434 2268 7452 2286
rect 7434 2286 7452 2304
rect 7434 2304 7452 2322
rect 7434 2322 7452 2340
rect 7434 2340 7452 2358
rect 7434 2358 7452 2376
rect 7434 2376 7452 2394
rect 7434 2394 7452 2412
rect 7434 2412 7452 2430
rect 7434 2430 7452 2448
rect 7434 2448 7452 2466
rect 7434 2466 7452 2484
rect 7434 2484 7452 2502
rect 7434 2502 7452 2520
rect 7434 2520 7452 2538
rect 7434 2538 7452 2556
rect 7434 2556 7452 2574
rect 7434 2574 7452 2592
rect 7434 2592 7452 2610
rect 7434 2610 7452 2628
rect 7434 2628 7452 2646
rect 7434 2646 7452 2664
rect 7434 2664 7452 2682
rect 7434 2682 7452 2700
rect 7434 2700 7452 2718
rect 7434 2718 7452 2736
rect 7434 2736 7452 2754
rect 7434 2754 7452 2772
rect 7434 2772 7452 2790
rect 7434 2790 7452 2808
rect 7434 2808 7452 2826
rect 7434 2826 7452 2844
rect 7434 2844 7452 2862
rect 7434 2862 7452 2880
rect 7434 2880 7452 2898
rect 7434 2898 7452 2916
rect 7434 2916 7452 2934
rect 7434 2934 7452 2952
rect 7434 2952 7452 2970
rect 7434 2970 7452 2988
rect 7434 2988 7452 3006
rect 7434 3006 7452 3024
rect 7434 3024 7452 3042
rect 7434 3042 7452 3060
rect 7434 3060 7452 3078
rect 7434 3078 7452 3096
rect 7434 3096 7452 3114
rect 7434 3114 7452 3132
rect 7434 3132 7452 3150
rect 7434 3150 7452 3168
rect 7434 3168 7452 3186
rect 7434 3186 7452 3204
rect 7434 3204 7452 3222
rect 7434 4554 7452 4572
rect 7434 4572 7452 4590
rect 7434 4590 7452 4608
rect 7434 4608 7452 4626
rect 7434 4626 7452 4644
rect 7434 4644 7452 4662
rect 7434 4662 7452 4680
rect 7434 4680 7452 4698
rect 7434 4698 7452 4716
rect 7434 4716 7452 4734
rect 7434 4734 7452 4752
rect 7434 4752 7452 4770
rect 7434 4770 7452 4788
rect 7434 4788 7452 4806
rect 7434 4806 7452 4824
rect 7434 4824 7452 4842
rect 7434 4842 7452 4860
rect 7434 4860 7452 4878
rect 7434 4878 7452 4896
rect 7434 4896 7452 4914
rect 7434 4914 7452 4932
rect 7434 4932 7452 4950
rect 7434 4950 7452 4968
rect 7434 4968 7452 4986
rect 7434 4986 7452 5004
rect 7434 5004 7452 5022
rect 7434 5022 7452 5040
rect 7434 5040 7452 5058
rect 7434 5058 7452 5076
rect 7434 5076 7452 5094
rect 7434 5094 7452 5112
rect 7434 5112 7452 5130
rect 7434 5130 7452 5148
rect 7434 5148 7452 5166
rect 7434 5166 7452 5184
rect 7434 5184 7452 5202
rect 7434 5202 7452 5220
rect 7434 5220 7452 5238
rect 7434 5238 7452 5256
rect 7434 5256 7452 5274
rect 7434 5274 7452 5292
rect 7434 5292 7452 5310
rect 7434 5310 7452 5328
rect 7434 5328 7452 5346
rect 7434 5346 7452 5364
rect 7434 5364 7452 5382
rect 7434 5382 7452 5400
rect 7434 5400 7452 5418
rect 7434 5418 7452 5436
rect 7434 5436 7452 5454
rect 7434 5454 7452 5472
rect 7434 5472 7452 5490
rect 7434 5490 7452 5508
rect 7434 5508 7452 5526
rect 7434 5526 7452 5544
rect 7434 5544 7452 5562
rect 7434 5562 7452 5580
rect 7434 5580 7452 5598
rect 7434 5598 7452 5616
rect 7434 5616 7452 5634
rect 7434 5634 7452 5652
rect 7434 5652 7452 5670
rect 7434 5670 7452 5688
rect 7434 5688 7452 5706
rect 7434 5706 7452 5724
rect 7434 5724 7452 5742
rect 7434 5742 7452 5760
rect 7434 5760 7452 5778
rect 7434 5778 7452 5796
rect 7434 5796 7452 5814
rect 7434 5814 7452 5832
rect 7434 5832 7452 5850
rect 7434 5850 7452 5868
rect 7434 5868 7452 5886
rect 7434 5886 7452 5904
rect 7434 5904 7452 5922
rect 7434 5922 7452 5940
rect 7434 5940 7452 5958
rect 7434 5958 7452 5976
rect 7434 5976 7452 5994
rect 7434 5994 7452 6012
rect 7434 6012 7452 6030
rect 7434 6030 7452 6048
rect 7434 6048 7452 6066
rect 7434 6066 7452 6084
rect 7434 6084 7452 6102
rect 7434 6102 7452 6120
rect 7434 6120 7452 6138
rect 7434 6138 7452 6156
rect 7434 6156 7452 6174
rect 7434 6174 7452 6192
rect 7434 6192 7452 6210
rect 7434 6210 7452 6228
rect 7434 6228 7452 6246
rect 7434 6246 7452 6264
rect 7434 6264 7452 6282
rect 7434 6282 7452 6300
rect 7434 6300 7452 6318
rect 7434 6318 7452 6336
rect 7434 6336 7452 6354
rect 7434 6354 7452 6372
rect 7434 6372 7452 6390
rect 7434 6390 7452 6408
rect 7434 6408 7452 6426
rect 7434 6426 7452 6444
rect 7434 6444 7452 6462
rect 7434 6462 7452 6480
rect 7434 6480 7452 6498
rect 7434 6498 7452 6516
rect 7434 6516 7452 6534
rect 7434 6534 7452 6552
rect 7434 6552 7452 6570
rect 7434 6570 7452 6588
rect 7434 6588 7452 6606
rect 7452 2052 7470 2070
rect 7452 2070 7470 2088
rect 7452 2088 7470 2106
rect 7452 2106 7470 2124
rect 7452 2124 7470 2142
rect 7452 2142 7470 2160
rect 7452 2160 7470 2178
rect 7452 2178 7470 2196
rect 7452 2196 7470 2214
rect 7452 2214 7470 2232
rect 7452 2232 7470 2250
rect 7452 2250 7470 2268
rect 7452 2268 7470 2286
rect 7452 2286 7470 2304
rect 7452 2304 7470 2322
rect 7452 2322 7470 2340
rect 7452 2340 7470 2358
rect 7452 2358 7470 2376
rect 7452 2376 7470 2394
rect 7452 2394 7470 2412
rect 7452 2412 7470 2430
rect 7452 2430 7470 2448
rect 7452 2448 7470 2466
rect 7452 2466 7470 2484
rect 7452 2484 7470 2502
rect 7452 2502 7470 2520
rect 7452 2520 7470 2538
rect 7452 2538 7470 2556
rect 7452 2556 7470 2574
rect 7452 2574 7470 2592
rect 7452 2592 7470 2610
rect 7452 2610 7470 2628
rect 7452 2628 7470 2646
rect 7452 2646 7470 2664
rect 7452 2664 7470 2682
rect 7452 2682 7470 2700
rect 7452 2700 7470 2718
rect 7452 2718 7470 2736
rect 7452 2736 7470 2754
rect 7452 2754 7470 2772
rect 7452 2772 7470 2790
rect 7452 2790 7470 2808
rect 7452 2808 7470 2826
rect 7452 2826 7470 2844
rect 7452 2844 7470 2862
rect 7452 2862 7470 2880
rect 7452 2880 7470 2898
rect 7452 2898 7470 2916
rect 7452 2916 7470 2934
rect 7452 2934 7470 2952
rect 7452 2952 7470 2970
rect 7452 2970 7470 2988
rect 7452 2988 7470 3006
rect 7452 3006 7470 3024
rect 7452 3024 7470 3042
rect 7452 3042 7470 3060
rect 7452 3060 7470 3078
rect 7452 3078 7470 3096
rect 7452 3096 7470 3114
rect 7452 3114 7470 3132
rect 7452 3132 7470 3150
rect 7452 3150 7470 3168
rect 7452 3168 7470 3186
rect 7452 3186 7470 3204
rect 7452 3204 7470 3222
rect 7452 4590 7470 4608
rect 7452 4608 7470 4626
rect 7452 4626 7470 4644
rect 7452 4644 7470 4662
rect 7452 4662 7470 4680
rect 7452 4680 7470 4698
rect 7452 4698 7470 4716
rect 7452 4716 7470 4734
rect 7452 4734 7470 4752
rect 7452 4752 7470 4770
rect 7452 4770 7470 4788
rect 7452 4788 7470 4806
rect 7452 4806 7470 4824
rect 7452 4824 7470 4842
rect 7452 4842 7470 4860
rect 7452 4860 7470 4878
rect 7452 4878 7470 4896
rect 7452 4896 7470 4914
rect 7452 4914 7470 4932
rect 7452 4932 7470 4950
rect 7452 4950 7470 4968
rect 7452 4968 7470 4986
rect 7452 4986 7470 5004
rect 7452 5004 7470 5022
rect 7452 5022 7470 5040
rect 7452 5040 7470 5058
rect 7452 5058 7470 5076
rect 7452 5076 7470 5094
rect 7452 5094 7470 5112
rect 7452 5112 7470 5130
rect 7452 5130 7470 5148
rect 7452 5148 7470 5166
rect 7452 5166 7470 5184
rect 7452 5184 7470 5202
rect 7452 5202 7470 5220
rect 7452 5220 7470 5238
rect 7452 5238 7470 5256
rect 7452 5256 7470 5274
rect 7452 5274 7470 5292
rect 7452 5292 7470 5310
rect 7452 5310 7470 5328
rect 7452 5328 7470 5346
rect 7452 5346 7470 5364
rect 7452 5364 7470 5382
rect 7452 5382 7470 5400
rect 7452 5400 7470 5418
rect 7452 5418 7470 5436
rect 7452 5436 7470 5454
rect 7452 5454 7470 5472
rect 7452 5472 7470 5490
rect 7452 5490 7470 5508
rect 7452 5508 7470 5526
rect 7452 5526 7470 5544
rect 7452 5544 7470 5562
rect 7452 5562 7470 5580
rect 7452 5580 7470 5598
rect 7452 5598 7470 5616
rect 7452 5616 7470 5634
rect 7452 5634 7470 5652
rect 7452 5652 7470 5670
rect 7452 5670 7470 5688
rect 7452 5688 7470 5706
rect 7452 5706 7470 5724
rect 7452 5724 7470 5742
rect 7452 5742 7470 5760
rect 7452 5760 7470 5778
rect 7452 5778 7470 5796
rect 7452 5796 7470 5814
rect 7452 5814 7470 5832
rect 7452 5832 7470 5850
rect 7452 5850 7470 5868
rect 7452 5868 7470 5886
rect 7452 5886 7470 5904
rect 7452 5904 7470 5922
rect 7452 5922 7470 5940
rect 7452 5940 7470 5958
rect 7452 5958 7470 5976
rect 7452 5976 7470 5994
rect 7452 5994 7470 6012
rect 7452 6012 7470 6030
rect 7452 6030 7470 6048
rect 7452 6048 7470 6066
rect 7452 6066 7470 6084
rect 7452 6084 7470 6102
rect 7452 6102 7470 6120
rect 7452 6120 7470 6138
rect 7452 6138 7470 6156
rect 7452 6156 7470 6174
rect 7452 6174 7470 6192
rect 7452 6192 7470 6210
rect 7452 6210 7470 6228
rect 7452 6228 7470 6246
rect 7452 6246 7470 6264
rect 7452 6264 7470 6282
rect 7452 6282 7470 6300
rect 7452 6300 7470 6318
rect 7452 6318 7470 6336
rect 7452 6336 7470 6354
rect 7452 6354 7470 6372
rect 7452 6372 7470 6390
rect 7452 6390 7470 6408
rect 7452 6408 7470 6426
rect 7452 6426 7470 6444
rect 7452 6444 7470 6462
rect 7452 6462 7470 6480
rect 7452 6480 7470 6498
rect 7452 6498 7470 6516
rect 7452 6516 7470 6534
rect 7452 6534 7470 6552
rect 7452 6552 7470 6570
rect 7452 6570 7470 6588
rect 7452 6588 7470 6606
rect 7452 6606 7470 6624
rect 7470 2070 7488 2088
rect 7470 2088 7488 2106
rect 7470 2106 7488 2124
rect 7470 2124 7488 2142
rect 7470 2142 7488 2160
rect 7470 2160 7488 2178
rect 7470 2178 7488 2196
rect 7470 2196 7488 2214
rect 7470 2214 7488 2232
rect 7470 2232 7488 2250
rect 7470 2250 7488 2268
rect 7470 2268 7488 2286
rect 7470 2286 7488 2304
rect 7470 2304 7488 2322
rect 7470 2322 7488 2340
rect 7470 2340 7488 2358
rect 7470 2358 7488 2376
rect 7470 2376 7488 2394
rect 7470 2394 7488 2412
rect 7470 2412 7488 2430
rect 7470 2430 7488 2448
rect 7470 2448 7488 2466
rect 7470 2466 7488 2484
rect 7470 2484 7488 2502
rect 7470 2502 7488 2520
rect 7470 2520 7488 2538
rect 7470 2538 7488 2556
rect 7470 2556 7488 2574
rect 7470 2574 7488 2592
rect 7470 2592 7488 2610
rect 7470 2610 7488 2628
rect 7470 2628 7488 2646
rect 7470 2646 7488 2664
rect 7470 2664 7488 2682
rect 7470 2682 7488 2700
rect 7470 2700 7488 2718
rect 7470 2718 7488 2736
rect 7470 2736 7488 2754
rect 7470 2754 7488 2772
rect 7470 2772 7488 2790
rect 7470 2790 7488 2808
rect 7470 2808 7488 2826
rect 7470 2826 7488 2844
rect 7470 2844 7488 2862
rect 7470 2862 7488 2880
rect 7470 2880 7488 2898
rect 7470 2898 7488 2916
rect 7470 2916 7488 2934
rect 7470 2934 7488 2952
rect 7470 2952 7488 2970
rect 7470 2970 7488 2988
rect 7470 2988 7488 3006
rect 7470 3006 7488 3024
rect 7470 3024 7488 3042
rect 7470 3042 7488 3060
rect 7470 3060 7488 3078
rect 7470 3078 7488 3096
rect 7470 3096 7488 3114
rect 7470 3114 7488 3132
rect 7470 3132 7488 3150
rect 7470 3150 7488 3168
rect 7470 3168 7488 3186
rect 7470 3186 7488 3204
rect 7470 3204 7488 3222
rect 7470 4608 7488 4626
rect 7470 4626 7488 4644
rect 7470 4644 7488 4662
rect 7470 4662 7488 4680
rect 7470 4680 7488 4698
rect 7470 4698 7488 4716
rect 7470 4716 7488 4734
rect 7470 4734 7488 4752
rect 7470 4752 7488 4770
rect 7470 4770 7488 4788
rect 7470 4788 7488 4806
rect 7470 4806 7488 4824
rect 7470 4824 7488 4842
rect 7470 4842 7488 4860
rect 7470 4860 7488 4878
rect 7470 4878 7488 4896
rect 7470 4896 7488 4914
rect 7470 4914 7488 4932
rect 7470 4932 7488 4950
rect 7470 4950 7488 4968
rect 7470 4968 7488 4986
rect 7470 4986 7488 5004
rect 7470 5004 7488 5022
rect 7470 5022 7488 5040
rect 7470 5040 7488 5058
rect 7470 5058 7488 5076
rect 7470 5076 7488 5094
rect 7470 5094 7488 5112
rect 7470 5112 7488 5130
rect 7470 5130 7488 5148
rect 7470 5148 7488 5166
rect 7470 5166 7488 5184
rect 7470 5184 7488 5202
rect 7470 5202 7488 5220
rect 7470 5220 7488 5238
rect 7470 5238 7488 5256
rect 7470 5256 7488 5274
rect 7470 5274 7488 5292
rect 7470 5292 7488 5310
rect 7470 5310 7488 5328
rect 7470 5328 7488 5346
rect 7470 5346 7488 5364
rect 7470 5364 7488 5382
rect 7470 5382 7488 5400
rect 7470 5400 7488 5418
rect 7470 5418 7488 5436
rect 7470 5436 7488 5454
rect 7470 5454 7488 5472
rect 7470 5472 7488 5490
rect 7470 5490 7488 5508
rect 7470 5508 7488 5526
rect 7470 5526 7488 5544
rect 7470 5544 7488 5562
rect 7470 5562 7488 5580
rect 7470 5580 7488 5598
rect 7470 5598 7488 5616
rect 7470 5616 7488 5634
rect 7470 5634 7488 5652
rect 7470 5652 7488 5670
rect 7470 5670 7488 5688
rect 7470 5688 7488 5706
rect 7470 5706 7488 5724
rect 7470 5724 7488 5742
rect 7470 5742 7488 5760
rect 7470 5760 7488 5778
rect 7470 5778 7488 5796
rect 7470 5796 7488 5814
rect 7470 5814 7488 5832
rect 7470 5832 7488 5850
rect 7470 5850 7488 5868
rect 7470 5868 7488 5886
rect 7470 5886 7488 5904
rect 7470 5904 7488 5922
rect 7470 5922 7488 5940
rect 7470 5940 7488 5958
rect 7470 5958 7488 5976
rect 7470 5976 7488 5994
rect 7470 5994 7488 6012
rect 7470 6012 7488 6030
rect 7470 6030 7488 6048
rect 7470 6048 7488 6066
rect 7470 6066 7488 6084
rect 7470 6084 7488 6102
rect 7470 6102 7488 6120
rect 7470 6120 7488 6138
rect 7470 6138 7488 6156
rect 7470 6156 7488 6174
rect 7470 6174 7488 6192
rect 7470 6192 7488 6210
rect 7470 6210 7488 6228
rect 7470 6228 7488 6246
rect 7470 6246 7488 6264
rect 7470 6264 7488 6282
rect 7470 6282 7488 6300
rect 7470 6300 7488 6318
rect 7470 6318 7488 6336
rect 7470 6336 7488 6354
rect 7470 6354 7488 6372
rect 7470 6372 7488 6390
rect 7470 6390 7488 6408
rect 7470 6408 7488 6426
rect 7470 6426 7488 6444
rect 7470 6444 7488 6462
rect 7470 6462 7488 6480
rect 7470 6480 7488 6498
rect 7470 6498 7488 6516
rect 7470 6516 7488 6534
rect 7470 6534 7488 6552
rect 7470 6552 7488 6570
rect 7470 6570 7488 6588
rect 7470 6588 7488 6606
rect 7470 6606 7488 6624
rect 7470 6624 7488 6642
rect 7488 2088 7506 2106
rect 7488 2106 7506 2124
rect 7488 2124 7506 2142
rect 7488 2142 7506 2160
rect 7488 2160 7506 2178
rect 7488 2178 7506 2196
rect 7488 2196 7506 2214
rect 7488 2214 7506 2232
rect 7488 2232 7506 2250
rect 7488 2250 7506 2268
rect 7488 2268 7506 2286
rect 7488 2286 7506 2304
rect 7488 2304 7506 2322
rect 7488 2322 7506 2340
rect 7488 2340 7506 2358
rect 7488 2358 7506 2376
rect 7488 2376 7506 2394
rect 7488 2394 7506 2412
rect 7488 2412 7506 2430
rect 7488 2430 7506 2448
rect 7488 2448 7506 2466
rect 7488 2466 7506 2484
rect 7488 2484 7506 2502
rect 7488 2502 7506 2520
rect 7488 2520 7506 2538
rect 7488 2538 7506 2556
rect 7488 2556 7506 2574
rect 7488 2574 7506 2592
rect 7488 2592 7506 2610
rect 7488 2610 7506 2628
rect 7488 2628 7506 2646
rect 7488 2646 7506 2664
rect 7488 2664 7506 2682
rect 7488 2682 7506 2700
rect 7488 2700 7506 2718
rect 7488 2718 7506 2736
rect 7488 2736 7506 2754
rect 7488 2754 7506 2772
rect 7488 2772 7506 2790
rect 7488 2790 7506 2808
rect 7488 2808 7506 2826
rect 7488 2826 7506 2844
rect 7488 2844 7506 2862
rect 7488 2862 7506 2880
rect 7488 2880 7506 2898
rect 7488 2898 7506 2916
rect 7488 2916 7506 2934
rect 7488 2934 7506 2952
rect 7488 2952 7506 2970
rect 7488 2970 7506 2988
rect 7488 2988 7506 3006
rect 7488 3006 7506 3024
rect 7488 3024 7506 3042
rect 7488 3042 7506 3060
rect 7488 3060 7506 3078
rect 7488 3078 7506 3096
rect 7488 3096 7506 3114
rect 7488 3114 7506 3132
rect 7488 3132 7506 3150
rect 7488 3150 7506 3168
rect 7488 3168 7506 3186
rect 7488 3186 7506 3204
rect 7488 3204 7506 3222
rect 7488 4626 7506 4644
rect 7488 4644 7506 4662
rect 7488 4662 7506 4680
rect 7488 4680 7506 4698
rect 7488 4698 7506 4716
rect 7488 4716 7506 4734
rect 7488 4734 7506 4752
rect 7488 4752 7506 4770
rect 7488 4770 7506 4788
rect 7488 4788 7506 4806
rect 7488 4806 7506 4824
rect 7488 4824 7506 4842
rect 7488 4842 7506 4860
rect 7488 4860 7506 4878
rect 7488 4878 7506 4896
rect 7488 4896 7506 4914
rect 7488 4914 7506 4932
rect 7488 4932 7506 4950
rect 7488 4950 7506 4968
rect 7488 4968 7506 4986
rect 7488 4986 7506 5004
rect 7488 5004 7506 5022
rect 7488 5022 7506 5040
rect 7488 5040 7506 5058
rect 7488 5058 7506 5076
rect 7488 5076 7506 5094
rect 7488 5094 7506 5112
rect 7488 5112 7506 5130
rect 7488 5130 7506 5148
rect 7488 5148 7506 5166
rect 7488 5166 7506 5184
rect 7488 5184 7506 5202
rect 7488 5202 7506 5220
rect 7488 5220 7506 5238
rect 7488 5238 7506 5256
rect 7488 5256 7506 5274
rect 7488 5274 7506 5292
rect 7488 5292 7506 5310
rect 7488 5310 7506 5328
rect 7488 5328 7506 5346
rect 7488 5346 7506 5364
rect 7488 5364 7506 5382
rect 7488 5382 7506 5400
rect 7488 5400 7506 5418
rect 7488 5418 7506 5436
rect 7488 5436 7506 5454
rect 7488 5454 7506 5472
rect 7488 5472 7506 5490
rect 7488 5490 7506 5508
rect 7488 5508 7506 5526
rect 7488 5526 7506 5544
rect 7488 5544 7506 5562
rect 7488 5562 7506 5580
rect 7488 5580 7506 5598
rect 7488 5598 7506 5616
rect 7488 5616 7506 5634
rect 7488 5634 7506 5652
rect 7488 5652 7506 5670
rect 7488 5670 7506 5688
rect 7488 5688 7506 5706
rect 7488 5706 7506 5724
rect 7488 5724 7506 5742
rect 7488 5742 7506 5760
rect 7488 5760 7506 5778
rect 7488 5778 7506 5796
rect 7488 5796 7506 5814
rect 7488 5814 7506 5832
rect 7488 5832 7506 5850
rect 7488 5850 7506 5868
rect 7488 5868 7506 5886
rect 7488 5886 7506 5904
rect 7488 5904 7506 5922
rect 7488 5922 7506 5940
rect 7488 5940 7506 5958
rect 7488 5958 7506 5976
rect 7488 5976 7506 5994
rect 7488 5994 7506 6012
rect 7488 6012 7506 6030
rect 7488 6030 7506 6048
rect 7488 6048 7506 6066
rect 7488 6066 7506 6084
rect 7488 6084 7506 6102
rect 7488 6102 7506 6120
rect 7488 6120 7506 6138
rect 7488 6138 7506 6156
rect 7488 6156 7506 6174
rect 7488 6174 7506 6192
rect 7488 6192 7506 6210
rect 7488 6210 7506 6228
rect 7488 6228 7506 6246
rect 7488 6246 7506 6264
rect 7488 6264 7506 6282
rect 7488 6282 7506 6300
rect 7488 6300 7506 6318
rect 7488 6318 7506 6336
rect 7488 6336 7506 6354
rect 7488 6354 7506 6372
rect 7488 6372 7506 6390
rect 7488 6390 7506 6408
rect 7488 6408 7506 6426
rect 7488 6426 7506 6444
rect 7488 6444 7506 6462
rect 7488 6462 7506 6480
rect 7488 6480 7506 6498
rect 7488 6498 7506 6516
rect 7488 6516 7506 6534
rect 7488 6534 7506 6552
rect 7488 6552 7506 6570
rect 7488 6570 7506 6588
rect 7488 6588 7506 6606
rect 7488 6606 7506 6624
rect 7488 6624 7506 6642
rect 7506 2088 7524 2106
rect 7506 2106 7524 2124
rect 7506 2124 7524 2142
rect 7506 2142 7524 2160
rect 7506 2160 7524 2178
rect 7506 2178 7524 2196
rect 7506 2196 7524 2214
rect 7506 2214 7524 2232
rect 7506 2232 7524 2250
rect 7506 2250 7524 2268
rect 7506 2268 7524 2286
rect 7506 2286 7524 2304
rect 7506 2304 7524 2322
rect 7506 2322 7524 2340
rect 7506 2340 7524 2358
rect 7506 2358 7524 2376
rect 7506 2376 7524 2394
rect 7506 2394 7524 2412
rect 7506 2412 7524 2430
rect 7506 2430 7524 2448
rect 7506 2448 7524 2466
rect 7506 2466 7524 2484
rect 7506 2484 7524 2502
rect 7506 2502 7524 2520
rect 7506 2520 7524 2538
rect 7506 2538 7524 2556
rect 7506 2556 7524 2574
rect 7506 2574 7524 2592
rect 7506 2592 7524 2610
rect 7506 2610 7524 2628
rect 7506 2628 7524 2646
rect 7506 2646 7524 2664
rect 7506 2664 7524 2682
rect 7506 2682 7524 2700
rect 7506 2700 7524 2718
rect 7506 2718 7524 2736
rect 7506 2736 7524 2754
rect 7506 2754 7524 2772
rect 7506 2772 7524 2790
rect 7506 2790 7524 2808
rect 7506 2808 7524 2826
rect 7506 2826 7524 2844
rect 7506 2844 7524 2862
rect 7506 2862 7524 2880
rect 7506 2880 7524 2898
rect 7506 2898 7524 2916
rect 7506 2916 7524 2934
rect 7506 2934 7524 2952
rect 7506 2952 7524 2970
rect 7506 2970 7524 2988
rect 7506 2988 7524 3006
rect 7506 3006 7524 3024
rect 7506 3024 7524 3042
rect 7506 3042 7524 3060
rect 7506 3060 7524 3078
rect 7506 3078 7524 3096
rect 7506 3096 7524 3114
rect 7506 3114 7524 3132
rect 7506 3132 7524 3150
rect 7506 3150 7524 3168
rect 7506 3168 7524 3186
rect 7506 3186 7524 3204
rect 7506 3204 7524 3222
rect 7506 3222 7524 3240
rect 7506 4644 7524 4662
rect 7506 4662 7524 4680
rect 7506 4680 7524 4698
rect 7506 4698 7524 4716
rect 7506 4716 7524 4734
rect 7506 4734 7524 4752
rect 7506 4752 7524 4770
rect 7506 4770 7524 4788
rect 7506 4788 7524 4806
rect 7506 4806 7524 4824
rect 7506 4824 7524 4842
rect 7506 4842 7524 4860
rect 7506 4860 7524 4878
rect 7506 4878 7524 4896
rect 7506 4896 7524 4914
rect 7506 4914 7524 4932
rect 7506 4932 7524 4950
rect 7506 4950 7524 4968
rect 7506 4968 7524 4986
rect 7506 4986 7524 5004
rect 7506 5004 7524 5022
rect 7506 5022 7524 5040
rect 7506 5040 7524 5058
rect 7506 5058 7524 5076
rect 7506 5076 7524 5094
rect 7506 5094 7524 5112
rect 7506 5112 7524 5130
rect 7506 5130 7524 5148
rect 7506 5148 7524 5166
rect 7506 5166 7524 5184
rect 7506 5184 7524 5202
rect 7506 5202 7524 5220
rect 7506 5220 7524 5238
rect 7506 5238 7524 5256
rect 7506 5256 7524 5274
rect 7506 5274 7524 5292
rect 7506 5292 7524 5310
rect 7506 5310 7524 5328
rect 7506 5328 7524 5346
rect 7506 5346 7524 5364
rect 7506 5364 7524 5382
rect 7506 5382 7524 5400
rect 7506 5400 7524 5418
rect 7506 5418 7524 5436
rect 7506 5436 7524 5454
rect 7506 5454 7524 5472
rect 7506 5472 7524 5490
rect 7506 5490 7524 5508
rect 7506 5508 7524 5526
rect 7506 5526 7524 5544
rect 7506 5544 7524 5562
rect 7506 5562 7524 5580
rect 7506 5580 7524 5598
rect 7506 5598 7524 5616
rect 7506 5616 7524 5634
rect 7506 5634 7524 5652
rect 7506 5652 7524 5670
rect 7506 5670 7524 5688
rect 7506 5688 7524 5706
rect 7506 5706 7524 5724
rect 7506 5724 7524 5742
rect 7506 5742 7524 5760
rect 7506 5760 7524 5778
rect 7506 5778 7524 5796
rect 7506 5796 7524 5814
rect 7506 5814 7524 5832
rect 7506 5832 7524 5850
rect 7506 5850 7524 5868
rect 7506 5868 7524 5886
rect 7506 5886 7524 5904
rect 7506 5904 7524 5922
rect 7506 5922 7524 5940
rect 7506 5940 7524 5958
rect 7506 5958 7524 5976
rect 7506 5976 7524 5994
rect 7506 5994 7524 6012
rect 7506 6012 7524 6030
rect 7506 6030 7524 6048
rect 7506 6048 7524 6066
rect 7506 6066 7524 6084
rect 7506 6084 7524 6102
rect 7506 6102 7524 6120
rect 7506 6120 7524 6138
rect 7506 6138 7524 6156
rect 7506 6156 7524 6174
rect 7506 6174 7524 6192
rect 7506 6192 7524 6210
rect 7506 6210 7524 6228
rect 7506 6228 7524 6246
rect 7506 6246 7524 6264
rect 7506 6264 7524 6282
rect 7506 6282 7524 6300
rect 7506 6300 7524 6318
rect 7506 6318 7524 6336
rect 7506 6336 7524 6354
rect 7506 6354 7524 6372
rect 7506 6372 7524 6390
rect 7506 6390 7524 6408
rect 7506 6408 7524 6426
rect 7506 6426 7524 6444
rect 7506 6444 7524 6462
rect 7506 6462 7524 6480
rect 7506 6480 7524 6498
rect 7506 6498 7524 6516
rect 7506 6516 7524 6534
rect 7506 6534 7524 6552
rect 7506 6552 7524 6570
rect 7506 6570 7524 6588
rect 7506 6588 7524 6606
rect 7506 6606 7524 6624
rect 7506 6624 7524 6642
rect 7506 6642 7524 6660
rect 7524 2106 7542 2124
rect 7524 2124 7542 2142
rect 7524 2142 7542 2160
rect 7524 2160 7542 2178
rect 7524 2178 7542 2196
rect 7524 2196 7542 2214
rect 7524 2214 7542 2232
rect 7524 2232 7542 2250
rect 7524 2250 7542 2268
rect 7524 2268 7542 2286
rect 7524 2286 7542 2304
rect 7524 2304 7542 2322
rect 7524 2322 7542 2340
rect 7524 2340 7542 2358
rect 7524 2358 7542 2376
rect 7524 2376 7542 2394
rect 7524 2394 7542 2412
rect 7524 2412 7542 2430
rect 7524 2430 7542 2448
rect 7524 2448 7542 2466
rect 7524 2466 7542 2484
rect 7524 2484 7542 2502
rect 7524 2502 7542 2520
rect 7524 2520 7542 2538
rect 7524 2538 7542 2556
rect 7524 2556 7542 2574
rect 7524 2574 7542 2592
rect 7524 2592 7542 2610
rect 7524 2610 7542 2628
rect 7524 2628 7542 2646
rect 7524 2646 7542 2664
rect 7524 2664 7542 2682
rect 7524 2682 7542 2700
rect 7524 2700 7542 2718
rect 7524 2718 7542 2736
rect 7524 2736 7542 2754
rect 7524 2754 7542 2772
rect 7524 2772 7542 2790
rect 7524 2790 7542 2808
rect 7524 2808 7542 2826
rect 7524 2826 7542 2844
rect 7524 2844 7542 2862
rect 7524 2862 7542 2880
rect 7524 2880 7542 2898
rect 7524 2898 7542 2916
rect 7524 2916 7542 2934
rect 7524 2934 7542 2952
rect 7524 2952 7542 2970
rect 7524 2970 7542 2988
rect 7524 2988 7542 3006
rect 7524 3006 7542 3024
rect 7524 3024 7542 3042
rect 7524 3042 7542 3060
rect 7524 3060 7542 3078
rect 7524 3078 7542 3096
rect 7524 3096 7542 3114
rect 7524 3114 7542 3132
rect 7524 3132 7542 3150
rect 7524 3150 7542 3168
rect 7524 3168 7542 3186
rect 7524 3186 7542 3204
rect 7524 3204 7542 3222
rect 7524 3222 7542 3240
rect 7524 4680 7542 4698
rect 7524 4698 7542 4716
rect 7524 4716 7542 4734
rect 7524 4734 7542 4752
rect 7524 4752 7542 4770
rect 7524 4770 7542 4788
rect 7524 4788 7542 4806
rect 7524 4806 7542 4824
rect 7524 4824 7542 4842
rect 7524 4842 7542 4860
rect 7524 4860 7542 4878
rect 7524 4878 7542 4896
rect 7524 4896 7542 4914
rect 7524 4914 7542 4932
rect 7524 4932 7542 4950
rect 7524 4950 7542 4968
rect 7524 4968 7542 4986
rect 7524 4986 7542 5004
rect 7524 5004 7542 5022
rect 7524 5022 7542 5040
rect 7524 5040 7542 5058
rect 7524 5058 7542 5076
rect 7524 5076 7542 5094
rect 7524 5094 7542 5112
rect 7524 5112 7542 5130
rect 7524 5130 7542 5148
rect 7524 5148 7542 5166
rect 7524 5166 7542 5184
rect 7524 5184 7542 5202
rect 7524 5202 7542 5220
rect 7524 5220 7542 5238
rect 7524 5238 7542 5256
rect 7524 5256 7542 5274
rect 7524 5274 7542 5292
rect 7524 5292 7542 5310
rect 7524 5310 7542 5328
rect 7524 5328 7542 5346
rect 7524 5346 7542 5364
rect 7524 5364 7542 5382
rect 7524 5382 7542 5400
rect 7524 5400 7542 5418
rect 7524 5418 7542 5436
rect 7524 5436 7542 5454
rect 7524 5454 7542 5472
rect 7524 5472 7542 5490
rect 7524 5490 7542 5508
rect 7524 5508 7542 5526
rect 7524 5526 7542 5544
rect 7524 5544 7542 5562
rect 7524 5562 7542 5580
rect 7524 5580 7542 5598
rect 7524 5598 7542 5616
rect 7524 5616 7542 5634
rect 7524 5634 7542 5652
rect 7524 5652 7542 5670
rect 7524 5670 7542 5688
rect 7524 5688 7542 5706
rect 7524 5706 7542 5724
rect 7524 5724 7542 5742
rect 7524 5742 7542 5760
rect 7524 5760 7542 5778
rect 7524 5778 7542 5796
rect 7524 5796 7542 5814
rect 7524 5814 7542 5832
rect 7524 5832 7542 5850
rect 7524 5850 7542 5868
rect 7524 5868 7542 5886
rect 7524 5886 7542 5904
rect 7524 5904 7542 5922
rect 7524 5922 7542 5940
rect 7524 5940 7542 5958
rect 7524 5958 7542 5976
rect 7524 5976 7542 5994
rect 7524 5994 7542 6012
rect 7524 6012 7542 6030
rect 7524 6030 7542 6048
rect 7524 6048 7542 6066
rect 7524 6066 7542 6084
rect 7524 6084 7542 6102
rect 7524 6102 7542 6120
rect 7524 6120 7542 6138
rect 7524 6138 7542 6156
rect 7524 6156 7542 6174
rect 7524 6174 7542 6192
rect 7524 6192 7542 6210
rect 7524 6210 7542 6228
rect 7524 6228 7542 6246
rect 7524 6246 7542 6264
rect 7524 6264 7542 6282
rect 7524 6282 7542 6300
rect 7524 6300 7542 6318
rect 7524 6318 7542 6336
rect 7524 6336 7542 6354
rect 7524 6354 7542 6372
rect 7524 6372 7542 6390
rect 7524 6390 7542 6408
rect 7524 6408 7542 6426
rect 7524 6426 7542 6444
rect 7524 6444 7542 6462
rect 7524 6462 7542 6480
rect 7524 6480 7542 6498
rect 7524 6498 7542 6516
rect 7524 6516 7542 6534
rect 7524 6534 7542 6552
rect 7524 6552 7542 6570
rect 7524 6570 7542 6588
rect 7524 6588 7542 6606
rect 7524 6606 7542 6624
rect 7524 6624 7542 6642
rect 7524 6642 7542 6660
rect 7524 6660 7542 6678
rect 7542 2106 7560 2124
rect 7542 2124 7560 2142
rect 7542 2142 7560 2160
rect 7542 2160 7560 2178
rect 7542 2178 7560 2196
rect 7542 2196 7560 2214
rect 7542 2214 7560 2232
rect 7542 2232 7560 2250
rect 7542 2250 7560 2268
rect 7542 2268 7560 2286
rect 7542 2286 7560 2304
rect 7542 2304 7560 2322
rect 7542 2322 7560 2340
rect 7542 2340 7560 2358
rect 7542 2358 7560 2376
rect 7542 2376 7560 2394
rect 7542 2394 7560 2412
rect 7542 2412 7560 2430
rect 7542 2430 7560 2448
rect 7542 2448 7560 2466
rect 7542 2466 7560 2484
rect 7542 2484 7560 2502
rect 7542 2502 7560 2520
rect 7542 2520 7560 2538
rect 7542 2538 7560 2556
rect 7542 2556 7560 2574
rect 7542 2574 7560 2592
rect 7542 2592 7560 2610
rect 7542 2610 7560 2628
rect 7542 2628 7560 2646
rect 7542 2646 7560 2664
rect 7542 2664 7560 2682
rect 7542 2682 7560 2700
rect 7542 2700 7560 2718
rect 7542 2718 7560 2736
rect 7542 2736 7560 2754
rect 7542 2754 7560 2772
rect 7542 2772 7560 2790
rect 7542 2790 7560 2808
rect 7542 2808 7560 2826
rect 7542 2826 7560 2844
rect 7542 2844 7560 2862
rect 7542 2862 7560 2880
rect 7542 2880 7560 2898
rect 7542 2898 7560 2916
rect 7542 2916 7560 2934
rect 7542 2934 7560 2952
rect 7542 2952 7560 2970
rect 7542 2970 7560 2988
rect 7542 2988 7560 3006
rect 7542 3006 7560 3024
rect 7542 3024 7560 3042
rect 7542 3042 7560 3060
rect 7542 3060 7560 3078
rect 7542 3078 7560 3096
rect 7542 3096 7560 3114
rect 7542 3114 7560 3132
rect 7542 3132 7560 3150
rect 7542 3150 7560 3168
rect 7542 3168 7560 3186
rect 7542 3186 7560 3204
rect 7542 3204 7560 3222
rect 7542 3222 7560 3240
rect 7542 4698 7560 4716
rect 7542 4716 7560 4734
rect 7542 4734 7560 4752
rect 7542 4752 7560 4770
rect 7542 4770 7560 4788
rect 7542 4788 7560 4806
rect 7542 4806 7560 4824
rect 7542 4824 7560 4842
rect 7542 4842 7560 4860
rect 7542 4860 7560 4878
rect 7542 4878 7560 4896
rect 7542 4896 7560 4914
rect 7542 4914 7560 4932
rect 7542 4932 7560 4950
rect 7542 4950 7560 4968
rect 7542 4968 7560 4986
rect 7542 4986 7560 5004
rect 7542 5004 7560 5022
rect 7542 5022 7560 5040
rect 7542 5040 7560 5058
rect 7542 5058 7560 5076
rect 7542 5076 7560 5094
rect 7542 5094 7560 5112
rect 7542 5112 7560 5130
rect 7542 5130 7560 5148
rect 7542 5148 7560 5166
rect 7542 5166 7560 5184
rect 7542 5184 7560 5202
rect 7542 5202 7560 5220
rect 7542 5220 7560 5238
rect 7542 5238 7560 5256
rect 7542 5256 7560 5274
rect 7542 5274 7560 5292
rect 7542 5292 7560 5310
rect 7542 5310 7560 5328
rect 7542 5328 7560 5346
rect 7542 5346 7560 5364
rect 7542 5364 7560 5382
rect 7542 5382 7560 5400
rect 7542 5400 7560 5418
rect 7542 5418 7560 5436
rect 7542 5436 7560 5454
rect 7542 5454 7560 5472
rect 7542 5472 7560 5490
rect 7542 5490 7560 5508
rect 7542 5508 7560 5526
rect 7542 5526 7560 5544
rect 7542 5544 7560 5562
rect 7542 5562 7560 5580
rect 7542 5580 7560 5598
rect 7542 5598 7560 5616
rect 7542 5616 7560 5634
rect 7542 5634 7560 5652
rect 7542 5652 7560 5670
rect 7542 5670 7560 5688
rect 7542 5688 7560 5706
rect 7542 5706 7560 5724
rect 7542 5724 7560 5742
rect 7542 5742 7560 5760
rect 7542 5760 7560 5778
rect 7542 5778 7560 5796
rect 7542 5796 7560 5814
rect 7542 5814 7560 5832
rect 7542 5832 7560 5850
rect 7542 5850 7560 5868
rect 7542 5868 7560 5886
rect 7542 5886 7560 5904
rect 7542 5904 7560 5922
rect 7542 5922 7560 5940
rect 7542 5940 7560 5958
rect 7542 5958 7560 5976
rect 7542 5976 7560 5994
rect 7542 5994 7560 6012
rect 7542 6012 7560 6030
rect 7542 6030 7560 6048
rect 7542 6048 7560 6066
rect 7542 6066 7560 6084
rect 7542 6084 7560 6102
rect 7542 6102 7560 6120
rect 7542 6120 7560 6138
rect 7542 6138 7560 6156
rect 7542 6156 7560 6174
rect 7542 6174 7560 6192
rect 7542 6192 7560 6210
rect 7542 6210 7560 6228
rect 7542 6228 7560 6246
rect 7542 6246 7560 6264
rect 7542 6264 7560 6282
rect 7542 6282 7560 6300
rect 7542 6300 7560 6318
rect 7542 6318 7560 6336
rect 7542 6336 7560 6354
rect 7542 6354 7560 6372
rect 7542 6372 7560 6390
rect 7542 6390 7560 6408
rect 7542 6408 7560 6426
rect 7542 6426 7560 6444
rect 7542 6444 7560 6462
rect 7542 6462 7560 6480
rect 7542 6480 7560 6498
rect 7542 6498 7560 6516
rect 7542 6516 7560 6534
rect 7542 6534 7560 6552
rect 7542 6552 7560 6570
rect 7542 6570 7560 6588
rect 7542 6588 7560 6606
rect 7542 6606 7560 6624
rect 7542 6624 7560 6642
rect 7542 6642 7560 6660
rect 7542 6660 7560 6678
rect 7542 6678 7560 6696
rect 7560 2124 7578 2142
rect 7560 2142 7578 2160
rect 7560 2160 7578 2178
rect 7560 2178 7578 2196
rect 7560 2196 7578 2214
rect 7560 2214 7578 2232
rect 7560 2232 7578 2250
rect 7560 2250 7578 2268
rect 7560 2268 7578 2286
rect 7560 2286 7578 2304
rect 7560 2304 7578 2322
rect 7560 2322 7578 2340
rect 7560 2340 7578 2358
rect 7560 2358 7578 2376
rect 7560 2376 7578 2394
rect 7560 2394 7578 2412
rect 7560 2412 7578 2430
rect 7560 2430 7578 2448
rect 7560 2448 7578 2466
rect 7560 2466 7578 2484
rect 7560 2484 7578 2502
rect 7560 2502 7578 2520
rect 7560 2520 7578 2538
rect 7560 2538 7578 2556
rect 7560 2556 7578 2574
rect 7560 2574 7578 2592
rect 7560 2592 7578 2610
rect 7560 2610 7578 2628
rect 7560 2628 7578 2646
rect 7560 2646 7578 2664
rect 7560 2664 7578 2682
rect 7560 2682 7578 2700
rect 7560 2700 7578 2718
rect 7560 2718 7578 2736
rect 7560 2736 7578 2754
rect 7560 2754 7578 2772
rect 7560 2772 7578 2790
rect 7560 2790 7578 2808
rect 7560 2808 7578 2826
rect 7560 2826 7578 2844
rect 7560 2844 7578 2862
rect 7560 2862 7578 2880
rect 7560 2880 7578 2898
rect 7560 2898 7578 2916
rect 7560 2916 7578 2934
rect 7560 2934 7578 2952
rect 7560 2952 7578 2970
rect 7560 2970 7578 2988
rect 7560 2988 7578 3006
rect 7560 3006 7578 3024
rect 7560 3024 7578 3042
rect 7560 3042 7578 3060
rect 7560 3060 7578 3078
rect 7560 3078 7578 3096
rect 7560 3096 7578 3114
rect 7560 3114 7578 3132
rect 7560 3132 7578 3150
rect 7560 3150 7578 3168
rect 7560 3168 7578 3186
rect 7560 3186 7578 3204
rect 7560 3204 7578 3222
rect 7560 3222 7578 3240
rect 7560 3240 7578 3258
rect 7560 4716 7578 4734
rect 7560 4734 7578 4752
rect 7560 4752 7578 4770
rect 7560 4770 7578 4788
rect 7560 4788 7578 4806
rect 7560 4806 7578 4824
rect 7560 4824 7578 4842
rect 7560 4842 7578 4860
rect 7560 4860 7578 4878
rect 7560 4878 7578 4896
rect 7560 4896 7578 4914
rect 7560 4914 7578 4932
rect 7560 4932 7578 4950
rect 7560 4950 7578 4968
rect 7560 4968 7578 4986
rect 7560 4986 7578 5004
rect 7560 5004 7578 5022
rect 7560 5022 7578 5040
rect 7560 5040 7578 5058
rect 7560 5058 7578 5076
rect 7560 5076 7578 5094
rect 7560 5094 7578 5112
rect 7560 5112 7578 5130
rect 7560 5130 7578 5148
rect 7560 5148 7578 5166
rect 7560 5166 7578 5184
rect 7560 5184 7578 5202
rect 7560 5202 7578 5220
rect 7560 5220 7578 5238
rect 7560 5238 7578 5256
rect 7560 5256 7578 5274
rect 7560 5274 7578 5292
rect 7560 5292 7578 5310
rect 7560 5310 7578 5328
rect 7560 5328 7578 5346
rect 7560 5346 7578 5364
rect 7560 5364 7578 5382
rect 7560 5382 7578 5400
rect 7560 5400 7578 5418
rect 7560 5418 7578 5436
rect 7560 5436 7578 5454
rect 7560 5454 7578 5472
rect 7560 5472 7578 5490
rect 7560 5490 7578 5508
rect 7560 5508 7578 5526
rect 7560 5526 7578 5544
rect 7560 5544 7578 5562
rect 7560 5562 7578 5580
rect 7560 5580 7578 5598
rect 7560 5598 7578 5616
rect 7560 5616 7578 5634
rect 7560 5634 7578 5652
rect 7560 5652 7578 5670
rect 7560 5670 7578 5688
rect 7560 5688 7578 5706
rect 7560 5706 7578 5724
rect 7560 5724 7578 5742
rect 7560 5742 7578 5760
rect 7560 5760 7578 5778
rect 7560 5778 7578 5796
rect 7560 5796 7578 5814
rect 7560 5814 7578 5832
rect 7560 5832 7578 5850
rect 7560 5850 7578 5868
rect 7560 5868 7578 5886
rect 7560 5886 7578 5904
rect 7560 5904 7578 5922
rect 7560 5922 7578 5940
rect 7560 5940 7578 5958
rect 7560 5958 7578 5976
rect 7560 5976 7578 5994
rect 7560 5994 7578 6012
rect 7560 6012 7578 6030
rect 7560 6030 7578 6048
rect 7560 6048 7578 6066
rect 7560 6066 7578 6084
rect 7560 6084 7578 6102
rect 7560 6102 7578 6120
rect 7560 6120 7578 6138
rect 7560 6138 7578 6156
rect 7560 6156 7578 6174
rect 7560 6174 7578 6192
rect 7560 6192 7578 6210
rect 7560 6210 7578 6228
rect 7560 6228 7578 6246
rect 7560 6246 7578 6264
rect 7560 6264 7578 6282
rect 7560 6282 7578 6300
rect 7560 6300 7578 6318
rect 7560 6318 7578 6336
rect 7560 6336 7578 6354
rect 7560 6354 7578 6372
rect 7560 6372 7578 6390
rect 7560 6390 7578 6408
rect 7560 6408 7578 6426
rect 7560 6426 7578 6444
rect 7560 6444 7578 6462
rect 7560 6462 7578 6480
rect 7560 6480 7578 6498
rect 7560 6498 7578 6516
rect 7560 6516 7578 6534
rect 7560 6534 7578 6552
rect 7560 6552 7578 6570
rect 7560 6570 7578 6588
rect 7560 6588 7578 6606
rect 7560 6606 7578 6624
rect 7560 6624 7578 6642
rect 7560 6642 7578 6660
rect 7560 6660 7578 6678
rect 7560 6678 7578 6696
rect 7578 2142 7596 2160
rect 7578 2160 7596 2178
rect 7578 2178 7596 2196
rect 7578 2196 7596 2214
rect 7578 2214 7596 2232
rect 7578 2232 7596 2250
rect 7578 2250 7596 2268
rect 7578 2268 7596 2286
rect 7578 2286 7596 2304
rect 7578 2304 7596 2322
rect 7578 2322 7596 2340
rect 7578 2340 7596 2358
rect 7578 2358 7596 2376
rect 7578 2376 7596 2394
rect 7578 2394 7596 2412
rect 7578 2412 7596 2430
rect 7578 2430 7596 2448
rect 7578 2448 7596 2466
rect 7578 2466 7596 2484
rect 7578 2484 7596 2502
rect 7578 2502 7596 2520
rect 7578 2520 7596 2538
rect 7578 2538 7596 2556
rect 7578 2556 7596 2574
rect 7578 2574 7596 2592
rect 7578 2592 7596 2610
rect 7578 2610 7596 2628
rect 7578 2628 7596 2646
rect 7578 2646 7596 2664
rect 7578 2664 7596 2682
rect 7578 2682 7596 2700
rect 7578 2700 7596 2718
rect 7578 2718 7596 2736
rect 7578 2736 7596 2754
rect 7578 2754 7596 2772
rect 7578 2772 7596 2790
rect 7578 2790 7596 2808
rect 7578 2808 7596 2826
rect 7578 2826 7596 2844
rect 7578 2844 7596 2862
rect 7578 2862 7596 2880
rect 7578 2880 7596 2898
rect 7578 2898 7596 2916
rect 7578 2916 7596 2934
rect 7578 2934 7596 2952
rect 7578 2952 7596 2970
rect 7578 2970 7596 2988
rect 7578 2988 7596 3006
rect 7578 3006 7596 3024
rect 7578 3024 7596 3042
rect 7578 3042 7596 3060
rect 7578 3060 7596 3078
rect 7578 3078 7596 3096
rect 7578 3096 7596 3114
rect 7578 3114 7596 3132
rect 7578 3132 7596 3150
rect 7578 3150 7596 3168
rect 7578 3168 7596 3186
rect 7578 3186 7596 3204
rect 7578 3204 7596 3222
rect 7578 3222 7596 3240
rect 7578 3240 7596 3258
rect 7578 4734 7596 4752
rect 7578 4752 7596 4770
rect 7578 4770 7596 4788
rect 7578 4788 7596 4806
rect 7578 4806 7596 4824
rect 7578 4824 7596 4842
rect 7578 4842 7596 4860
rect 7578 4860 7596 4878
rect 7578 4878 7596 4896
rect 7578 4896 7596 4914
rect 7578 4914 7596 4932
rect 7578 4932 7596 4950
rect 7578 4950 7596 4968
rect 7578 4968 7596 4986
rect 7578 4986 7596 5004
rect 7578 5004 7596 5022
rect 7578 5022 7596 5040
rect 7578 5040 7596 5058
rect 7578 5058 7596 5076
rect 7578 5076 7596 5094
rect 7578 5094 7596 5112
rect 7578 5112 7596 5130
rect 7578 5130 7596 5148
rect 7578 5148 7596 5166
rect 7578 5166 7596 5184
rect 7578 5184 7596 5202
rect 7578 5202 7596 5220
rect 7578 5220 7596 5238
rect 7578 5238 7596 5256
rect 7578 5256 7596 5274
rect 7578 5274 7596 5292
rect 7578 5292 7596 5310
rect 7578 5310 7596 5328
rect 7578 5328 7596 5346
rect 7578 5346 7596 5364
rect 7578 5364 7596 5382
rect 7578 5382 7596 5400
rect 7578 5400 7596 5418
rect 7578 5418 7596 5436
rect 7578 5436 7596 5454
rect 7578 5454 7596 5472
rect 7578 5472 7596 5490
rect 7578 5490 7596 5508
rect 7578 5508 7596 5526
rect 7578 5526 7596 5544
rect 7578 5544 7596 5562
rect 7578 5562 7596 5580
rect 7578 5580 7596 5598
rect 7578 5598 7596 5616
rect 7578 5616 7596 5634
rect 7578 5634 7596 5652
rect 7578 5652 7596 5670
rect 7578 5670 7596 5688
rect 7578 5688 7596 5706
rect 7578 5706 7596 5724
rect 7578 5724 7596 5742
rect 7578 5742 7596 5760
rect 7578 5760 7596 5778
rect 7578 5778 7596 5796
rect 7578 5796 7596 5814
rect 7578 5814 7596 5832
rect 7578 5832 7596 5850
rect 7578 5850 7596 5868
rect 7578 5868 7596 5886
rect 7578 5886 7596 5904
rect 7578 5904 7596 5922
rect 7578 5922 7596 5940
rect 7578 5940 7596 5958
rect 7578 5958 7596 5976
rect 7578 5976 7596 5994
rect 7578 5994 7596 6012
rect 7578 6012 7596 6030
rect 7578 6030 7596 6048
rect 7578 6048 7596 6066
rect 7578 6066 7596 6084
rect 7578 6084 7596 6102
rect 7578 6102 7596 6120
rect 7578 6120 7596 6138
rect 7578 6138 7596 6156
rect 7578 6156 7596 6174
rect 7578 6174 7596 6192
rect 7578 6192 7596 6210
rect 7578 6210 7596 6228
rect 7578 6228 7596 6246
rect 7578 6246 7596 6264
rect 7578 6264 7596 6282
rect 7578 6282 7596 6300
rect 7578 6300 7596 6318
rect 7578 6318 7596 6336
rect 7578 6336 7596 6354
rect 7578 6354 7596 6372
rect 7578 6372 7596 6390
rect 7578 6390 7596 6408
rect 7578 6408 7596 6426
rect 7578 6426 7596 6444
rect 7578 6444 7596 6462
rect 7578 6462 7596 6480
rect 7578 6480 7596 6498
rect 7578 6498 7596 6516
rect 7578 6516 7596 6534
rect 7578 6534 7596 6552
rect 7578 6552 7596 6570
rect 7578 6570 7596 6588
rect 7578 6588 7596 6606
rect 7578 6606 7596 6624
rect 7578 6624 7596 6642
rect 7578 6642 7596 6660
rect 7578 6660 7596 6678
rect 7578 6678 7596 6696
rect 7578 6696 7596 6714
rect 7596 2142 7614 2160
rect 7596 2160 7614 2178
rect 7596 2178 7614 2196
rect 7596 2196 7614 2214
rect 7596 2214 7614 2232
rect 7596 2232 7614 2250
rect 7596 2250 7614 2268
rect 7596 2268 7614 2286
rect 7596 2286 7614 2304
rect 7596 2304 7614 2322
rect 7596 2322 7614 2340
rect 7596 2340 7614 2358
rect 7596 2358 7614 2376
rect 7596 2376 7614 2394
rect 7596 2394 7614 2412
rect 7596 2412 7614 2430
rect 7596 2430 7614 2448
rect 7596 2448 7614 2466
rect 7596 2466 7614 2484
rect 7596 2484 7614 2502
rect 7596 2502 7614 2520
rect 7596 2520 7614 2538
rect 7596 2538 7614 2556
rect 7596 2556 7614 2574
rect 7596 2574 7614 2592
rect 7596 2592 7614 2610
rect 7596 2610 7614 2628
rect 7596 2628 7614 2646
rect 7596 2646 7614 2664
rect 7596 2664 7614 2682
rect 7596 2682 7614 2700
rect 7596 2700 7614 2718
rect 7596 2718 7614 2736
rect 7596 2736 7614 2754
rect 7596 2754 7614 2772
rect 7596 2772 7614 2790
rect 7596 2790 7614 2808
rect 7596 2808 7614 2826
rect 7596 2826 7614 2844
rect 7596 2844 7614 2862
rect 7596 2862 7614 2880
rect 7596 2880 7614 2898
rect 7596 2898 7614 2916
rect 7596 2916 7614 2934
rect 7596 2934 7614 2952
rect 7596 2952 7614 2970
rect 7596 2970 7614 2988
rect 7596 2988 7614 3006
rect 7596 3006 7614 3024
rect 7596 3024 7614 3042
rect 7596 3042 7614 3060
rect 7596 3060 7614 3078
rect 7596 3078 7614 3096
rect 7596 3096 7614 3114
rect 7596 3114 7614 3132
rect 7596 3132 7614 3150
rect 7596 3150 7614 3168
rect 7596 3168 7614 3186
rect 7596 3186 7614 3204
rect 7596 3204 7614 3222
rect 7596 3222 7614 3240
rect 7596 3240 7614 3258
rect 7596 4770 7614 4788
rect 7596 4788 7614 4806
rect 7596 4806 7614 4824
rect 7596 4824 7614 4842
rect 7596 4842 7614 4860
rect 7596 4860 7614 4878
rect 7596 4878 7614 4896
rect 7596 4896 7614 4914
rect 7596 4914 7614 4932
rect 7596 4932 7614 4950
rect 7596 4950 7614 4968
rect 7596 4968 7614 4986
rect 7596 4986 7614 5004
rect 7596 5004 7614 5022
rect 7596 5022 7614 5040
rect 7596 5040 7614 5058
rect 7596 5058 7614 5076
rect 7596 5076 7614 5094
rect 7596 5094 7614 5112
rect 7596 5112 7614 5130
rect 7596 5130 7614 5148
rect 7596 5148 7614 5166
rect 7596 5166 7614 5184
rect 7596 5184 7614 5202
rect 7596 5202 7614 5220
rect 7596 5220 7614 5238
rect 7596 5238 7614 5256
rect 7596 5256 7614 5274
rect 7596 5274 7614 5292
rect 7596 5292 7614 5310
rect 7596 5310 7614 5328
rect 7596 5328 7614 5346
rect 7596 5346 7614 5364
rect 7596 5364 7614 5382
rect 7596 5382 7614 5400
rect 7596 5400 7614 5418
rect 7596 5418 7614 5436
rect 7596 5436 7614 5454
rect 7596 5454 7614 5472
rect 7596 5472 7614 5490
rect 7596 5490 7614 5508
rect 7596 5508 7614 5526
rect 7596 5526 7614 5544
rect 7596 5544 7614 5562
rect 7596 5562 7614 5580
rect 7596 5580 7614 5598
rect 7596 5598 7614 5616
rect 7596 5616 7614 5634
rect 7596 5634 7614 5652
rect 7596 5652 7614 5670
rect 7596 5670 7614 5688
rect 7596 5688 7614 5706
rect 7596 5706 7614 5724
rect 7596 5724 7614 5742
rect 7596 5742 7614 5760
rect 7596 5760 7614 5778
rect 7596 5778 7614 5796
rect 7596 5796 7614 5814
rect 7596 5814 7614 5832
rect 7596 5832 7614 5850
rect 7596 5850 7614 5868
rect 7596 5868 7614 5886
rect 7596 5886 7614 5904
rect 7596 5904 7614 5922
rect 7596 5922 7614 5940
rect 7596 5940 7614 5958
rect 7596 5958 7614 5976
rect 7596 5976 7614 5994
rect 7596 5994 7614 6012
rect 7596 6012 7614 6030
rect 7596 6030 7614 6048
rect 7596 6048 7614 6066
rect 7596 6066 7614 6084
rect 7596 6084 7614 6102
rect 7596 6102 7614 6120
rect 7596 6120 7614 6138
rect 7596 6138 7614 6156
rect 7596 6156 7614 6174
rect 7596 6174 7614 6192
rect 7596 6192 7614 6210
rect 7596 6210 7614 6228
rect 7596 6228 7614 6246
rect 7596 6246 7614 6264
rect 7596 6264 7614 6282
rect 7596 6282 7614 6300
rect 7596 6300 7614 6318
rect 7596 6318 7614 6336
rect 7596 6336 7614 6354
rect 7596 6354 7614 6372
rect 7596 6372 7614 6390
rect 7596 6390 7614 6408
rect 7596 6408 7614 6426
rect 7596 6426 7614 6444
rect 7596 6444 7614 6462
rect 7596 6462 7614 6480
rect 7596 6480 7614 6498
rect 7596 6498 7614 6516
rect 7596 6516 7614 6534
rect 7596 6534 7614 6552
rect 7596 6552 7614 6570
rect 7596 6570 7614 6588
rect 7596 6588 7614 6606
rect 7596 6606 7614 6624
rect 7596 6624 7614 6642
rect 7596 6642 7614 6660
rect 7596 6660 7614 6678
rect 7596 6678 7614 6696
rect 7596 6696 7614 6714
rect 7596 6714 7614 6732
rect 7614 2160 7632 2178
rect 7614 2178 7632 2196
rect 7614 2196 7632 2214
rect 7614 2214 7632 2232
rect 7614 2232 7632 2250
rect 7614 2250 7632 2268
rect 7614 2268 7632 2286
rect 7614 2286 7632 2304
rect 7614 2304 7632 2322
rect 7614 2322 7632 2340
rect 7614 2340 7632 2358
rect 7614 2358 7632 2376
rect 7614 2376 7632 2394
rect 7614 2394 7632 2412
rect 7614 2412 7632 2430
rect 7614 2430 7632 2448
rect 7614 2448 7632 2466
rect 7614 2466 7632 2484
rect 7614 2484 7632 2502
rect 7614 2502 7632 2520
rect 7614 2520 7632 2538
rect 7614 2538 7632 2556
rect 7614 2556 7632 2574
rect 7614 2574 7632 2592
rect 7614 2592 7632 2610
rect 7614 2610 7632 2628
rect 7614 2628 7632 2646
rect 7614 2646 7632 2664
rect 7614 2664 7632 2682
rect 7614 2682 7632 2700
rect 7614 2700 7632 2718
rect 7614 2718 7632 2736
rect 7614 2736 7632 2754
rect 7614 2754 7632 2772
rect 7614 2772 7632 2790
rect 7614 2790 7632 2808
rect 7614 2808 7632 2826
rect 7614 2826 7632 2844
rect 7614 2844 7632 2862
rect 7614 2862 7632 2880
rect 7614 2880 7632 2898
rect 7614 2898 7632 2916
rect 7614 2916 7632 2934
rect 7614 2934 7632 2952
rect 7614 2952 7632 2970
rect 7614 2970 7632 2988
rect 7614 2988 7632 3006
rect 7614 3006 7632 3024
rect 7614 3024 7632 3042
rect 7614 3042 7632 3060
rect 7614 3060 7632 3078
rect 7614 3078 7632 3096
rect 7614 3096 7632 3114
rect 7614 3114 7632 3132
rect 7614 3132 7632 3150
rect 7614 3150 7632 3168
rect 7614 3168 7632 3186
rect 7614 3186 7632 3204
rect 7614 3204 7632 3222
rect 7614 3222 7632 3240
rect 7614 3240 7632 3258
rect 7614 4788 7632 4806
rect 7614 4806 7632 4824
rect 7614 4824 7632 4842
rect 7614 4842 7632 4860
rect 7614 4860 7632 4878
rect 7614 4878 7632 4896
rect 7614 4896 7632 4914
rect 7614 4914 7632 4932
rect 7614 4932 7632 4950
rect 7614 4950 7632 4968
rect 7614 4968 7632 4986
rect 7614 4986 7632 5004
rect 7614 5004 7632 5022
rect 7614 5022 7632 5040
rect 7614 5040 7632 5058
rect 7614 5058 7632 5076
rect 7614 5076 7632 5094
rect 7614 5094 7632 5112
rect 7614 5112 7632 5130
rect 7614 5130 7632 5148
rect 7614 5148 7632 5166
rect 7614 5166 7632 5184
rect 7614 5184 7632 5202
rect 7614 5202 7632 5220
rect 7614 5220 7632 5238
rect 7614 5238 7632 5256
rect 7614 5256 7632 5274
rect 7614 5274 7632 5292
rect 7614 5292 7632 5310
rect 7614 5310 7632 5328
rect 7614 5328 7632 5346
rect 7614 5346 7632 5364
rect 7614 5364 7632 5382
rect 7614 5382 7632 5400
rect 7614 5400 7632 5418
rect 7614 5418 7632 5436
rect 7614 5436 7632 5454
rect 7614 5454 7632 5472
rect 7614 5472 7632 5490
rect 7614 5490 7632 5508
rect 7614 5508 7632 5526
rect 7614 5526 7632 5544
rect 7614 5544 7632 5562
rect 7614 5562 7632 5580
rect 7614 5580 7632 5598
rect 7614 5598 7632 5616
rect 7614 5616 7632 5634
rect 7614 5634 7632 5652
rect 7614 5652 7632 5670
rect 7614 5670 7632 5688
rect 7614 5688 7632 5706
rect 7614 5706 7632 5724
rect 7614 5724 7632 5742
rect 7614 5742 7632 5760
rect 7614 5760 7632 5778
rect 7614 5778 7632 5796
rect 7614 5796 7632 5814
rect 7614 5814 7632 5832
rect 7614 5832 7632 5850
rect 7614 5850 7632 5868
rect 7614 5868 7632 5886
rect 7614 5886 7632 5904
rect 7614 5904 7632 5922
rect 7614 5922 7632 5940
rect 7614 5940 7632 5958
rect 7614 5958 7632 5976
rect 7614 5976 7632 5994
rect 7614 5994 7632 6012
rect 7614 6012 7632 6030
rect 7614 6030 7632 6048
rect 7614 6048 7632 6066
rect 7614 6066 7632 6084
rect 7614 6084 7632 6102
rect 7614 6102 7632 6120
rect 7614 6120 7632 6138
rect 7614 6138 7632 6156
rect 7614 6156 7632 6174
rect 7614 6174 7632 6192
rect 7614 6192 7632 6210
rect 7614 6210 7632 6228
rect 7614 6228 7632 6246
rect 7614 6246 7632 6264
rect 7614 6264 7632 6282
rect 7614 6282 7632 6300
rect 7614 6300 7632 6318
rect 7614 6318 7632 6336
rect 7614 6336 7632 6354
rect 7614 6354 7632 6372
rect 7614 6372 7632 6390
rect 7614 6390 7632 6408
rect 7614 6408 7632 6426
rect 7614 6426 7632 6444
rect 7614 6444 7632 6462
rect 7614 6462 7632 6480
rect 7614 6480 7632 6498
rect 7614 6498 7632 6516
rect 7614 6516 7632 6534
rect 7614 6534 7632 6552
rect 7614 6552 7632 6570
rect 7614 6570 7632 6588
rect 7614 6588 7632 6606
rect 7614 6606 7632 6624
rect 7614 6624 7632 6642
rect 7614 6642 7632 6660
rect 7614 6660 7632 6678
rect 7614 6678 7632 6696
rect 7614 6696 7632 6714
rect 7614 6714 7632 6732
rect 7614 6732 7632 6750
rect 7632 2160 7650 2178
rect 7632 2178 7650 2196
rect 7632 2196 7650 2214
rect 7632 2214 7650 2232
rect 7632 2232 7650 2250
rect 7632 2250 7650 2268
rect 7632 2268 7650 2286
rect 7632 2286 7650 2304
rect 7632 2304 7650 2322
rect 7632 2322 7650 2340
rect 7632 2340 7650 2358
rect 7632 2358 7650 2376
rect 7632 2376 7650 2394
rect 7632 2394 7650 2412
rect 7632 2412 7650 2430
rect 7632 2430 7650 2448
rect 7632 2448 7650 2466
rect 7632 2466 7650 2484
rect 7632 2484 7650 2502
rect 7632 2502 7650 2520
rect 7632 2520 7650 2538
rect 7632 2538 7650 2556
rect 7632 2556 7650 2574
rect 7632 2574 7650 2592
rect 7632 2592 7650 2610
rect 7632 2610 7650 2628
rect 7632 2628 7650 2646
rect 7632 2646 7650 2664
rect 7632 2664 7650 2682
rect 7632 2682 7650 2700
rect 7632 2700 7650 2718
rect 7632 2718 7650 2736
rect 7632 2736 7650 2754
rect 7632 2754 7650 2772
rect 7632 2772 7650 2790
rect 7632 2790 7650 2808
rect 7632 2808 7650 2826
rect 7632 2826 7650 2844
rect 7632 2844 7650 2862
rect 7632 2862 7650 2880
rect 7632 2880 7650 2898
rect 7632 2898 7650 2916
rect 7632 2916 7650 2934
rect 7632 2934 7650 2952
rect 7632 2952 7650 2970
rect 7632 2970 7650 2988
rect 7632 2988 7650 3006
rect 7632 3006 7650 3024
rect 7632 3024 7650 3042
rect 7632 3042 7650 3060
rect 7632 3060 7650 3078
rect 7632 3078 7650 3096
rect 7632 3096 7650 3114
rect 7632 3114 7650 3132
rect 7632 3132 7650 3150
rect 7632 3150 7650 3168
rect 7632 3168 7650 3186
rect 7632 3186 7650 3204
rect 7632 3204 7650 3222
rect 7632 3222 7650 3240
rect 7632 3240 7650 3258
rect 7632 3258 7650 3276
rect 7632 4806 7650 4824
rect 7632 4824 7650 4842
rect 7632 4842 7650 4860
rect 7632 4860 7650 4878
rect 7632 4878 7650 4896
rect 7632 4896 7650 4914
rect 7632 4914 7650 4932
rect 7632 4932 7650 4950
rect 7632 4950 7650 4968
rect 7632 4968 7650 4986
rect 7632 4986 7650 5004
rect 7632 5004 7650 5022
rect 7632 5022 7650 5040
rect 7632 5040 7650 5058
rect 7632 5058 7650 5076
rect 7632 5076 7650 5094
rect 7632 5094 7650 5112
rect 7632 5112 7650 5130
rect 7632 5130 7650 5148
rect 7632 5148 7650 5166
rect 7632 5166 7650 5184
rect 7632 5184 7650 5202
rect 7632 5202 7650 5220
rect 7632 5220 7650 5238
rect 7632 5238 7650 5256
rect 7632 5256 7650 5274
rect 7632 5274 7650 5292
rect 7632 5292 7650 5310
rect 7632 5310 7650 5328
rect 7632 5328 7650 5346
rect 7632 5346 7650 5364
rect 7632 5364 7650 5382
rect 7632 5382 7650 5400
rect 7632 5400 7650 5418
rect 7632 5418 7650 5436
rect 7632 5436 7650 5454
rect 7632 5454 7650 5472
rect 7632 5472 7650 5490
rect 7632 5490 7650 5508
rect 7632 5508 7650 5526
rect 7632 5526 7650 5544
rect 7632 5544 7650 5562
rect 7632 5562 7650 5580
rect 7632 5580 7650 5598
rect 7632 5598 7650 5616
rect 7632 5616 7650 5634
rect 7632 5634 7650 5652
rect 7632 5652 7650 5670
rect 7632 5670 7650 5688
rect 7632 5688 7650 5706
rect 7632 5706 7650 5724
rect 7632 5724 7650 5742
rect 7632 5742 7650 5760
rect 7632 5760 7650 5778
rect 7632 5778 7650 5796
rect 7632 5796 7650 5814
rect 7632 5814 7650 5832
rect 7632 5832 7650 5850
rect 7632 5850 7650 5868
rect 7632 5868 7650 5886
rect 7632 5886 7650 5904
rect 7632 5904 7650 5922
rect 7632 5922 7650 5940
rect 7632 5940 7650 5958
rect 7632 5958 7650 5976
rect 7632 5976 7650 5994
rect 7632 5994 7650 6012
rect 7632 6012 7650 6030
rect 7632 6030 7650 6048
rect 7632 6048 7650 6066
rect 7632 6066 7650 6084
rect 7632 6084 7650 6102
rect 7632 6102 7650 6120
rect 7632 6120 7650 6138
rect 7632 6138 7650 6156
rect 7632 6156 7650 6174
rect 7632 6174 7650 6192
rect 7632 6192 7650 6210
rect 7632 6210 7650 6228
rect 7632 6228 7650 6246
rect 7632 6246 7650 6264
rect 7632 6264 7650 6282
rect 7632 6282 7650 6300
rect 7632 6300 7650 6318
rect 7632 6318 7650 6336
rect 7632 6336 7650 6354
rect 7632 6354 7650 6372
rect 7632 6372 7650 6390
rect 7632 6390 7650 6408
rect 7632 6408 7650 6426
rect 7632 6426 7650 6444
rect 7632 6444 7650 6462
rect 7632 6462 7650 6480
rect 7632 6480 7650 6498
rect 7632 6498 7650 6516
rect 7632 6516 7650 6534
rect 7632 6534 7650 6552
rect 7632 6552 7650 6570
rect 7632 6570 7650 6588
rect 7632 6588 7650 6606
rect 7632 6606 7650 6624
rect 7632 6624 7650 6642
rect 7632 6642 7650 6660
rect 7632 6660 7650 6678
rect 7632 6678 7650 6696
rect 7632 6696 7650 6714
rect 7632 6714 7650 6732
rect 7632 6732 7650 6750
rect 7650 2178 7668 2196
rect 7650 2196 7668 2214
rect 7650 2214 7668 2232
rect 7650 2232 7668 2250
rect 7650 2250 7668 2268
rect 7650 2268 7668 2286
rect 7650 2286 7668 2304
rect 7650 2304 7668 2322
rect 7650 2322 7668 2340
rect 7650 2340 7668 2358
rect 7650 2358 7668 2376
rect 7650 2376 7668 2394
rect 7650 2394 7668 2412
rect 7650 2412 7668 2430
rect 7650 2430 7668 2448
rect 7650 2448 7668 2466
rect 7650 2466 7668 2484
rect 7650 2484 7668 2502
rect 7650 2502 7668 2520
rect 7650 2520 7668 2538
rect 7650 2538 7668 2556
rect 7650 2556 7668 2574
rect 7650 2574 7668 2592
rect 7650 2592 7668 2610
rect 7650 2610 7668 2628
rect 7650 2628 7668 2646
rect 7650 2646 7668 2664
rect 7650 2664 7668 2682
rect 7650 2682 7668 2700
rect 7650 2700 7668 2718
rect 7650 2718 7668 2736
rect 7650 2736 7668 2754
rect 7650 2754 7668 2772
rect 7650 2772 7668 2790
rect 7650 2790 7668 2808
rect 7650 2808 7668 2826
rect 7650 2826 7668 2844
rect 7650 2844 7668 2862
rect 7650 2862 7668 2880
rect 7650 2880 7668 2898
rect 7650 2898 7668 2916
rect 7650 2916 7668 2934
rect 7650 2934 7668 2952
rect 7650 2952 7668 2970
rect 7650 2970 7668 2988
rect 7650 2988 7668 3006
rect 7650 3006 7668 3024
rect 7650 3024 7668 3042
rect 7650 3042 7668 3060
rect 7650 3060 7668 3078
rect 7650 3078 7668 3096
rect 7650 3096 7668 3114
rect 7650 3114 7668 3132
rect 7650 3132 7668 3150
rect 7650 3150 7668 3168
rect 7650 3168 7668 3186
rect 7650 3186 7668 3204
rect 7650 3204 7668 3222
rect 7650 3222 7668 3240
rect 7650 3240 7668 3258
rect 7650 3258 7668 3276
rect 7650 4824 7668 4842
rect 7650 4842 7668 4860
rect 7650 4860 7668 4878
rect 7650 4878 7668 4896
rect 7650 4896 7668 4914
rect 7650 4914 7668 4932
rect 7650 4932 7668 4950
rect 7650 4950 7668 4968
rect 7650 4968 7668 4986
rect 7650 4986 7668 5004
rect 7650 5004 7668 5022
rect 7650 5022 7668 5040
rect 7650 5040 7668 5058
rect 7650 5058 7668 5076
rect 7650 5076 7668 5094
rect 7650 5094 7668 5112
rect 7650 5112 7668 5130
rect 7650 5130 7668 5148
rect 7650 5148 7668 5166
rect 7650 5166 7668 5184
rect 7650 5184 7668 5202
rect 7650 5202 7668 5220
rect 7650 5220 7668 5238
rect 7650 5238 7668 5256
rect 7650 5256 7668 5274
rect 7650 5274 7668 5292
rect 7650 5292 7668 5310
rect 7650 5310 7668 5328
rect 7650 5328 7668 5346
rect 7650 5346 7668 5364
rect 7650 5364 7668 5382
rect 7650 5382 7668 5400
rect 7650 5400 7668 5418
rect 7650 5418 7668 5436
rect 7650 5436 7668 5454
rect 7650 5454 7668 5472
rect 7650 5472 7668 5490
rect 7650 5490 7668 5508
rect 7650 5508 7668 5526
rect 7650 5526 7668 5544
rect 7650 5544 7668 5562
rect 7650 5562 7668 5580
rect 7650 5580 7668 5598
rect 7650 5598 7668 5616
rect 7650 5616 7668 5634
rect 7650 5634 7668 5652
rect 7650 5652 7668 5670
rect 7650 5670 7668 5688
rect 7650 5688 7668 5706
rect 7650 5706 7668 5724
rect 7650 5724 7668 5742
rect 7650 5742 7668 5760
rect 7650 5760 7668 5778
rect 7650 5778 7668 5796
rect 7650 5796 7668 5814
rect 7650 5814 7668 5832
rect 7650 5832 7668 5850
rect 7650 5850 7668 5868
rect 7650 5868 7668 5886
rect 7650 5886 7668 5904
rect 7650 5904 7668 5922
rect 7650 5922 7668 5940
rect 7650 5940 7668 5958
rect 7650 5958 7668 5976
rect 7650 5976 7668 5994
rect 7650 5994 7668 6012
rect 7650 6012 7668 6030
rect 7650 6030 7668 6048
rect 7650 6048 7668 6066
rect 7650 6066 7668 6084
rect 7650 6084 7668 6102
rect 7650 6102 7668 6120
rect 7650 6120 7668 6138
rect 7650 6138 7668 6156
rect 7650 6156 7668 6174
rect 7650 6174 7668 6192
rect 7650 6192 7668 6210
rect 7650 6210 7668 6228
rect 7650 6228 7668 6246
rect 7650 6246 7668 6264
rect 7650 6264 7668 6282
rect 7650 6282 7668 6300
rect 7650 6300 7668 6318
rect 7650 6318 7668 6336
rect 7650 6336 7668 6354
rect 7650 6354 7668 6372
rect 7650 6372 7668 6390
rect 7650 6390 7668 6408
rect 7650 6408 7668 6426
rect 7650 6426 7668 6444
rect 7650 6444 7668 6462
rect 7650 6462 7668 6480
rect 7650 6480 7668 6498
rect 7650 6498 7668 6516
rect 7650 6516 7668 6534
rect 7650 6534 7668 6552
rect 7650 6552 7668 6570
rect 7650 6570 7668 6588
rect 7650 6588 7668 6606
rect 7650 6606 7668 6624
rect 7650 6624 7668 6642
rect 7650 6642 7668 6660
rect 7650 6660 7668 6678
rect 7650 6678 7668 6696
rect 7650 6696 7668 6714
rect 7650 6714 7668 6732
rect 7650 6732 7668 6750
rect 7650 6750 7668 6768
rect 7668 2196 7686 2214
rect 7668 2214 7686 2232
rect 7668 2232 7686 2250
rect 7668 2250 7686 2268
rect 7668 2268 7686 2286
rect 7668 2286 7686 2304
rect 7668 2304 7686 2322
rect 7668 2322 7686 2340
rect 7668 2340 7686 2358
rect 7668 2358 7686 2376
rect 7668 2376 7686 2394
rect 7668 2394 7686 2412
rect 7668 2412 7686 2430
rect 7668 2430 7686 2448
rect 7668 2448 7686 2466
rect 7668 2466 7686 2484
rect 7668 2484 7686 2502
rect 7668 2502 7686 2520
rect 7668 2520 7686 2538
rect 7668 2538 7686 2556
rect 7668 2556 7686 2574
rect 7668 2574 7686 2592
rect 7668 2592 7686 2610
rect 7668 2610 7686 2628
rect 7668 2628 7686 2646
rect 7668 2646 7686 2664
rect 7668 2664 7686 2682
rect 7668 2682 7686 2700
rect 7668 2700 7686 2718
rect 7668 2718 7686 2736
rect 7668 2736 7686 2754
rect 7668 2754 7686 2772
rect 7668 2772 7686 2790
rect 7668 2790 7686 2808
rect 7668 2808 7686 2826
rect 7668 2826 7686 2844
rect 7668 2844 7686 2862
rect 7668 2862 7686 2880
rect 7668 2880 7686 2898
rect 7668 2898 7686 2916
rect 7668 2916 7686 2934
rect 7668 2934 7686 2952
rect 7668 2952 7686 2970
rect 7668 2970 7686 2988
rect 7668 2988 7686 3006
rect 7668 3006 7686 3024
rect 7668 3024 7686 3042
rect 7668 3042 7686 3060
rect 7668 3060 7686 3078
rect 7668 3078 7686 3096
rect 7668 3096 7686 3114
rect 7668 3114 7686 3132
rect 7668 3132 7686 3150
rect 7668 3150 7686 3168
rect 7668 3168 7686 3186
rect 7668 3186 7686 3204
rect 7668 3204 7686 3222
rect 7668 3222 7686 3240
rect 7668 3240 7686 3258
rect 7668 3258 7686 3276
rect 7668 4842 7686 4860
rect 7668 4860 7686 4878
rect 7668 4878 7686 4896
rect 7668 4896 7686 4914
rect 7668 4914 7686 4932
rect 7668 4932 7686 4950
rect 7668 4950 7686 4968
rect 7668 4968 7686 4986
rect 7668 4986 7686 5004
rect 7668 5004 7686 5022
rect 7668 5022 7686 5040
rect 7668 5040 7686 5058
rect 7668 5058 7686 5076
rect 7668 5076 7686 5094
rect 7668 5094 7686 5112
rect 7668 5112 7686 5130
rect 7668 5130 7686 5148
rect 7668 5148 7686 5166
rect 7668 5166 7686 5184
rect 7668 5184 7686 5202
rect 7668 5202 7686 5220
rect 7668 5220 7686 5238
rect 7668 5238 7686 5256
rect 7668 5256 7686 5274
rect 7668 5274 7686 5292
rect 7668 5292 7686 5310
rect 7668 5310 7686 5328
rect 7668 5328 7686 5346
rect 7668 5346 7686 5364
rect 7668 5364 7686 5382
rect 7668 5382 7686 5400
rect 7668 5400 7686 5418
rect 7668 5418 7686 5436
rect 7668 5436 7686 5454
rect 7668 5454 7686 5472
rect 7668 5472 7686 5490
rect 7668 5490 7686 5508
rect 7668 5508 7686 5526
rect 7668 5526 7686 5544
rect 7668 5544 7686 5562
rect 7668 5562 7686 5580
rect 7668 5580 7686 5598
rect 7668 5598 7686 5616
rect 7668 5616 7686 5634
rect 7668 5634 7686 5652
rect 7668 5652 7686 5670
rect 7668 5670 7686 5688
rect 7668 5688 7686 5706
rect 7668 5706 7686 5724
rect 7668 5724 7686 5742
rect 7668 5742 7686 5760
rect 7668 5760 7686 5778
rect 7668 5778 7686 5796
rect 7668 5796 7686 5814
rect 7668 5814 7686 5832
rect 7668 5832 7686 5850
rect 7668 5850 7686 5868
rect 7668 5868 7686 5886
rect 7668 5886 7686 5904
rect 7668 5904 7686 5922
rect 7668 5922 7686 5940
rect 7668 5940 7686 5958
rect 7668 5958 7686 5976
rect 7668 5976 7686 5994
rect 7668 5994 7686 6012
rect 7668 6012 7686 6030
rect 7668 6030 7686 6048
rect 7668 6048 7686 6066
rect 7668 6066 7686 6084
rect 7668 6084 7686 6102
rect 7668 6102 7686 6120
rect 7668 6120 7686 6138
rect 7668 6138 7686 6156
rect 7668 6156 7686 6174
rect 7668 6174 7686 6192
rect 7668 6192 7686 6210
rect 7668 6210 7686 6228
rect 7668 6228 7686 6246
rect 7668 6246 7686 6264
rect 7668 6264 7686 6282
rect 7668 6282 7686 6300
rect 7668 6300 7686 6318
rect 7668 6318 7686 6336
rect 7668 6336 7686 6354
rect 7668 6354 7686 6372
rect 7668 6372 7686 6390
rect 7668 6390 7686 6408
rect 7668 6408 7686 6426
rect 7668 6426 7686 6444
rect 7668 6444 7686 6462
rect 7668 6462 7686 6480
rect 7668 6480 7686 6498
rect 7668 6498 7686 6516
rect 7668 6516 7686 6534
rect 7668 6534 7686 6552
rect 7668 6552 7686 6570
rect 7668 6570 7686 6588
rect 7668 6588 7686 6606
rect 7668 6606 7686 6624
rect 7668 6624 7686 6642
rect 7668 6642 7686 6660
rect 7668 6660 7686 6678
rect 7668 6678 7686 6696
rect 7668 6696 7686 6714
rect 7668 6714 7686 6732
rect 7668 6732 7686 6750
rect 7668 6750 7686 6768
rect 7668 6768 7686 6786
rect 7686 2196 7704 2214
rect 7686 2214 7704 2232
rect 7686 2232 7704 2250
rect 7686 2250 7704 2268
rect 7686 2268 7704 2286
rect 7686 2286 7704 2304
rect 7686 2304 7704 2322
rect 7686 2322 7704 2340
rect 7686 2340 7704 2358
rect 7686 2358 7704 2376
rect 7686 2376 7704 2394
rect 7686 2394 7704 2412
rect 7686 2412 7704 2430
rect 7686 2430 7704 2448
rect 7686 2448 7704 2466
rect 7686 2466 7704 2484
rect 7686 2484 7704 2502
rect 7686 2502 7704 2520
rect 7686 2520 7704 2538
rect 7686 2538 7704 2556
rect 7686 2556 7704 2574
rect 7686 2574 7704 2592
rect 7686 2592 7704 2610
rect 7686 2610 7704 2628
rect 7686 2628 7704 2646
rect 7686 2646 7704 2664
rect 7686 2664 7704 2682
rect 7686 2682 7704 2700
rect 7686 2700 7704 2718
rect 7686 2718 7704 2736
rect 7686 2736 7704 2754
rect 7686 2754 7704 2772
rect 7686 2772 7704 2790
rect 7686 2790 7704 2808
rect 7686 2808 7704 2826
rect 7686 2826 7704 2844
rect 7686 2844 7704 2862
rect 7686 2862 7704 2880
rect 7686 2880 7704 2898
rect 7686 2898 7704 2916
rect 7686 2916 7704 2934
rect 7686 2934 7704 2952
rect 7686 2952 7704 2970
rect 7686 2970 7704 2988
rect 7686 2988 7704 3006
rect 7686 3006 7704 3024
rect 7686 3024 7704 3042
rect 7686 3042 7704 3060
rect 7686 3060 7704 3078
rect 7686 3078 7704 3096
rect 7686 3096 7704 3114
rect 7686 3114 7704 3132
rect 7686 3132 7704 3150
rect 7686 3150 7704 3168
rect 7686 3168 7704 3186
rect 7686 3186 7704 3204
rect 7686 3204 7704 3222
rect 7686 3222 7704 3240
rect 7686 3240 7704 3258
rect 7686 3258 7704 3276
rect 7686 4878 7704 4896
rect 7686 4896 7704 4914
rect 7686 4914 7704 4932
rect 7686 4932 7704 4950
rect 7686 4950 7704 4968
rect 7686 4968 7704 4986
rect 7686 4986 7704 5004
rect 7686 5004 7704 5022
rect 7686 5022 7704 5040
rect 7686 5040 7704 5058
rect 7686 5058 7704 5076
rect 7686 5076 7704 5094
rect 7686 5094 7704 5112
rect 7686 5112 7704 5130
rect 7686 5130 7704 5148
rect 7686 5148 7704 5166
rect 7686 5166 7704 5184
rect 7686 5184 7704 5202
rect 7686 5202 7704 5220
rect 7686 5220 7704 5238
rect 7686 5238 7704 5256
rect 7686 5256 7704 5274
rect 7686 5274 7704 5292
rect 7686 5292 7704 5310
rect 7686 5310 7704 5328
rect 7686 5328 7704 5346
rect 7686 5346 7704 5364
rect 7686 5364 7704 5382
rect 7686 5382 7704 5400
rect 7686 5400 7704 5418
rect 7686 5418 7704 5436
rect 7686 5436 7704 5454
rect 7686 5454 7704 5472
rect 7686 5472 7704 5490
rect 7686 5490 7704 5508
rect 7686 5508 7704 5526
rect 7686 5526 7704 5544
rect 7686 5544 7704 5562
rect 7686 5562 7704 5580
rect 7686 5580 7704 5598
rect 7686 5598 7704 5616
rect 7686 5616 7704 5634
rect 7686 5634 7704 5652
rect 7686 5652 7704 5670
rect 7686 5670 7704 5688
rect 7686 5688 7704 5706
rect 7686 5706 7704 5724
rect 7686 5724 7704 5742
rect 7686 5742 7704 5760
rect 7686 5760 7704 5778
rect 7686 5778 7704 5796
rect 7686 5796 7704 5814
rect 7686 5814 7704 5832
rect 7686 5832 7704 5850
rect 7686 5850 7704 5868
rect 7686 5868 7704 5886
rect 7686 5886 7704 5904
rect 7686 5904 7704 5922
rect 7686 5922 7704 5940
rect 7686 5940 7704 5958
rect 7686 5958 7704 5976
rect 7686 5976 7704 5994
rect 7686 5994 7704 6012
rect 7686 6012 7704 6030
rect 7686 6030 7704 6048
rect 7686 6048 7704 6066
rect 7686 6066 7704 6084
rect 7686 6084 7704 6102
rect 7686 6102 7704 6120
rect 7686 6120 7704 6138
rect 7686 6138 7704 6156
rect 7686 6156 7704 6174
rect 7686 6174 7704 6192
rect 7686 6192 7704 6210
rect 7686 6210 7704 6228
rect 7686 6228 7704 6246
rect 7686 6246 7704 6264
rect 7686 6264 7704 6282
rect 7686 6282 7704 6300
rect 7686 6300 7704 6318
rect 7686 6318 7704 6336
rect 7686 6336 7704 6354
rect 7686 6354 7704 6372
rect 7686 6372 7704 6390
rect 7686 6390 7704 6408
rect 7686 6408 7704 6426
rect 7686 6426 7704 6444
rect 7686 6444 7704 6462
rect 7686 6462 7704 6480
rect 7686 6480 7704 6498
rect 7686 6498 7704 6516
rect 7686 6516 7704 6534
rect 7686 6534 7704 6552
rect 7686 6552 7704 6570
rect 7686 6570 7704 6588
rect 7686 6588 7704 6606
rect 7686 6606 7704 6624
rect 7686 6624 7704 6642
rect 7686 6642 7704 6660
rect 7686 6660 7704 6678
rect 7686 6678 7704 6696
rect 7686 6696 7704 6714
rect 7686 6714 7704 6732
rect 7686 6732 7704 6750
rect 7686 6750 7704 6768
rect 7686 6768 7704 6786
rect 7686 6786 7704 6804
rect 7704 2214 7722 2232
rect 7704 2232 7722 2250
rect 7704 2250 7722 2268
rect 7704 2268 7722 2286
rect 7704 2286 7722 2304
rect 7704 2304 7722 2322
rect 7704 2322 7722 2340
rect 7704 2340 7722 2358
rect 7704 2358 7722 2376
rect 7704 2376 7722 2394
rect 7704 2394 7722 2412
rect 7704 2412 7722 2430
rect 7704 2430 7722 2448
rect 7704 2448 7722 2466
rect 7704 2466 7722 2484
rect 7704 2484 7722 2502
rect 7704 2502 7722 2520
rect 7704 2520 7722 2538
rect 7704 2538 7722 2556
rect 7704 2556 7722 2574
rect 7704 2574 7722 2592
rect 7704 2592 7722 2610
rect 7704 2610 7722 2628
rect 7704 2628 7722 2646
rect 7704 2646 7722 2664
rect 7704 2664 7722 2682
rect 7704 2682 7722 2700
rect 7704 2700 7722 2718
rect 7704 2718 7722 2736
rect 7704 2736 7722 2754
rect 7704 2754 7722 2772
rect 7704 2772 7722 2790
rect 7704 2790 7722 2808
rect 7704 2808 7722 2826
rect 7704 2826 7722 2844
rect 7704 2844 7722 2862
rect 7704 2862 7722 2880
rect 7704 2880 7722 2898
rect 7704 2898 7722 2916
rect 7704 2916 7722 2934
rect 7704 2934 7722 2952
rect 7704 2952 7722 2970
rect 7704 2970 7722 2988
rect 7704 2988 7722 3006
rect 7704 3006 7722 3024
rect 7704 3024 7722 3042
rect 7704 3042 7722 3060
rect 7704 3060 7722 3078
rect 7704 3078 7722 3096
rect 7704 3096 7722 3114
rect 7704 3114 7722 3132
rect 7704 3132 7722 3150
rect 7704 3150 7722 3168
rect 7704 3168 7722 3186
rect 7704 3186 7722 3204
rect 7704 3204 7722 3222
rect 7704 3222 7722 3240
rect 7704 3240 7722 3258
rect 7704 3258 7722 3276
rect 7704 3276 7722 3294
rect 7704 4896 7722 4914
rect 7704 4914 7722 4932
rect 7704 4932 7722 4950
rect 7704 4950 7722 4968
rect 7704 4968 7722 4986
rect 7704 4986 7722 5004
rect 7704 5004 7722 5022
rect 7704 5022 7722 5040
rect 7704 5040 7722 5058
rect 7704 5058 7722 5076
rect 7704 5076 7722 5094
rect 7704 5094 7722 5112
rect 7704 5112 7722 5130
rect 7704 5130 7722 5148
rect 7704 5148 7722 5166
rect 7704 5166 7722 5184
rect 7704 5184 7722 5202
rect 7704 5202 7722 5220
rect 7704 5220 7722 5238
rect 7704 5238 7722 5256
rect 7704 5256 7722 5274
rect 7704 5274 7722 5292
rect 7704 5292 7722 5310
rect 7704 5310 7722 5328
rect 7704 5328 7722 5346
rect 7704 5346 7722 5364
rect 7704 5364 7722 5382
rect 7704 5382 7722 5400
rect 7704 5400 7722 5418
rect 7704 5418 7722 5436
rect 7704 5436 7722 5454
rect 7704 5454 7722 5472
rect 7704 5472 7722 5490
rect 7704 5490 7722 5508
rect 7704 5508 7722 5526
rect 7704 5526 7722 5544
rect 7704 5544 7722 5562
rect 7704 5562 7722 5580
rect 7704 5580 7722 5598
rect 7704 5598 7722 5616
rect 7704 5616 7722 5634
rect 7704 5634 7722 5652
rect 7704 5652 7722 5670
rect 7704 5670 7722 5688
rect 7704 5688 7722 5706
rect 7704 5706 7722 5724
rect 7704 5724 7722 5742
rect 7704 5742 7722 5760
rect 7704 5760 7722 5778
rect 7704 5778 7722 5796
rect 7704 5796 7722 5814
rect 7704 5814 7722 5832
rect 7704 5832 7722 5850
rect 7704 5850 7722 5868
rect 7704 5868 7722 5886
rect 7704 5886 7722 5904
rect 7704 5904 7722 5922
rect 7704 5922 7722 5940
rect 7704 5940 7722 5958
rect 7704 5958 7722 5976
rect 7704 5976 7722 5994
rect 7704 5994 7722 6012
rect 7704 6012 7722 6030
rect 7704 6030 7722 6048
rect 7704 6048 7722 6066
rect 7704 6066 7722 6084
rect 7704 6084 7722 6102
rect 7704 6102 7722 6120
rect 7704 6120 7722 6138
rect 7704 6138 7722 6156
rect 7704 6156 7722 6174
rect 7704 6174 7722 6192
rect 7704 6192 7722 6210
rect 7704 6210 7722 6228
rect 7704 6228 7722 6246
rect 7704 6246 7722 6264
rect 7704 6264 7722 6282
rect 7704 6282 7722 6300
rect 7704 6300 7722 6318
rect 7704 6318 7722 6336
rect 7704 6336 7722 6354
rect 7704 6354 7722 6372
rect 7704 6372 7722 6390
rect 7704 6390 7722 6408
rect 7704 6408 7722 6426
rect 7704 6426 7722 6444
rect 7704 6444 7722 6462
rect 7704 6462 7722 6480
rect 7704 6480 7722 6498
rect 7704 6498 7722 6516
rect 7704 6516 7722 6534
rect 7704 6534 7722 6552
rect 7704 6552 7722 6570
rect 7704 6570 7722 6588
rect 7704 6588 7722 6606
rect 7704 6606 7722 6624
rect 7704 6624 7722 6642
rect 7704 6642 7722 6660
rect 7704 6660 7722 6678
rect 7704 6678 7722 6696
rect 7704 6696 7722 6714
rect 7704 6714 7722 6732
rect 7704 6732 7722 6750
rect 7704 6750 7722 6768
rect 7704 6768 7722 6786
rect 7704 6786 7722 6804
rect 7722 2232 7740 2250
rect 7722 2250 7740 2268
rect 7722 2268 7740 2286
rect 7722 2286 7740 2304
rect 7722 2304 7740 2322
rect 7722 2322 7740 2340
rect 7722 2340 7740 2358
rect 7722 2358 7740 2376
rect 7722 2376 7740 2394
rect 7722 2394 7740 2412
rect 7722 2412 7740 2430
rect 7722 2430 7740 2448
rect 7722 2448 7740 2466
rect 7722 2466 7740 2484
rect 7722 2484 7740 2502
rect 7722 2502 7740 2520
rect 7722 2520 7740 2538
rect 7722 2538 7740 2556
rect 7722 2556 7740 2574
rect 7722 2574 7740 2592
rect 7722 2592 7740 2610
rect 7722 2610 7740 2628
rect 7722 2628 7740 2646
rect 7722 2646 7740 2664
rect 7722 2664 7740 2682
rect 7722 2682 7740 2700
rect 7722 2700 7740 2718
rect 7722 2718 7740 2736
rect 7722 2736 7740 2754
rect 7722 2754 7740 2772
rect 7722 2772 7740 2790
rect 7722 2790 7740 2808
rect 7722 2808 7740 2826
rect 7722 2826 7740 2844
rect 7722 2844 7740 2862
rect 7722 2862 7740 2880
rect 7722 2880 7740 2898
rect 7722 2898 7740 2916
rect 7722 2916 7740 2934
rect 7722 2934 7740 2952
rect 7722 2952 7740 2970
rect 7722 2970 7740 2988
rect 7722 2988 7740 3006
rect 7722 3006 7740 3024
rect 7722 3024 7740 3042
rect 7722 3042 7740 3060
rect 7722 3060 7740 3078
rect 7722 3078 7740 3096
rect 7722 3096 7740 3114
rect 7722 3114 7740 3132
rect 7722 3132 7740 3150
rect 7722 3150 7740 3168
rect 7722 3168 7740 3186
rect 7722 3186 7740 3204
rect 7722 3204 7740 3222
rect 7722 3222 7740 3240
rect 7722 3240 7740 3258
rect 7722 3258 7740 3276
rect 7722 3276 7740 3294
rect 7722 4914 7740 4932
rect 7722 4932 7740 4950
rect 7722 4950 7740 4968
rect 7722 4968 7740 4986
rect 7722 4986 7740 5004
rect 7722 5004 7740 5022
rect 7722 5022 7740 5040
rect 7722 5040 7740 5058
rect 7722 5058 7740 5076
rect 7722 5076 7740 5094
rect 7722 5094 7740 5112
rect 7722 5112 7740 5130
rect 7722 5130 7740 5148
rect 7722 5148 7740 5166
rect 7722 5166 7740 5184
rect 7722 5184 7740 5202
rect 7722 5202 7740 5220
rect 7722 5220 7740 5238
rect 7722 5238 7740 5256
rect 7722 5256 7740 5274
rect 7722 5274 7740 5292
rect 7722 5292 7740 5310
rect 7722 5310 7740 5328
rect 7722 5328 7740 5346
rect 7722 5346 7740 5364
rect 7722 5364 7740 5382
rect 7722 5382 7740 5400
rect 7722 5400 7740 5418
rect 7722 5418 7740 5436
rect 7722 5436 7740 5454
rect 7722 5454 7740 5472
rect 7722 5472 7740 5490
rect 7722 5490 7740 5508
rect 7722 5508 7740 5526
rect 7722 5526 7740 5544
rect 7722 5544 7740 5562
rect 7722 5562 7740 5580
rect 7722 5580 7740 5598
rect 7722 5598 7740 5616
rect 7722 5616 7740 5634
rect 7722 5634 7740 5652
rect 7722 5652 7740 5670
rect 7722 5670 7740 5688
rect 7722 5688 7740 5706
rect 7722 5706 7740 5724
rect 7722 5724 7740 5742
rect 7722 5742 7740 5760
rect 7722 5760 7740 5778
rect 7722 5778 7740 5796
rect 7722 5796 7740 5814
rect 7722 5814 7740 5832
rect 7722 5832 7740 5850
rect 7722 5850 7740 5868
rect 7722 5868 7740 5886
rect 7722 5886 7740 5904
rect 7722 5904 7740 5922
rect 7722 5922 7740 5940
rect 7722 5940 7740 5958
rect 7722 5958 7740 5976
rect 7722 5976 7740 5994
rect 7722 5994 7740 6012
rect 7722 6012 7740 6030
rect 7722 6030 7740 6048
rect 7722 6048 7740 6066
rect 7722 6066 7740 6084
rect 7722 6084 7740 6102
rect 7722 6102 7740 6120
rect 7722 6120 7740 6138
rect 7722 6138 7740 6156
rect 7722 6156 7740 6174
rect 7722 6174 7740 6192
rect 7722 6192 7740 6210
rect 7722 6210 7740 6228
rect 7722 6228 7740 6246
rect 7722 6246 7740 6264
rect 7722 6264 7740 6282
rect 7722 6282 7740 6300
rect 7722 6300 7740 6318
rect 7722 6318 7740 6336
rect 7722 6336 7740 6354
rect 7722 6354 7740 6372
rect 7722 6372 7740 6390
rect 7722 6390 7740 6408
rect 7722 6408 7740 6426
rect 7722 6426 7740 6444
rect 7722 6444 7740 6462
rect 7722 6462 7740 6480
rect 7722 6480 7740 6498
rect 7722 6498 7740 6516
rect 7722 6516 7740 6534
rect 7722 6534 7740 6552
rect 7722 6552 7740 6570
rect 7722 6570 7740 6588
rect 7722 6588 7740 6606
rect 7722 6606 7740 6624
rect 7722 6624 7740 6642
rect 7722 6642 7740 6660
rect 7722 6660 7740 6678
rect 7722 6678 7740 6696
rect 7722 6696 7740 6714
rect 7722 6714 7740 6732
rect 7722 6732 7740 6750
rect 7722 6750 7740 6768
rect 7722 6768 7740 6786
rect 7722 6786 7740 6804
rect 7722 6804 7740 6822
rect 7740 2232 7758 2250
rect 7740 2250 7758 2268
rect 7740 2268 7758 2286
rect 7740 2286 7758 2304
rect 7740 2304 7758 2322
rect 7740 2322 7758 2340
rect 7740 2340 7758 2358
rect 7740 2358 7758 2376
rect 7740 2376 7758 2394
rect 7740 2394 7758 2412
rect 7740 2412 7758 2430
rect 7740 2430 7758 2448
rect 7740 2448 7758 2466
rect 7740 2466 7758 2484
rect 7740 2484 7758 2502
rect 7740 2502 7758 2520
rect 7740 2520 7758 2538
rect 7740 2538 7758 2556
rect 7740 2556 7758 2574
rect 7740 2574 7758 2592
rect 7740 2592 7758 2610
rect 7740 2610 7758 2628
rect 7740 2628 7758 2646
rect 7740 2646 7758 2664
rect 7740 2664 7758 2682
rect 7740 2682 7758 2700
rect 7740 2700 7758 2718
rect 7740 2718 7758 2736
rect 7740 2736 7758 2754
rect 7740 2754 7758 2772
rect 7740 2772 7758 2790
rect 7740 2790 7758 2808
rect 7740 2808 7758 2826
rect 7740 2826 7758 2844
rect 7740 2844 7758 2862
rect 7740 2862 7758 2880
rect 7740 2880 7758 2898
rect 7740 2898 7758 2916
rect 7740 2916 7758 2934
rect 7740 2934 7758 2952
rect 7740 2952 7758 2970
rect 7740 2970 7758 2988
rect 7740 2988 7758 3006
rect 7740 3006 7758 3024
rect 7740 3024 7758 3042
rect 7740 3042 7758 3060
rect 7740 3060 7758 3078
rect 7740 3078 7758 3096
rect 7740 3096 7758 3114
rect 7740 3114 7758 3132
rect 7740 3132 7758 3150
rect 7740 3150 7758 3168
rect 7740 3168 7758 3186
rect 7740 3186 7758 3204
rect 7740 3204 7758 3222
rect 7740 3222 7758 3240
rect 7740 3240 7758 3258
rect 7740 3258 7758 3276
rect 7740 3276 7758 3294
rect 7740 4932 7758 4950
rect 7740 4950 7758 4968
rect 7740 4968 7758 4986
rect 7740 4986 7758 5004
rect 7740 5004 7758 5022
rect 7740 5022 7758 5040
rect 7740 5040 7758 5058
rect 7740 5058 7758 5076
rect 7740 5076 7758 5094
rect 7740 5094 7758 5112
rect 7740 5112 7758 5130
rect 7740 5130 7758 5148
rect 7740 5148 7758 5166
rect 7740 5166 7758 5184
rect 7740 5184 7758 5202
rect 7740 5202 7758 5220
rect 7740 5220 7758 5238
rect 7740 5238 7758 5256
rect 7740 5256 7758 5274
rect 7740 5274 7758 5292
rect 7740 5292 7758 5310
rect 7740 5310 7758 5328
rect 7740 5328 7758 5346
rect 7740 5346 7758 5364
rect 7740 5364 7758 5382
rect 7740 5382 7758 5400
rect 7740 5400 7758 5418
rect 7740 5418 7758 5436
rect 7740 5436 7758 5454
rect 7740 5454 7758 5472
rect 7740 5472 7758 5490
rect 7740 5490 7758 5508
rect 7740 5508 7758 5526
rect 7740 5526 7758 5544
rect 7740 5544 7758 5562
rect 7740 5562 7758 5580
rect 7740 5580 7758 5598
rect 7740 5598 7758 5616
rect 7740 5616 7758 5634
rect 7740 5634 7758 5652
rect 7740 5652 7758 5670
rect 7740 5670 7758 5688
rect 7740 5688 7758 5706
rect 7740 5706 7758 5724
rect 7740 5724 7758 5742
rect 7740 5742 7758 5760
rect 7740 5760 7758 5778
rect 7740 5778 7758 5796
rect 7740 5796 7758 5814
rect 7740 5814 7758 5832
rect 7740 5832 7758 5850
rect 7740 5850 7758 5868
rect 7740 5868 7758 5886
rect 7740 5886 7758 5904
rect 7740 5904 7758 5922
rect 7740 5922 7758 5940
rect 7740 5940 7758 5958
rect 7740 5958 7758 5976
rect 7740 5976 7758 5994
rect 7740 5994 7758 6012
rect 7740 6012 7758 6030
rect 7740 6030 7758 6048
rect 7740 6048 7758 6066
rect 7740 6066 7758 6084
rect 7740 6084 7758 6102
rect 7740 6102 7758 6120
rect 7740 6120 7758 6138
rect 7740 6138 7758 6156
rect 7740 6156 7758 6174
rect 7740 6174 7758 6192
rect 7740 6192 7758 6210
rect 7740 6210 7758 6228
rect 7740 6228 7758 6246
rect 7740 6246 7758 6264
rect 7740 6264 7758 6282
rect 7740 6282 7758 6300
rect 7740 6300 7758 6318
rect 7740 6318 7758 6336
rect 7740 6336 7758 6354
rect 7740 6354 7758 6372
rect 7740 6372 7758 6390
rect 7740 6390 7758 6408
rect 7740 6408 7758 6426
rect 7740 6426 7758 6444
rect 7740 6444 7758 6462
rect 7740 6462 7758 6480
rect 7740 6480 7758 6498
rect 7740 6498 7758 6516
rect 7740 6516 7758 6534
rect 7740 6534 7758 6552
rect 7740 6552 7758 6570
rect 7740 6570 7758 6588
rect 7740 6588 7758 6606
rect 7740 6606 7758 6624
rect 7740 6624 7758 6642
rect 7740 6642 7758 6660
rect 7740 6660 7758 6678
rect 7740 6678 7758 6696
rect 7740 6696 7758 6714
rect 7740 6714 7758 6732
rect 7740 6732 7758 6750
rect 7740 6750 7758 6768
rect 7740 6768 7758 6786
rect 7740 6786 7758 6804
rect 7740 6804 7758 6822
rect 7740 6822 7758 6840
rect 7758 2250 7776 2268
rect 7758 2268 7776 2286
rect 7758 2286 7776 2304
rect 7758 2304 7776 2322
rect 7758 2322 7776 2340
rect 7758 2340 7776 2358
rect 7758 2358 7776 2376
rect 7758 2376 7776 2394
rect 7758 2394 7776 2412
rect 7758 2412 7776 2430
rect 7758 2430 7776 2448
rect 7758 2448 7776 2466
rect 7758 2466 7776 2484
rect 7758 2484 7776 2502
rect 7758 2502 7776 2520
rect 7758 2520 7776 2538
rect 7758 2538 7776 2556
rect 7758 2556 7776 2574
rect 7758 2574 7776 2592
rect 7758 2592 7776 2610
rect 7758 2610 7776 2628
rect 7758 2628 7776 2646
rect 7758 2646 7776 2664
rect 7758 2664 7776 2682
rect 7758 2682 7776 2700
rect 7758 2700 7776 2718
rect 7758 2718 7776 2736
rect 7758 2736 7776 2754
rect 7758 2754 7776 2772
rect 7758 2772 7776 2790
rect 7758 2790 7776 2808
rect 7758 2808 7776 2826
rect 7758 2826 7776 2844
rect 7758 2844 7776 2862
rect 7758 2862 7776 2880
rect 7758 2880 7776 2898
rect 7758 2898 7776 2916
rect 7758 2916 7776 2934
rect 7758 2934 7776 2952
rect 7758 2952 7776 2970
rect 7758 2970 7776 2988
rect 7758 2988 7776 3006
rect 7758 3006 7776 3024
rect 7758 3024 7776 3042
rect 7758 3042 7776 3060
rect 7758 3060 7776 3078
rect 7758 3078 7776 3096
rect 7758 3096 7776 3114
rect 7758 3114 7776 3132
rect 7758 3132 7776 3150
rect 7758 3150 7776 3168
rect 7758 3168 7776 3186
rect 7758 3186 7776 3204
rect 7758 3204 7776 3222
rect 7758 3222 7776 3240
rect 7758 3240 7776 3258
rect 7758 3258 7776 3276
rect 7758 3276 7776 3294
rect 7758 4968 7776 4986
rect 7758 4986 7776 5004
rect 7758 5004 7776 5022
rect 7758 5022 7776 5040
rect 7758 5040 7776 5058
rect 7758 5058 7776 5076
rect 7758 5076 7776 5094
rect 7758 5094 7776 5112
rect 7758 5112 7776 5130
rect 7758 5130 7776 5148
rect 7758 5148 7776 5166
rect 7758 5166 7776 5184
rect 7758 5184 7776 5202
rect 7758 5202 7776 5220
rect 7758 5220 7776 5238
rect 7758 5238 7776 5256
rect 7758 5256 7776 5274
rect 7758 5274 7776 5292
rect 7758 5292 7776 5310
rect 7758 5310 7776 5328
rect 7758 5328 7776 5346
rect 7758 5346 7776 5364
rect 7758 5364 7776 5382
rect 7758 5382 7776 5400
rect 7758 5400 7776 5418
rect 7758 5418 7776 5436
rect 7758 5436 7776 5454
rect 7758 5454 7776 5472
rect 7758 5472 7776 5490
rect 7758 5490 7776 5508
rect 7758 5508 7776 5526
rect 7758 5526 7776 5544
rect 7758 5544 7776 5562
rect 7758 5562 7776 5580
rect 7758 5580 7776 5598
rect 7758 5598 7776 5616
rect 7758 5616 7776 5634
rect 7758 5634 7776 5652
rect 7758 5652 7776 5670
rect 7758 5670 7776 5688
rect 7758 5688 7776 5706
rect 7758 5706 7776 5724
rect 7758 5724 7776 5742
rect 7758 5742 7776 5760
rect 7758 5760 7776 5778
rect 7758 5778 7776 5796
rect 7758 5796 7776 5814
rect 7758 5814 7776 5832
rect 7758 5832 7776 5850
rect 7758 5850 7776 5868
rect 7758 5868 7776 5886
rect 7758 5886 7776 5904
rect 7758 5904 7776 5922
rect 7758 5922 7776 5940
rect 7758 5940 7776 5958
rect 7758 5958 7776 5976
rect 7758 5976 7776 5994
rect 7758 5994 7776 6012
rect 7758 6012 7776 6030
rect 7758 6030 7776 6048
rect 7758 6048 7776 6066
rect 7758 6066 7776 6084
rect 7758 6084 7776 6102
rect 7758 6102 7776 6120
rect 7758 6120 7776 6138
rect 7758 6138 7776 6156
rect 7758 6156 7776 6174
rect 7758 6174 7776 6192
rect 7758 6192 7776 6210
rect 7758 6210 7776 6228
rect 7758 6228 7776 6246
rect 7758 6246 7776 6264
rect 7758 6264 7776 6282
rect 7758 6282 7776 6300
rect 7758 6300 7776 6318
rect 7758 6318 7776 6336
rect 7758 6336 7776 6354
rect 7758 6354 7776 6372
rect 7758 6372 7776 6390
rect 7758 6390 7776 6408
rect 7758 6408 7776 6426
rect 7758 6426 7776 6444
rect 7758 6444 7776 6462
rect 7758 6462 7776 6480
rect 7758 6480 7776 6498
rect 7758 6498 7776 6516
rect 7758 6516 7776 6534
rect 7758 6534 7776 6552
rect 7758 6552 7776 6570
rect 7758 6570 7776 6588
rect 7758 6588 7776 6606
rect 7758 6606 7776 6624
rect 7758 6624 7776 6642
rect 7758 6642 7776 6660
rect 7758 6660 7776 6678
rect 7758 6678 7776 6696
rect 7758 6696 7776 6714
rect 7758 6714 7776 6732
rect 7758 6732 7776 6750
rect 7758 6750 7776 6768
rect 7758 6768 7776 6786
rect 7758 6786 7776 6804
rect 7758 6804 7776 6822
rect 7758 6822 7776 6840
rect 7758 6840 7776 6858
rect 7776 2268 7794 2286
rect 7776 2286 7794 2304
rect 7776 2304 7794 2322
rect 7776 2322 7794 2340
rect 7776 2340 7794 2358
rect 7776 2358 7794 2376
rect 7776 2376 7794 2394
rect 7776 2394 7794 2412
rect 7776 2412 7794 2430
rect 7776 2430 7794 2448
rect 7776 2448 7794 2466
rect 7776 2466 7794 2484
rect 7776 2484 7794 2502
rect 7776 2502 7794 2520
rect 7776 2520 7794 2538
rect 7776 2538 7794 2556
rect 7776 2556 7794 2574
rect 7776 2574 7794 2592
rect 7776 2592 7794 2610
rect 7776 2610 7794 2628
rect 7776 2628 7794 2646
rect 7776 2646 7794 2664
rect 7776 2664 7794 2682
rect 7776 2682 7794 2700
rect 7776 2700 7794 2718
rect 7776 2718 7794 2736
rect 7776 2736 7794 2754
rect 7776 2754 7794 2772
rect 7776 2772 7794 2790
rect 7776 2790 7794 2808
rect 7776 2808 7794 2826
rect 7776 2826 7794 2844
rect 7776 2844 7794 2862
rect 7776 2862 7794 2880
rect 7776 2880 7794 2898
rect 7776 2898 7794 2916
rect 7776 2916 7794 2934
rect 7776 2934 7794 2952
rect 7776 2952 7794 2970
rect 7776 2970 7794 2988
rect 7776 2988 7794 3006
rect 7776 3006 7794 3024
rect 7776 3024 7794 3042
rect 7776 3042 7794 3060
rect 7776 3060 7794 3078
rect 7776 3078 7794 3096
rect 7776 3096 7794 3114
rect 7776 3114 7794 3132
rect 7776 3132 7794 3150
rect 7776 3150 7794 3168
rect 7776 3168 7794 3186
rect 7776 3186 7794 3204
rect 7776 3204 7794 3222
rect 7776 3222 7794 3240
rect 7776 3240 7794 3258
rect 7776 3258 7794 3276
rect 7776 3276 7794 3294
rect 7776 3294 7794 3312
rect 7776 4986 7794 5004
rect 7776 5004 7794 5022
rect 7776 5022 7794 5040
rect 7776 5040 7794 5058
rect 7776 5058 7794 5076
rect 7776 5076 7794 5094
rect 7776 5094 7794 5112
rect 7776 5112 7794 5130
rect 7776 5130 7794 5148
rect 7776 5148 7794 5166
rect 7776 5166 7794 5184
rect 7776 5184 7794 5202
rect 7776 5202 7794 5220
rect 7776 5220 7794 5238
rect 7776 5238 7794 5256
rect 7776 5256 7794 5274
rect 7776 5274 7794 5292
rect 7776 5292 7794 5310
rect 7776 5310 7794 5328
rect 7776 5328 7794 5346
rect 7776 5346 7794 5364
rect 7776 5364 7794 5382
rect 7776 5382 7794 5400
rect 7776 5400 7794 5418
rect 7776 5418 7794 5436
rect 7776 5436 7794 5454
rect 7776 5454 7794 5472
rect 7776 5472 7794 5490
rect 7776 5490 7794 5508
rect 7776 5508 7794 5526
rect 7776 5526 7794 5544
rect 7776 5544 7794 5562
rect 7776 5562 7794 5580
rect 7776 5580 7794 5598
rect 7776 5598 7794 5616
rect 7776 5616 7794 5634
rect 7776 5634 7794 5652
rect 7776 5652 7794 5670
rect 7776 5670 7794 5688
rect 7776 5688 7794 5706
rect 7776 5706 7794 5724
rect 7776 5724 7794 5742
rect 7776 5742 7794 5760
rect 7776 5760 7794 5778
rect 7776 5778 7794 5796
rect 7776 5796 7794 5814
rect 7776 5814 7794 5832
rect 7776 5832 7794 5850
rect 7776 5850 7794 5868
rect 7776 5868 7794 5886
rect 7776 5886 7794 5904
rect 7776 5904 7794 5922
rect 7776 5922 7794 5940
rect 7776 5940 7794 5958
rect 7776 5958 7794 5976
rect 7776 5976 7794 5994
rect 7776 5994 7794 6012
rect 7776 6012 7794 6030
rect 7776 6030 7794 6048
rect 7776 6048 7794 6066
rect 7776 6066 7794 6084
rect 7776 6084 7794 6102
rect 7776 6102 7794 6120
rect 7776 6120 7794 6138
rect 7776 6138 7794 6156
rect 7776 6156 7794 6174
rect 7776 6174 7794 6192
rect 7776 6192 7794 6210
rect 7776 6210 7794 6228
rect 7776 6228 7794 6246
rect 7776 6246 7794 6264
rect 7776 6264 7794 6282
rect 7776 6282 7794 6300
rect 7776 6300 7794 6318
rect 7776 6318 7794 6336
rect 7776 6336 7794 6354
rect 7776 6354 7794 6372
rect 7776 6372 7794 6390
rect 7776 6390 7794 6408
rect 7776 6408 7794 6426
rect 7776 6426 7794 6444
rect 7776 6444 7794 6462
rect 7776 6462 7794 6480
rect 7776 6480 7794 6498
rect 7776 6498 7794 6516
rect 7776 6516 7794 6534
rect 7776 6534 7794 6552
rect 7776 6552 7794 6570
rect 7776 6570 7794 6588
rect 7776 6588 7794 6606
rect 7776 6606 7794 6624
rect 7776 6624 7794 6642
rect 7776 6642 7794 6660
rect 7776 6660 7794 6678
rect 7776 6678 7794 6696
rect 7776 6696 7794 6714
rect 7776 6714 7794 6732
rect 7776 6732 7794 6750
rect 7776 6750 7794 6768
rect 7776 6768 7794 6786
rect 7776 6786 7794 6804
rect 7776 6804 7794 6822
rect 7776 6822 7794 6840
rect 7776 6840 7794 6858
rect 7794 2268 7812 2286
rect 7794 2286 7812 2304
rect 7794 2304 7812 2322
rect 7794 2322 7812 2340
rect 7794 2340 7812 2358
rect 7794 2358 7812 2376
rect 7794 2376 7812 2394
rect 7794 2394 7812 2412
rect 7794 2412 7812 2430
rect 7794 2430 7812 2448
rect 7794 2448 7812 2466
rect 7794 2466 7812 2484
rect 7794 2484 7812 2502
rect 7794 2502 7812 2520
rect 7794 2520 7812 2538
rect 7794 2538 7812 2556
rect 7794 2556 7812 2574
rect 7794 2574 7812 2592
rect 7794 2592 7812 2610
rect 7794 2610 7812 2628
rect 7794 2628 7812 2646
rect 7794 2646 7812 2664
rect 7794 2664 7812 2682
rect 7794 2682 7812 2700
rect 7794 2700 7812 2718
rect 7794 2718 7812 2736
rect 7794 2736 7812 2754
rect 7794 2754 7812 2772
rect 7794 2772 7812 2790
rect 7794 2790 7812 2808
rect 7794 2808 7812 2826
rect 7794 2826 7812 2844
rect 7794 2844 7812 2862
rect 7794 2862 7812 2880
rect 7794 2880 7812 2898
rect 7794 2898 7812 2916
rect 7794 2916 7812 2934
rect 7794 2934 7812 2952
rect 7794 2952 7812 2970
rect 7794 2970 7812 2988
rect 7794 2988 7812 3006
rect 7794 3006 7812 3024
rect 7794 3024 7812 3042
rect 7794 3042 7812 3060
rect 7794 3060 7812 3078
rect 7794 3078 7812 3096
rect 7794 3096 7812 3114
rect 7794 3114 7812 3132
rect 7794 3132 7812 3150
rect 7794 3150 7812 3168
rect 7794 3168 7812 3186
rect 7794 3186 7812 3204
rect 7794 3204 7812 3222
rect 7794 3222 7812 3240
rect 7794 3240 7812 3258
rect 7794 3258 7812 3276
rect 7794 3276 7812 3294
rect 7794 3294 7812 3312
rect 7794 5004 7812 5022
rect 7794 5022 7812 5040
rect 7794 5040 7812 5058
rect 7794 5058 7812 5076
rect 7794 5076 7812 5094
rect 7794 5094 7812 5112
rect 7794 5112 7812 5130
rect 7794 5130 7812 5148
rect 7794 5148 7812 5166
rect 7794 5166 7812 5184
rect 7794 5184 7812 5202
rect 7794 5202 7812 5220
rect 7794 5220 7812 5238
rect 7794 5238 7812 5256
rect 7794 5256 7812 5274
rect 7794 5274 7812 5292
rect 7794 5292 7812 5310
rect 7794 5310 7812 5328
rect 7794 5328 7812 5346
rect 7794 5346 7812 5364
rect 7794 5364 7812 5382
rect 7794 5382 7812 5400
rect 7794 5400 7812 5418
rect 7794 5418 7812 5436
rect 7794 5436 7812 5454
rect 7794 5454 7812 5472
rect 7794 5472 7812 5490
rect 7794 5490 7812 5508
rect 7794 5508 7812 5526
rect 7794 5526 7812 5544
rect 7794 5544 7812 5562
rect 7794 5562 7812 5580
rect 7794 5580 7812 5598
rect 7794 5598 7812 5616
rect 7794 5616 7812 5634
rect 7794 5634 7812 5652
rect 7794 5652 7812 5670
rect 7794 5670 7812 5688
rect 7794 5688 7812 5706
rect 7794 5706 7812 5724
rect 7794 5724 7812 5742
rect 7794 5742 7812 5760
rect 7794 5760 7812 5778
rect 7794 5778 7812 5796
rect 7794 5796 7812 5814
rect 7794 5814 7812 5832
rect 7794 5832 7812 5850
rect 7794 5850 7812 5868
rect 7794 5868 7812 5886
rect 7794 5886 7812 5904
rect 7794 5904 7812 5922
rect 7794 5922 7812 5940
rect 7794 5940 7812 5958
rect 7794 5958 7812 5976
rect 7794 5976 7812 5994
rect 7794 5994 7812 6012
rect 7794 6012 7812 6030
rect 7794 6030 7812 6048
rect 7794 6048 7812 6066
rect 7794 6066 7812 6084
rect 7794 6084 7812 6102
rect 7794 6102 7812 6120
rect 7794 6120 7812 6138
rect 7794 6138 7812 6156
rect 7794 6156 7812 6174
rect 7794 6174 7812 6192
rect 7794 6192 7812 6210
rect 7794 6210 7812 6228
rect 7794 6228 7812 6246
rect 7794 6246 7812 6264
rect 7794 6264 7812 6282
rect 7794 6282 7812 6300
rect 7794 6300 7812 6318
rect 7794 6318 7812 6336
rect 7794 6336 7812 6354
rect 7794 6354 7812 6372
rect 7794 6372 7812 6390
rect 7794 6390 7812 6408
rect 7794 6408 7812 6426
rect 7794 6426 7812 6444
rect 7794 6444 7812 6462
rect 7794 6462 7812 6480
rect 7794 6480 7812 6498
rect 7794 6498 7812 6516
rect 7794 6516 7812 6534
rect 7794 6534 7812 6552
rect 7794 6552 7812 6570
rect 7794 6570 7812 6588
rect 7794 6588 7812 6606
rect 7794 6606 7812 6624
rect 7794 6624 7812 6642
rect 7794 6642 7812 6660
rect 7794 6660 7812 6678
rect 7794 6678 7812 6696
rect 7794 6696 7812 6714
rect 7794 6714 7812 6732
rect 7794 6732 7812 6750
rect 7794 6750 7812 6768
rect 7794 6768 7812 6786
rect 7794 6786 7812 6804
rect 7794 6804 7812 6822
rect 7794 6822 7812 6840
rect 7794 6840 7812 6858
rect 7794 6858 7812 6876
rect 7812 2286 7830 2304
rect 7812 2304 7830 2322
rect 7812 2322 7830 2340
rect 7812 2340 7830 2358
rect 7812 2358 7830 2376
rect 7812 2376 7830 2394
rect 7812 2394 7830 2412
rect 7812 2412 7830 2430
rect 7812 2430 7830 2448
rect 7812 2448 7830 2466
rect 7812 2466 7830 2484
rect 7812 2484 7830 2502
rect 7812 2502 7830 2520
rect 7812 2520 7830 2538
rect 7812 2538 7830 2556
rect 7812 2556 7830 2574
rect 7812 2574 7830 2592
rect 7812 2592 7830 2610
rect 7812 2610 7830 2628
rect 7812 2628 7830 2646
rect 7812 2646 7830 2664
rect 7812 2664 7830 2682
rect 7812 2682 7830 2700
rect 7812 2700 7830 2718
rect 7812 2718 7830 2736
rect 7812 2736 7830 2754
rect 7812 2754 7830 2772
rect 7812 2772 7830 2790
rect 7812 2790 7830 2808
rect 7812 2808 7830 2826
rect 7812 2826 7830 2844
rect 7812 2844 7830 2862
rect 7812 2862 7830 2880
rect 7812 2880 7830 2898
rect 7812 2898 7830 2916
rect 7812 2916 7830 2934
rect 7812 2934 7830 2952
rect 7812 2952 7830 2970
rect 7812 2970 7830 2988
rect 7812 2988 7830 3006
rect 7812 3006 7830 3024
rect 7812 3024 7830 3042
rect 7812 3042 7830 3060
rect 7812 3060 7830 3078
rect 7812 3078 7830 3096
rect 7812 3096 7830 3114
rect 7812 3114 7830 3132
rect 7812 3132 7830 3150
rect 7812 3150 7830 3168
rect 7812 3168 7830 3186
rect 7812 3186 7830 3204
rect 7812 3204 7830 3222
rect 7812 3222 7830 3240
rect 7812 3240 7830 3258
rect 7812 3258 7830 3276
rect 7812 3276 7830 3294
rect 7812 3294 7830 3312
rect 7812 5022 7830 5040
rect 7812 5040 7830 5058
rect 7812 5058 7830 5076
rect 7812 5076 7830 5094
rect 7812 5094 7830 5112
rect 7812 5112 7830 5130
rect 7812 5130 7830 5148
rect 7812 5148 7830 5166
rect 7812 5166 7830 5184
rect 7812 5184 7830 5202
rect 7812 5202 7830 5220
rect 7812 5220 7830 5238
rect 7812 5238 7830 5256
rect 7812 5256 7830 5274
rect 7812 5274 7830 5292
rect 7812 5292 7830 5310
rect 7812 5310 7830 5328
rect 7812 5328 7830 5346
rect 7812 5346 7830 5364
rect 7812 5364 7830 5382
rect 7812 5382 7830 5400
rect 7812 5400 7830 5418
rect 7812 5418 7830 5436
rect 7812 5436 7830 5454
rect 7812 5454 7830 5472
rect 7812 5472 7830 5490
rect 7812 5490 7830 5508
rect 7812 5508 7830 5526
rect 7812 5526 7830 5544
rect 7812 5544 7830 5562
rect 7812 5562 7830 5580
rect 7812 5580 7830 5598
rect 7812 5598 7830 5616
rect 7812 5616 7830 5634
rect 7812 5634 7830 5652
rect 7812 5652 7830 5670
rect 7812 5670 7830 5688
rect 7812 5688 7830 5706
rect 7812 5706 7830 5724
rect 7812 5724 7830 5742
rect 7812 5742 7830 5760
rect 7812 5760 7830 5778
rect 7812 5778 7830 5796
rect 7812 5796 7830 5814
rect 7812 5814 7830 5832
rect 7812 5832 7830 5850
rect 7812 5850 7830 5868
rect 7812 5868 7830 5886
rect 7812 5886 7830 5904
rect 7812 5904 7830 5922
rect 7812 5922 7830 5940
rect 7812 5940 7830 5958
rect 7812 5958 7830 5976
rect 7812 5976 7830 5994
rect 7812 5994 7830 6012
rect 7812 6012 7830 6030
rect 7812 6030 7830 6048
rect 7812 6048 7830 6066
rect 7812 6066 7830 6084
rect 7812 6084 7830 6102
rect 7812 6102 7830 6120
rect 7812 6120 7830 6138
rect 7812 6138 7830 6156
rect 7812 6156 7830 6174
rect 7812 6174 7830 6192
rect 7812 6192 7830 6210
rect 7812 6210 7830 6228
rect 7812 6228 7830 6246
rect 7812 6246 7830 6264
rect 7812 6264 7830 6282
rect 7812 6282 7830 6300
rect 7812 6300 7830 6318
rect 7812 6318 7830 6336
rect 7812 6336 7830 6354
rect 7812 6354 7830 6372
rect 7812 6372 7830 6390
rect 7812 6390 7830 6408
rect 7812 6408 7830 6426
rect 7812 6426 7830 6444
rect 7812 6444 7830 6462
rect 7812 6462 7830 6480
rect 7812 6480 7830 6498
rect 7812 6498 7830 6516
rect 7812 6516 7830 6534
rect 7812 6534 7830 6552
rect 7812 6552 7830 6570
rect 7812 6570 7830 6588
rect 7812 6588 7830 6606
rect 7812 6606 7830 6624
rect 7812 6624 7830 6642
rect 7812 6642 7830 6660
rect 7812 6660 7830 6678
rect 7812 6678 7830 6696
rect 7812 6696 7830 6714
rect 7812 6714 7830 6732
rect 7812 6732 7830 6750
rect 7812 6750 7830 6768
rect 7812 6768 7830 6786
rect 7812 6786 7830 6804
rect 7812 6804 7830 6822
rect 7812 6822 7830 6840
rect 7812 6840 7830 6858
rect 7812 6858 7830 6876
rect 7812 6876 7830 6894
rect 7830 2304 7848 2322
rect 7830 2322 7848 2340
rect 7830 2340 7848 2358
rect 7830 2358 7848 2376
rect 7830 2376 7848 2394
rect 7830 2394 7848 2412
rect 7830 2412 7848 2430
rect 7830 2430 7848 2448
rect 7830 2448 7848 2466
rect 7830 2466 7848 2484
rect 7830 2484 7848 2502
rect 7830 2502 7848 2520
rect 7830 2520 7848 2538
rect 7830 2538 7848 2556
rect 7830 2556 7848 2574
rect 7830 2574 7848 2592
rect 7830 2592 7848 2610
rect 7830 2610 7848 2628
rect 7830 2628 7848 2646
rect 7830 2646 7848 2664
rect 7830 2664 7848 2682
rect 7830 2682 7848 2700
rect 7830 2700 7848 2718
rect 7830 2718 7848 2736
rect 7830 2736 7848 2754
rect 7830 2754 7848 2772
rect 7830 2772 7848 2790
rect 7830 2790 7848 2808
rect 7830 2808 7848 2826
rect 7830 2826 7848 2844
rect 7830 2844 7848 2862
rect 7830 2862 7848 2880
rect 7830 2880 7848 2898
rect 7830 2898 7848 2916
rect 7830 2916 7848 2934
rect 7830 2934 7848 2952
rect 7830 2952 7848 2970
rect 7830 2970 7848 2988
rect 7830 2988 7848 3006
rect 7830 3006 7848 3024
rect 7830 3024 7848 3042
rect 7830 3042 7848 3060
rect 7830 3060 7848 3078
rect 7830 3078 7848 3096
rect 7830 3096 7848 3114
rect 7830 3114 7848 3132
rect 7830 3132 7848 3150
rect 7830 3150 7848 3168
rect 7830 3168 7848 3186
rect 7830 3186 7848 3204
rect 7830 3204 7848 3222
rect 7830 3222 7848 3240
rect 7830 3240 7848 3258
rect 7830 3258 7848 3276
rect 7830 3276 7848 3294
rect 7830 3294 7848 3312
rect 7830 3312 7848 3330
rect 7830 5058 7848 5076
rect 7830 5076 7848 5094
rect 7830 5094 7848 5112
rect 7830 5112 7848 5130
rect 7830 5130 7848 5148
rect 7830 5148 7848 5166
rect 7830 5166 7848 5184
rect 7830 5184 7848 5202
rect 7830 5202 7848 5220
rect 7830 5220 7848 5238
rect 7830 5238 7848 5256
rect 7830 5256 7848 5274
rect 7830 5274 7848 5292
rect 7830 5292 7848 5310
rect 7830 5310 7848 5328
rect 7830 5328 7848 5346
rect 7830 5346 7848 5364
rect 7830 5364 7848 5382
rect 7830 5382 7848 5400
rect 7830 5400 7848 5418
rect 7830 5418 7848 5436
rect 7830 5436 7848 5454
rect 7830 5454 7848 5472
rect 7830 5472 7848 5490
rect 7830 5490 7848 5508
rect 7830 5508 7848 5526
rect 7830 5526 7848 5544
rect 7830 5544 7848 5562
rect 7830 5562 7848 5580
rect 7830 5580 7848 5598
rect 7830 5598 7848 5616
rect 7830 5616 7848 5634
rect 7830 5634 7848 5652
rect 7830 5652 7848 5670
rect 7830 5670 7848 5688
rect 7830 5688 7848 5706
rect 7830 5706 7848 5724
rect 7830 5724 7848 5742
rect 7830 5742 7848 5760
rect 7830 5760 7848 5778
rect 7830 5778 7848 5796
rect 7830 5796 7848 5814
rect 7830 5814 7848 5832
rect 7830 5832 7848 5850
rect 7830 5850 7848 5868
rect 7830 5868 7848 5886
rect 7830 5886 7848 5904
rect 7830 5904 7848 5922
rect 7830 5922 7848 5940
rect 7830 5940 7848 5958
rect 7830 5958 7848 5976
rect 7830 5976 7848 5994
rect 7830 5994 7848 6012
rect 7830 6012 7848 6030
rect 7830 6030 7848 6048
rect 7830 6048 7848 6066
rect 7830 6066 7848 6084
rect 7830 6084 7848 6102
rect 7830 6102 7848 6120
rect 7830 6120 7848 6138
rect 7830 6138 7848 6156
rect 7830 6156 7848 6174
rect 7830 6174 7848 6192
rect 7830 6192 7848 6210
rect 7830 6210 7848 6228
rect 7830 6228 7848 6246
rect 7830 6246 7848 6264
rect 7830 6264 7848 6282
rect 7830 6282 7848 6300
rect 7830 6300 7848 6318
rect 7830 6318 7848 6336
rect 7830 6336 7848 6354
rect 7830 6354 7848 6372
rect 7830 6372 7848 6390
rect 7830 6390 7848 6408
rect 7830 6408 7848 6426
rect 7830 6426 7848 6444
rect 7830 6444 7848 6462
rect 7830 6462 7848 6480
rect 7830 6480 7848 6498
rect 7830 6498 7848 6516
rect 7830 6516 7848 6534
rect 7830 6534 7848 6552
rect 7830 6552 7848 6570
rect 7830 6570 7848 6588
rect 7830 6588 7848 6606
rect 7830 6606 7848 6624
rect 7830 6624 7848 6642
rect 7830 6642 7848 6660
rect 7830 6660 7848 6678
rect 7830 6678 7848 6696
rect 7830 6696 7848 6714
rect 7830 6714 7848 6732
rect 7830 6732 7848 6750
rect 7830 6750 7848 6768
rect 7830 6768 7848 6786
rect 7830 6786 7848 6804
rect 7830 6804 7848 6822
rect 7830 6822 7848 6840
rect 7830 6840 7848 6858
rect 7830 6858 7848 6876
rect 7830 6876 7848 6894
rect 7830 6894 7848 6912
rect 7848 2304 7866 2322
rect 7848 2322 7866 2340
rect 7848 2340 7866 2358
rect 7848 2358 7866 2376
rect 7848 2376 7866 2394
rect 7848 2394 7866 2412
rect 7848 2412 7866 2430
rect 7848 2430 7866 2448
rect 7848 2448 7866 2466
rect 7848 2466 7866 2484
rect 7848 2484 7866 2502
rect 7848 2502 7866 2520
rect 7848 2520 7866 2538
rect 7848 2538 7866 2556
rect 7848 2556 7866 2574
rect 7848 2574 7866 2592
rect 7848 2592 7866 2610
rect 7848 2610 7866 2628
rect 7848 2628 7866 2646
rect 7848 2646 7866 2664
rect 7848 2664 7866 2682
rect 7848 2682 7866 2700
rect 7848 2700 7866 2718
rect 7848 2718 7866 2736
rect 7848 2736 7866 2754
rect 7848 2754 7866 2772
rect 7848 2772 7866 2790
rect 7848 2790 7866 2808
rect 7848 2808 7866 2826
rect 7848 2826 7866 2844
rect 7848 2844 7866 2862
rect 7848 2862 7866 2880
rect 7848 2880 7866 2898
rect 7848 2898 7866 2916
rect 7848 2916 7866 2934
rect 7848 2934 7866 2952
rect 7848 2952 7866 2970
rect 7848 2970 7866 2988
rect 7848 2988 7866 3006
rect 7848 3006 7866 3024
rect 7848 3024 7866 3042
rect 7848 3042 7866 3060
rect 7848 3060 7866 3078
rect 7848 3078 7866 3096
rect 7848 3096 7866 3114
rect 7848 3114 7866 3132
rect 7848 3132 7866 3150
rect 7848 3150 7866 3168
rect 7848 3168 7866 3186
rect 7848 3186 7866 3204
rect 7848 3204 7866 3222
rect 7848 3222 7866 3240
rect 7848 3240 7866 3258
rect 7848 3258 7866 3276
rect 7848 3276 7866 3294
rect 7848 3294 7866 3312
rect 7848 3312 7866 3330
rect 7848 5076 7866 5094
rect 7848 5094 7866 5112
rect 7848 5112 7866 5130
rect 7848 5130 7866 5148
rect 7848 5148 7866 5166
rect 7848 5166 7866 5184
rect 7848 5184 7866 5202
rect 7848 5202 7866 5220
rect 7848 5220 7866 5238
rect 7848 5238 7866 5256
rect 7848 5256 7866 5274
rect 7848 5274 7866 5292
rect 7848 5292 7866 5310
rect 7848 5310 7866 5328
rect 7848 5328 7866 5346
rect 7848 5346 7866 5364
rect 7848 5364 7866 5382
rect 7848 5382 7866 5400
rect 7848 5400 7866 5418
rect 7848 5418 7866 5436
rect 7848 5436 7866 5454
rect 7848 5454 7866 5472
rect 7848 5472 7866 5490
rect 7848 5490 7866 5508
rect 7848 5508 7866 5526
rect 7848 5526 7866 5544
rect 7848 5544 7866 5562
rect 7848 5562 7866 5580
rect 7848 5580 7866 5598
rect 7848 5598 7866 5616
rect 7848 5616 7866 5634
rect 7848 5634 7866 5652
rect 7848 5652 7866 5670
rect 7848 5670 7866 5688
rect 7848 5688 7866 5706
rect 7848 5706 7866 5724
rect 7848 5724 7866 5742
rect 7848 5742 7866 5760
rect 7848 5760 7866 5778
rect 7848 5778 7866 5796
rect 7848 5796 7866 5814
rect 7848 5814 7866 5832
rect 7848 5832 7866 5850
rect 7848 5850 7866 5868
rect 7848 5868 7866 5886
rect 7848 5886 7866 5904
rect 7848 5904 7866 5922
rect 7848 5922 7866 5940
rect 7848 5940 7866 5958
rect 7848 5958 7866 5976
rect 7848 5976 7866 5994
rect 7848 5994 7866 6012
rect 7848 6012 7866 6030
rect 7848 6030 7866 6048
rect 7848 6048 7866 6066
rect 7848 6066 7866 6084
rect 7848 6084 7866 6102
rect 7848 6102 7866 6120
rect 7848 6120 7866 6138
rect 7848 6138 7866 6156
rect 7848 6156 7866 6174
rect 7848 6174 7866 6192
rect 7848 6192 7866 6210
rect 7848 6210 7866 6228
rect 7848 6228 7866 6246
rect 7848 6246 7866 6264
rect 7848 6264 7866 6282
rect 7848 6282 7866 6300
rect 7848 6300 7866 6318
rect 7848 6318 7866 6336
rect 7848 6336 7866 6354
rect 7848 6354 7866 6372
rect 7848 6372 7866 6390
rect 7848 6390 7866 6408
rect 7848 6408 7866 6426
rect 7848 6426 7866 6444
rect 7848 6444 7866 6462
rect 7848 6462 7866 6480
rect 7848 6480 7866 6498
rect 7848 6498 7866 6516
rect 7848 6516 7866 6534
rect 7848 6534 7866 6552
rect 7848 6552 7866 6570
rect 7848 6570 7866 6588
rect 7848 6588 7866 6606
rect 7848 6606 7866 6624
rect 7848 6624 7866 6642
rect 7848 6642 7866 6660
rect 7848 6660 7866 6678
rect 7848 6678 7866 6696
rect 7848 6696 7866 6714
rect 7848 6714 7866 6732
rect 7848 6732 7866 6750
rect 7848 6750 7866 6768
rect 7848 6768 7866 6786
rect 7848 6786 7866 6804
rect 7848 6804 7866 6822
rect 7848 6822 7866 6840
rect 7848 6840 7866 6858
rect 7848 6858 7866 6876
rect 7848 6876 7866 6894
rect 7848 6894 7866 6912
rect 7866 2322 7884 2340
rect 7866 2340 7884 2358
rect 7866 2358 7884 2376
rect 7866 2376 7884 2394
rect 7866 2394 7884 2412
rect 7866 2412 7884 2430
rect 7866 2430 7884 2448
rect 7866 2448 7884 2466
rect 7866 2466 7884 2484
rect 7866 2484 7884 2502
rect 7866 2502 7884 2520
rect 7866 2520 7884 2538
rect 7866 2538 7884 2556
rect 7866 2556 7884 2574
rect 7866 2574 7884 2592
rect 7866 2592 7884 2610
rect 7866 2610 7884 2628
rect 7866 2628 7884 2646
rect 7866 2646 7884 2664
rect 7866 2664 7884 2682
rect 7866 2682 7884 2700
rect 7866 2700 7884 2718
rect 7866 2718 7884 2736
rect 7866 2736 7884 2754
rect 7866 2754 7884 2772
rect 7866 2772 7884 2790
rect 7866 2790 7884 2808
rect 7866 2808 7884 2826
rect 7866 2826 7884 2844
rect 7866 2844 7884 2862
rect 7866 2862 7884 2880
rect 7866 2880 7884 2898
rect 7866 2898 7884 2916
rect 7866 2916 7884 2934
rect 7866 2934 7884 2952
rect 7866 2952 7884 2970
rect 7866 2970 7884 2988
rect 7866 2988 7884 3006
rect 7866 3006 7884 3024
rect 7866 3024 7884 3042
rect 7866 3042 7884 3060
rect 7866 3060 7884 3078
rect 7866 3078 7884 3096
rect 7866 3096 7884 3114
rect 7866 3114 7884 3132
rect 7866 3132 7884 3150
rect 7866 3150 7884 3168
rect 7866 3168 7884 3186
rect 7866 3186 7884 3204
rect 7866 3204 7884 3222
rect 7866 3222 7884 3240
rect 7866 3240 7884 3258
rect 7866 3258 7884 3276
rect 7866 3276 7884 3294
rect 7866 3294 7884 3312
rect 7866 3312 7884 3330
rect 7866 5094 7884 5112
rect 7866 5112 7884 5130
rect 7866 5130 7884 5148
rect 7866 5148 7884 5166
rect 7866 5166 7884 5184
rect 7866 5184 7884 5202
rect 7866 5202 7884 5220
rect 7866 5220 7884 5238
rect 7866 5238 7884 5256
rect 7866 5256 7884 5274
rect 7866 5274 7884 5292
rect 7866 5292 7884 5310
rect 7866 5310 7884 5328
rect 7866 5328 7884 5346
rect 7866 5346 7884 5364
rect 7866 5364 7884 5382
rect 7866 5382 7884 5400
rect 7866 5400 7884 5418
rect 7866 5418 7884 5436
rect 7866 5436 7884 5454
rect 7866 5454 7884 5472
rect 7866 5472 7884 5490
rect 7866 5490 7884 5508
rect 7866 5508 7884 5526
rect 7866 5526 7884 5544
rect 7866 5544 7884 5562
rect 7866 5562 7884 5580
rect 7866 5580 7884 5598
rect 7866 5598 7884 5616
rect 7866 5616 7884 5634
rect 7866 5634 7884 5652
rect 7866 5652 7884 5670
rect 7866 5670 7884 5688
rect 7866 5688 7884 5706
rect 7866 5706 7884 5724
rect 7866 5724 7884 5742
rect 7866 5742 7884 5760
rect 7866 5760 7884 5778
rect 7866 5778 7884 5796
rect 7866 5796 7884 5814
rect 7866 5814 7884 5832
rect 7866 5832 7884 5850
rect 7866 5850 7884 5868
rect 7866 5868 7884 5886
rect 7866 5886 7884 5904
rect 7866 5904 7884 5922
rect 7866 5922 7884 5940
rect 7866 5940 7884 5958
rect 7866 5958 7884 5976
rect 7866 5976 7884 5994
rect 7866 5994 7884 6012
rect 7866 6012 7884 6030
rect 7866 6030 7884 6048
rect 7866 6048 7884 6066
rect 7866 6066 7884 6084
rect 7866 6084 7884 6102
rect 7866 6102 7884 6120
rect 7866 6120 7884 6138
rect 7866 6138 7884 6156
rect 7866 6156 7884 6174
rect 7866 6174 7884 6192
rect 7866 6192 7884 6210
rect 7866 6210 7884 6228
rect 7866 6228 7884 6246
rect 7866 6246 7884 6264
rect 7866 6264 7884 6282
rect 7866 6282 7884 6300
rect 7866 6300 7884 6318
rect 7866 6318 7884 6336
rect 7866 6336 7884 6354
rect 7866 6354 7884 6372
rect 7866 6372 7884 6390
rect 7866 6390 7884 6408
rect 7866 6408 7884 6426
rect 7866 6426 7884 6444
rect 7866 6444 7884 6462
rect 7866 6462 7884 6480
rect 7866 6480 7884 6498
rect 7866 6498 7884 6516
rect 7866 6516 7884 6534
rect 7866 6534 7884 6552
rect 7866 6552 7884 6570
rect 7866 6570 7884 6588
rect 7866 6588 7884 6606
rect 7866 6606 7884 6624
rect 7866 6624 7884 6642
rect 7866 6642 7884 6660
rect 7866 6660 7884 6678
rect 7866 6678 7884 6696
rect 7866 6696 7884 6714
rect 7866 6714 7884 6732
rect 7866 6732 7884 6750
rect 7866 6750 7884 6768
rect 7866 6768 7884 6786
rect 7866 6786 7884 6804
rect 7866 6804 7884 6822
rect 7866 6822 7884 6840
rect 7866 6840 7884 6858
rect 7866 6858 7884 6876
rect 7866 6876 7884 6894
rect 7866 6894 7884 6912
rect 7866 6912 7884 6930
rect 7884 2322 7902 2340
rect 7884 2340 7902 2358
rect 7884 2358 7902 2376
rect 7884 2376 7902 2394
rect 7884 2394 7902 2412
rect 7884 2412 7902 2430
rect 7884 2430 7902 2448
rect 7884 2448 7902 2466
rect 7884 2466 7902 2484
rect 7884 2484 7902 2502
rect 7884 2502 7902 2520
rect 7884 2520 7902 2538
rect 7884 2538 7902 2556
rect 7884 2556 7902 2574
rect 7884 2574 7902 2592
rect 7884 2592 7902 2610
rect 7884 2610 7902 2628
rect 7884 2628 7902 2646
rect 7884 2646 7902 2664
rect 7884 2664 7902 2682
rect 7884 2682 7902 2700
rect 7884 2700 7902 2718
rect 7884 2718 7902 2736
rect 7884 2736 7902 2754
rect 7884 2754 7902 2772
rect 7884 2772 7902 2790
rect 7884 2790 7902 2808
rect 7884 2808 7902 2826
rect 7884 2826 7902 2844
rect 7884 2844 7902 2862
rect 7884 2862 7902 2880
rect 7884 2880 7902 2898
rect 7884 2898 7902 2916
rect 7884 2916 7902 2934
rect 7884 2934 7902 2952
rect 7884 2952 7902 2970
rect 7884 2970 7902 2988
rect 7884 2988 7902 3006
rect 7884 3006 7902 3024
rect 7884 3024 7902 3042
rect 7884 3042 7902 3060
rect 7884 3060 7902 3078
rect 7884 3078 7902 3096
rect 7884 3096 7902 3114
rect 7884 3114 7902 3132
rect 7884 3132 7902 3150
rect 7884 3150 7902 3168
rect 7884 3168 7902 3186
rect 7884 3186 7902 3204
rect 7884 3204 7902 3222
rect 7884 3222 7902 3240
rect 7884 3240 7902 3258
rect 7884 3258 7902 3276
rect 7884 3276 7902 3294
rect 7884 3294 7902 3312
rect 7884 3312 7902 3330
rect 7884 5112 7902 5130
rect 7884 5130 7902 5148
rect 7884 5148 7902 5166
rect 7884 5166 7902 5184
rect 7884 5184 7902 5202
rect 7884 5202 7902 5220
rect 7884 5220 7902 5238
rect 7884 5238 7902 5256
rect 7884 5256 7902 5274
rect 7884 5274 7902 5292
rect 7884 5292 7902 5310
rect 7884 5310 7902 5328
rect 7884 5328 7902 5346
rect 7884 5346 7902 5364
rect 7884 5364 7902 5382
rect 7884 5382 7902 5400
rect 7884 5400 7902 5418
rect 7884 5418 7902 5436
rect 7884 5436 7902 5454
rect 7884 5454 7902 5472
rect 7884 5472 7902 5490
rect 7884 5490 7902 5508
rect 7884 5508 7902 5526
rect 7884 5526 7902 5544
rect 7884 5544 7902 5562
rect 7884 5562 7902 5580
rect 7884 5580 7902 5598
rect 7884 5598 7902 5616
rect 7884 5616 7902 5634
rect 7884 5634 7902 5652
rect 7884 5652 7902 5670
rect 7884 5670 7902 5688
rect 7884 5688 7902 5706
rect 7884 5706 7902 5724
rect 7884 5724 7902 5742
rect 7884 5742 7902 5760
rect 7884 5760 7902 5778
rect 7884 5778 7902 5796
rect 7884 5796 7902 5814
rect 7884 5814 7902 5832
rect 7884 5832 7902 5850
rect 7884 5850 7902 5868
rect 7884 5868 7902 5886
rect 7884 5886 7902 5904
rect 7884 5904 7902 5922
rect 7884 5922 7902 5940
rect 7884 5940 7902 5958
rect 7884 5958 7902 5976
rect 7884 5976 7902 5994
rect 7884 5994 7902 6012
rect 7884 6012 7902 6030
rect 7884 6030 7902 6048
rect 7884 6048 7902 6066
rect 7884 6066 7902 6084
rect 7884 6084 7902 6102
rect 7884 6102 7902 6120
rect 7884 6120 7902 6138
rect 7884 6138 7902 6156
rect 7884 6156 7902 6174
rect 7884 6174 7902 6192
rect 7884 6192 7902 6210
rect 7884 6210 7902 6228
rect 7884 6228 7902 6246
rect 7884 6246 7902 6264
rect 7884 6264 7902 6282
rect 7884 6282 7902 6300
rect 7884 6300 7902 6318
rect 7884 6318 7902 6336
rect 7884 6336 7902 6354
rect 7884 6354 7902 6372
rect 7884 6372 7902 6390
rect 7884 6390 7902 6408
rect 7884 6408 7902 6426
rect 7884 6426 7902 6444
rect 7884 6444 7902 6462
rect 7884 6462 7902 6480
rect 7884 6480 7902 6498
rect 7884 6498 7902 6516
rect 7884 6516 7902 6534
rect 7884 6534 7902 6552
rect 7884 6552 7902 6570
rect 7884 6570 7902 6588
rect 7884 6588 7902 6606
rect 7884 6606 7902 6624
rect 7884 6624 7902 6642
rect 7884 6642 7902 6660
rect 7884 6660 7902 6678
rect 7884 6678 7902 6696
rect 7884 6696 7902 6714
rect 7884 6714 7902 6732
rect 7884 6732 7902 6750
rect 7884 6750 7902 6768
rect 7884 6768 7902 6786
rect 7884 6786 7902 6804
rect 7884 6804 7902 6822
rect 7884 6822 7902 6840
rect 7884 6840 7902 6858
rect 7884 6858 7902 6876
rect 7884 6876 7902 6894
rect 7884 6894 7902 6912
rect 7884 6912 7902 6930
rect 7884 6930 7902 6948
rect 7902 2340 7920 2358
rect 7902 2358 7920 2376
rect 7902 2376 7920 2394
rect 7902 2394 7920 2412
rect 7902 2412 7920 2430
rect 7902 2430 7920 2448
rect 7902 2448 7920 2466
rect 7902 2466 7920 2484
rect 7902 2484 7920 2502
rect 7902 2502 7920 2520
rect 7902 2520 7920 2538
rect 7902 2538 7920 2556
rect 7902 2556 7920 2574
rect 7902 2574 7920 2592
rect 7902 2592 7920 2610
rect 7902 2610 7920 2628
rect 7902 2628 7920 2646
rect 7902 2646 7920 2664
rect 7902 2664 7920 2682
rect 7902 2682 7920 2700
rect 7902 2700 7920 2718
rect 7902 2718 7920 2736
rect 7902 2736 7920 2754
rect 7902 2754 7920 2772
rect 7902 2772 7920 2790
rect 7902 2790 7920 2808
rect 7902 2808 7920 2826
rect 7902 2826 7920 2844
rect 7902 2844 7920 2862
rect 7902 2862 7920 2880
rect 7902 2880 7920 2898
rect 7902 2898 7920 2916
rect 7902 2916 7920 2934
rect 7902 2934 7920 2952
rect 7902 2952 7920 2970
rect 7902 2970 7920 2988
rect 7902 2988 7920 3006
rect 7902 3006 7920 3024
rect 7902 3024 7920 3042
rect 7902 3042 7920 3060
rect 7902 3060 7920 3078
rect 7902 3078 7920 3096
rect 7902 3096 7920 3114
rect 7902 3114 7920 3132
rect 7902 3132 7920 3150
rect 7902 3150 7920 3168
rect 7902 3168 7920 3186
rect 7902 3186 7920 3204
rect 7902 3204 7920 3222
rect 7902 3222 7920 3240
rect 7902 3240 7920 3258
rect 7902 3258 7920 3276
rect 7902 3276 7920 3294
rect 7902 3294 7920 3312
rect 7902 3312 7920 3330
rect 7902 3330 7920 3348
rect 7902 5148 7920 5166
rect 7902 5166 7920 5184
rect 7902 5184 7920 5202
rect 7902 5202 7920 5220
rect 7902 5220 7920 5238
rect 7902 5238 7920 5256
rect 7902 5256 7920 5274
rect 7902 5274 7920 5292
rect 7902 5292 7920 5310
rect 7902 5310 7920 5328
rect 7902 5328 7920 5346
rect 7902 5346 7920 5364
rect 7902 5364 7920 5382
rect 7902 5382 7920 5400
rect 7902 5400 7920 5418
rect 7902 5418 7920 5436
rect 7902 5436 7920 5454
rect 7902 5454 7920 5472
rect 7902 5472 7920 5490
rect 7902 5490 7920 5508
rect 7902 5508 7920 5526
rect 7902 5526 7920 5544
rect 7902 5544 7920 5562
rect 7902 5562 7920 5580
rect 7902 5580 7920 5598
rect 7902 5598 7920 5616
rect 7902 5616 7920 5634
rect 7902 5634 7920 5652
rect 7902 5652 7920 5670
rect 7902 5670 7920 5688
rect 7902 5688 7920 5706
rect 7902 5706 7920 5724
rect 7902 5724 7920 5742
rect 7902 5742 7920 5760
rect 7902 5760 7920 5778
rect 7902 5778 7920 5796
rect 7902 5796 7920 5814
rect 7902 5814 7920 5832
rect 7902 5832 7920 5850
rect 7902 5850 7920 5868
rect 7902 5868 7920 5886
rect 7902 5886 7920 5904
rect 7902 5904 7920 5922
rect 7902 5922 7920 5940
rect 7902 5940 7920 5958
rect 7902 5958 7920 5976
rect 7902 5976 7920 5994
rect 7902 5994 7920 6012
rect 7902 6012 7920 6030
rect 7902 6030 7920 6048
rect 7902 6048 7920 6066
rect 7902 6066 7920 6084
rect 7902 6084 7920 6102
rect 7902 6102 7920 6120
rect 7902 6120 7920 6138
rect 7902 6138 7920 6156
rect 7902 6156 7920 6174
rect 7902 6174 7920 6192
rect 7902 6192 7920 6210
rect 7902 6210 7920 6228
rect 7902 6228 7920 6246
rect 7902 6246 7920 6264
rect 7902 6264 7920 6282
rect 7902 6282 7920 6300
rect 7902 6300 7920 6318
rect 7902 6318 7920 6336
rect 7902 6336 7920 6354
rect 7902 6354 7920 6372
rect 7902 6372 7920 6390
rect 7902 6390 7920 6408
rect 7902 6408 7920 6426
rect 7902 6426 7920 6444
rect 7902 6444 7920 6462
rect 7902 6462 7920 6480
rect 7902 6480 7920 6498
rect 7902 6498 7920 6516
rect 7902 6516 7920 6534
rect 7902 6534 7920 6552
rect 7902 6552 7920 6570
rect 7902 6570 7920 6588
rect 7902 6588 7920 6606
rect 7902 6606 7920 6624
rect 7902 6624 7920 6642
rect 7902 6642 7920 6660
rect 7902 6660 7920 6678
rect 7902 6678 7920 6696
rect 7902 6696 7920 6714
rect 7902 6714 7920 6732
rect 7902 6732 7920 6750
rect 7902 6750 7920 6768
rect 7902 6768 7920 6786
rect 7902 6786 7920 6804
rect 7902 6804 7920 6822
rect 7902 6822 7920 6840
rect 7902 6840 7920 6858
rect 7902 6858 7920 6876
rect 7902 6876 7920 6894
rect 7902 6894 7920 6912
rect 7902 6912 7920 6930
rect 7902 6930 7920 6948
rect 7920 2358 7938 2376
rect 7920 2376 7938 2394
rect 7920 2394 7938 2412
rect 7920 2412 7938 2430
rect 7920 2430 7938 2448
rect 7920 2448 7938 2466
rect 7920 2466 7938 2484
rect 7920 2484 7938 2502
rect 7920 2502 7938 2520
rect 7920 2520 7938 2538
rect 7920 2538 7938 2556
rect 7920 2556 7938 2574
rect 7920 2574 7938 2592
rect 7920 2592 7938 2610
rect 7920 2610 7938 2628
rect 7920 2628 7938 2646
rect 7920 2646 7938 2664
rect 7920 2664 7938 2682
rect 7920 2682 7938 2700
rect 7920 2700 7938 2718
rect 7920 2718 7938 2736
rect 7920 2736 7938 2754
rect 7920 2754 7938 2772
rect 7920 2772 7938 2790
rect 7920 2790 7938 2808
rect 7920 2808 7938 2826
rect 7920 2826 7938 2844
rect 7920 2844 7938 2862
rect 7920 2862 7938 2880
rect 7920 2880 7938 2898
rect 7920 2898 7938 2916
rect 7920 2916 7938 2934
rect 7920 2934 7938 2952
rect 7920 2952 7938 2970
rect 7920 2970 7938 2988
rect 7920 2988 7938 3006
rect 7920 3006 7938 3024
rect 7920 3024 7938 3042
rect 7920 3042 7938 3060
rect 7920 3060 7938 3078
rect 7920 3078 7938 3096
rect 7920 3096 7938 3114
rect 7920 3114 7938 3132
rect 7920 3132 7938 3150
rect 7920 3150 7938 3168
rect 7920 3168 7938 3186
rect 7920 3186 7938 3204
rect 7920 3204 7938 3222
rect 7920 3222 7938 3240
rect 7920 3240 7938 3258
rect 7920 3258 7938 3276
rect 7920 3276 7938 3294
rect 7920 3294 7938 3312
rect 7920 3312 7938 3330
rect 7920 3330 7938 3348
rect 7920 5166 7938 5184
rect 7920 5184 7938 5202
rect 7920 5202 7938 5220
rect 7920 5220 7938 5238
rect 7920 5238 7938 5256
rect 7920 5256 7938 5274
rect 7920 5274 7938 5292
rect 7920 5292 7938 5310
rect 7920 5310 7938 5328
rect 7920 5328 7938 5346
rect 7920 5346 7938 5364
rect 7920 5364 7938 5382
rect 7920 5382 7938 5400
rect 7920 5400 7938 5418
rect 7920 5418 7938 5436
rect 7920 5436 7938 5454
rect 7920 5454 7938 5472
rect 7920 5472 7938 5490
rect 7920 5490 7938 5508
rect 7920 5508 7938 5526
rect 7920 5526 7938 5544
rect 7920 5544 7938 5562
rect 7920 5562 7938 5580
rect 7920 5580 7938 5598
rect 7920 5598 7938 5616
rect 7920 5616 7938 5634
rect 7920 5634 7938 5652
rect 7920 5652 7938 5670
rect 7920 5670 7938 5688
rect 7920 5688 7938 5706
rect 7920 5706 7938 5724
rect 7920 5724 7938 5742
rect 7920 5742 7938 5760
rect 7920 5760 7938 5778
rect 7920 5778 7938 5796
rect 7920 5796 7938 5814
rect 7920 5814 7938 5832
rect 7920 5832 7938 5850
rect 7920 5850 7938 5868
rect 7920 5868 7938 5886
rect 7920 5886 7938 5904
rect 7920 5904 7938 5922
rect 7920 5922 7938 5940
rect 7920 5940 7938 5958
rect 7920 5958 7938 5976
rect 7920 5976 7938 5994
rect 7920 5994 7938 6012
rect 7920 6012 7938 6030
rect 7920 6030 7938 6048
rect 7920 6048 7938 6066
rect 7920 6066 7938 6084
rect 7920 6084 7938 6102
rect 7920 6102 7938 6120
rect 7920 6120 7938 6138
rect 7920 6138 7938 6156
rect 7920 6156 7938 6174
rect 7920 6174 7938 6192
rect 7920 6192 7938 6210
rect 7920 6210 7938 6228
rect 7920 6228 7938 6246
rect 7920 6246 7938 6264
rect 7920 6264 7938 6282
rect 7920 6282 7938 6300
rect 7920 6300 7938 6318
rect 7920 6318 7938 6336
rect 7920 6336 7938 6354
rect 7920 6354 7938 6372
rect 7920 6372 7938 6390
rect 7920 6390 7938 6408
rect 7920 6408 7938 6426
rect 7920 6426 7938 6444
rect 7920 6444 7938 6462
rect 7920 6462 7938 6480
rect 7920 6480 7938 6498
rect 7920 6498 7938 6516
rect 7920 6516 7938 6534
rect 7920 6534 7938 6552
rect 7920 6552 7938 6570
rect 7920 6570 7938 6588
rect 7920 6588 7938 6606
rect 7920 6606 7938 6624
rect 7920 6624 7938 6642
rect 7920 6642 7938 6660
rect 7920 6660 7938 6678
rect 7920 6678 7938 6696
rect 7920 6696 7938 6714
rect 7920 6714 7938 6732
rect 7920 6732 7938 6750
rect 7920 6750 7938 6768
rect 7920 6768 7938 6786
rect 7920 6786 7938 6804
rect 7920 6804 7938 6822
rect 7920 6822 7938 6840
rect 7920 6840 7938 6858
rect 7920 6858 7938 6876
rect 7920 6876 7938 6894
rect 7920 6894 7938 6912
rect 7920 6912 7938 6930
rect 7920 6930 7938 6948
rect 7920 6948 7938 6966
rect 7938 2358 7956 2376
rect 7938 2376 7956 2394
rect 7938 2394 7956 2412
rect 7938 2412 7956 2430
rect 7938 2430 7956 2448
rect 7938 2448 7956 2466
rect 7938 2466 7956 2484
rect 7938 2484 7956 2502
rect 7938 2502 7956 2520
rect 7938 2520 7956 2538
rect 7938 2538 7956 2556
rect 7938 2556 7956 2574
rect 7938 2574 7956 2592
rect 7938 2592 7956 2610
rect 7938 2610 7956 2628
rect 7938 2628 7956 2646
rect 7938 2646 7956 2664
rect 7938 2664 7956 2682
rect 7938 2682 7956 2700
rect 7938 2700 7956 2718
rect 7938 2718 7956 2736
rect 7938 2736 7956 2754
rect 7938 2754 7956 2772
rect 7938 2772 7956 2790
rect 7938 2790 7956 2808
rect 7938 2808 7956 2826
rect 7938 2826 7956 2844
rect 7938 2844 7956 2862
rect 7938 2862 7956 2880
rect 7938 2880 7956 2898
rect 7938 2898 7956 2916
rect 7938 2916 7956 2934
rect 7938 2934 7956 2952
rect 7938 2952 7956 2970
rect 7938 2970 7956 2988
rect 7938 2988 7956 3006
rect 7938 3006 7956 3024
rect 7938 3024 7956 3042
rect 7938 3042 7956 3060
rect 7938 3060 7956 3078
rect 7938 3078 7956 3096
rect 7938 3096 7956 3114
rect 7938 3114 7956 3132
rect 7938 3132 7956 3150
rect 7938 3150 7956 3168
rect 7938 3168 7956 3186
rect 7938 3186 7956 3204
rect 7938 3204 7956 3222
rect 7938 3222 7956 3240
rect 7938 3240 7956 3258
rect 7938 3258 7956 3276
rect 7938 3276 7956 3294
rect 7938 3294 7956 3312
rect 7938 3312 7956 3330
rect 7938 3330 7956 3348
rect 7938 5184 7956 5202
rect 7938 5202 7956 5220
rect 7938 5220 7956 5238
rect 7938 5238 7956 5256
rect 7938 5256 7956 5274
rect 7938 5274 7956 5292
rect 7938 5292 7956 5310
rect 7938 5310 7956 5328
rect 7938 5328 7956 5346
rect 7938 5346 7956 5364
rect 7938 5364 7956 5382
rect 7938 5382 7956 5400
rect 7938 5400 7956 5418
rect 7938 5418 7956 5436
rect 7938 5436 7956 5454
rect 7938 5454 7956 5472
rect 7938 5472 7956 5490
rect 7938 5490 7956 5508
rect 7938 5508 7956 5526
rect 7938 5526 7956 5544
rect 7938 5544 7956 5562
rect 7938 5562 7956 5580
rect 7938 5580 7956 5598
rect 7938 5598 7956 5616
rect 7938 5616 7956 5634
rect 7938 5634 7956 5652
rect 7938 5652 7956 5670
rect 7938 5670 7956 5688
rect 7938 5688 7956 5706
rect 7938 5706 7956 5724
rect 7938 5724 7956 5742
rect 7938 5742 7956 5760
rect 7938 5760 7956 5778
rect 7938 5778 7956 5796
rect 7938 5796 7956 5814
rect 7938 5814 7956 5832
rect 7938 5832 7956 5850
rect 7938 5850 7956 5868
rect 7938 5868 7956 5886
rect 7938 5886 7956 5904
rect 7938 5904 7956 5922
rect 7938 5922 7956 5940
rect 7938 5940 7956 5958
rect 7938 5958 7956 5976
rect 7938 5976 7956 5994
rect 7938 5994 7956 6012
rect 7938 6012 7956 6030
rect 7938 6030 7956 6048
rect 7938 6048 7956 6066
rect 7938 6066 7956 6084
rect 7938 6084 7956 6102
rect 7938 6102 7956 6120
rect 7938 6120 7956 6138
rect 7938 6138 7956 6156
rect 7938 6156 7956 6174
rect 7938 6174 7956 6192
rect 7938 6192 7956 6210
rect 7938 6210 7956 6228
rect 7938 6228 7956 6246
rect 7938 6246 7956 6264
rect 7938 6264 7956 6282
rect 7938 6282 7956 6300
rect 7938 6300 7956 6318
rect 7938 6318 7956 6336
rect 7938 6336 7956 6354
rect 7938 6354 7956 6372
rect 7938 6372 7956 6390
rect 7938 6390 7956 6408
rect 7938 6408 7956 6426
rect 7938 6426 7956 6444
rect 7938 6444 7956 6462
rect 7938 6462 7956 6480
rect 7938 6480 7956 6498
rect 7938 6498 7956 6516
rect 7938 6516 7956 6534
rect 7938 6534 7956 6552
rect 7938 6552 7956 6570
rect 7938 6570 7956 6588
rect 7938 6588 7956 6606
rect 7938 6606 7956 6624
rect 7938 6624 7956 6642
rect 7938 6642 7956 6660
rect 7938 6660 7956 6678
rect 7938 6678 7956 6696
rect 7938 6696 7956 6714
rect 7938 6714 7956 6732
rect 7938 6732 7956 6750
rect 7938 6750 7956 6768
rect 7938 6768 7956 6786
rect 7938 6786 7956 6804
rect 7938 6804 7956 6822
rect 7938 6822 7956 6840
rect 7938 6840 7956 6858
rect 7938 6858 7956 6876
rect 7938 6876 7956 6894
rect 7938 6894 7956 6912
rect 7938 6912 7956 6930
rect 7938 6930 7956 6948
rect 7938 6948 7956 6966
rect 7938 6966 7956 6984
rect 7956 2376 7974 2394
rect 7956 2394 7974 2412
rect 7956 2412 7974 2430
rect 7956 2430 7974 2448
rect 7956 2448 7974 2466
rect 7956 2466 7974 2484
rect 7956 2484 7974 2502
rect 7956 2502 7974 2520
rect 7956 2520 7974 2538
rect 7956 2538 7974 2556
rect 7956 2556 7974 2574
rect 7956 2574 7974 2592
rect 7956 2592 7974 2610
rect 7956 2610 7974 2628
rect 7956 2628 7974 2646
rect 7956 2646 7974 2664
rect 7956 2664 7974 2682
rect 7956 2682 7974 2700
rect 7956 2700 7974 2718
rect 7956 2718 7974 2736
rect 7956 2736 7974 2754
rect 7956 2754 7974 2772
rect 7956 2772 7974 2790
rect 7956 2790 7974 2808
rect 7956 2808 7974 2826
rect 7956 2826 7974 2844
rect 7956 2844 7974 2862
rect 7956 2862 7974 2880
rect 7956 2880 7974 2898
rect 7956 2898 7974 2916
rect 7956 2916 7974 2934
rect 7956 2934 7974 2952
rect 7956 2952 7974 2970
rect 7956 2970 7974 2988
rect 7956 2988 7974 3006
rect 7956 3006 7974 3024
rect 7956 3024 7974 3042
rect 7956 3042 7974 3060
rect 7956 3060 7974 3078
rect 7956 3078 7974 3096
rect 7956 3096 7974 3114
rect 7956 3114 7974 3132
rect 7956 3132 7974 3150
rect 7956 3150 7974 3168
rect 7956 3168 7974 3186
rect 7956 3186 7974 3204
rect 7956 3204 7974 3222
rect 7956 3222 7974 3240
rect 7956 3240 7974 3258
rect 7956 3258 7974 3276
rect 7956 3276 7974 3294
rect 7956 3294 7974 3312
rect 7956 3312 7974 3330
rect 7956 3330 7974 3348
rect 7956 5220 7974 5238
rect 7956 5238 7974 5256
rect 7956 5256 7974 5274
rect 7956 5274 7974 5292
rect 7956 5292 7974 5310
rect 7956 5310 7974 5328
rect 7956 5328 7974 5346
rect 7956 5346 7974 5364
rect 7956 5364 7974 5382
rect 7956 5382 7974 5400
rect 7956 5400 7974 5418
rect 7956 5418 7974 5436
rect 7956 5436 7974 5454
rect 7956 5454 7974 5472
rect 7956 5472 7974 5490
rect 7956 5490 7974 5508
rect 7956 5508 7974 5526
rect 7956 5526 7974 5544
rect 7956 5544 7974 5562
rect 7956 5562 7974 5580
rect 7956 5580 7974 5598
rect 7956 5598 7974 5616
rect 7956 5616 7974 5634
rect 7956 5634 7974 5652
rect 7956 5652 7974 5670
rect 7956 5670 7974 5688
rect 7956 5688 7974 5706
rect 7956 5706 7974 5724
rect 7956 5724 7974 5742
rect 7956 5742 7974 5760
rect 7956 5760 7974 5778
rect 7956 5778 7974 5796
rect 7956 5796 7974 5814
rect 7956 5814 7974 5832
rect 7956 5832 7974 5850
rect 7956 5850 7974 5868
rect 7956 5868 7974 5886
rect 7956 5886 7974 5904
rect 7956 5904 7974 5922
rect 7956 5922 7974 5940
rect 7956 5940 7974 5958
rect 7956 5958 7974 5976
rect 7956 5976 7974 5994
rect 7956 5994 7974 6012
rect 7956 6012 7974 6030
rect 7956 6030 7974 6048
rect 7956 6048 7974 6066
rect 7956 6066 7974 6084
rect 7956 6084 7974 6102
rect 7956 6102 7974 6120
rect 7956 6120 7974 6138
rect 7956 6138 7974 6156
rect 7956 6156 7974 6174
rect 7956 6174 7974 6192
rect 7956 6192 7974 6210
rect 7956 6210 7974 6228
rect 7956 6228 7974 6246
rect 7956 6246 7974 6264
rect 7956 6264 7974 6282
rect 7956 6282 7974 6300
rect 7956 6300 7974 6318
rect 7956 6318 7974 6336
rect 7956 6336 7974 6354
rect 7956 6354 7974 6372
rect 7956 6372 7974 6390
rect 7956 6390 7974 6408
rect 7956 6408 7974 6426
rect 7956 6426 7974 6444
rect 7956 6444 7974 6462
rect 7956 6462 7974 6480
rect 7956 6480 7974 6498
rect 7956 6498 7974 6516
rect 7956 6516 7974 6534
rect 7956 6534 7974 6552
rect 7956 6552 7974 6570
rect 7956 6570 7974 6588
rect 7956 6588 7974 6606
rect 7956 6606 7974 6624
rect 7956 6624 7974 6642
rect 7956 6642 7974 6660
rect 7956 6660 7974 6678
rect 7956 6678 7974 6696
rect 7956 6696 7974 6714
rect 7956 6714 7974 6732
rect 7956 6732 7974 6750
rect 7956 6750 7974 6768
rect 7956 6768 7974 6786
rect 7956 6786 7974 6804
rect 7956 6804 7974 6822
rect 7956 6822 7974 6840
rect 7956 6840 7974 6858
rect 7956 6858 7974 6876
rect 7956 6876 7974 6894
rect 7956 6894 7974 6912
rect 7956 6912 7974 6930
rect 7956 6930 7974 6948
rect 7956 6948 7974 6966
rect 7956 6966 7974 6984
rect 7956 6984 7974 7002
rect 7974 2394 7992 2412
rect 7974 2412 7992 2430
rect 7974 2430 7992 2448
rect 7974 2448 7992 2466
rect 7974 2466 7992 2484
rect 7974 2484 7992 2502
rect 7974 2502 7992 2520
rect 7974 2520 7992 2538
rect 7974 2538 7992 2556
rect 7974 2556 7992 2574
rect 7974 2574 7992 2592
rect 7974 2592 7992 2610
rect 7974 2610 7992 2628
rect 7974 2628 7992 2646
rect 7974 2646 7992 2664
rect 7974 2664 7992 2682
rect 7974 2682 7992 2700
rect 7974 2700 7992 2718
rect 7974 2718 7992 2736
rect 7974 2736 7992 2754
rect 7974 2754 7992 2772
rect 7974 2772 7992 2790
rect 7974 2790 7992 2808
rect 7974 2808 7992 2826
rect 7974 2826 7992 2844
rect 7974 2844 7992 2862
rect 7974 2862 7992 2880
rect 7974 2880 7992 2898
rect 7974 2898 7992 2916
rect 7974 2916 7992 2934
rect 7974 2934 7992 2952
rect 7974 2952 7992 2970
rect 7974 2970 7992 2988
rect 7974 2988 7992 3006
rect 7974 3006 7992 3024
rect 7974 3024 7992 3042
rect 7974 3042 7992 3060
rect 7974 3060 7992 3078
rect 7974 3078 7992 3096
rect 7974 3096 7992 3114
rect 7974 3114 7992 3132
rect 7974 3132 7992 3150
rect 7974 3150 7992 3168
rect 7974 3168 7992 3186
rect 7974 3186 7992 3204
rect 7974 3204 7992 3222
rect 7974 3222 7992 3240
rect 7974 3240 7992 3258
rect 7974 3258 7992 3276
rect 7974 3276 7992 3294
rect 7974 3294 7992 3312
rect 7974 3312 7992 3330
rect 7974 3330 7992 3348
rect 7974 3348 7992 3366
rect 7974 5238 7992 5256
rect 7974 5256 7992 5274
rect 7974 5274 7992 5292
rect 7974 5292 7992 5310
rect 7974 5310 7992 5328
rect 7974 5328 7992 5346
rect 7974 5346 7992 5364
rect 7974 5364 7992 5382
rect 7974 5382 7992 5400
rect 7974 5400 7992 5418
rect 7974 5418 7992 5436
rect 7974 5436 7992 5454
rect 7974 5454 7992 5472
rect 7974 5472 7992 5490
rect 7974 5490 7992 5508
rect 7974 5508 7992 5526
rect 7974 5526 7992 5544
rect 7974 5544 7992 5562
rect 7974 5562 7992 5580
rect 7974 5580 7992 5598
rect 7974 5598 7992 5616
rect 7974 5616 7992 5634
rect 7974 5634 7992 5652
rect 7974 5652 7992 5670
rect 7974 5670 7992 5688
rect 7974 5688 7992 5706
rect 7974 5706 7992 5724
rect 7974 5724 7992 5742
rect 7974 5742 7992 5760
rect 7974 5760 7992 5778
rect 7974 5778 7992 5796
rect 7974 5796 7992 5814
rect 7974 5814 7992 5832
rect 7974 5832 7992 5850
rect 7974 5850 7992 5868
rect 7974 5868 7992 5886
rect 7974 5886 7992 5904
rect 7974 5904 7992 5922
rect 7974 5922 7992 5940
rect 7974 5940 7992 5958
rect 7974 5958 7992 5976
rect 7974 5976 7992 5994
rect 7974 5994 7992 6012
rect 7974 6012 7992 6030
rect 7974 6030 7992 6048
rect 7974 6048 7992 6066
rect 7974 6066 7992 6084
rect 7974 6084 7992 6102
rect 7974 6102 7992 6120
rect 7974 6120 7992 6138
rect 7974 6138 7992 6156
rect 7974 6156 7992 6174
rect 7974 6174 7992 6192
rect 7974 6192 7992 6210
rect 7974 6210 7992 6228
rect 7974 6228 7992 6246
rect 7974 6246 7992 6264
rect 7974 6264 7992 6282
rect 7974 6282 7992 6300
rect 7974 6300 7992 6318
rect 7974 6318 7992 6336
rect 7974 6336 7992 6354
rect 7974 6354 7992 6372
rect 7974 6372 7992 6390
rect 7974 6390 7992 6408
rect 7974 6408 7992 6426
rect 7974 6426 7992 6444
rect 7974 6444 7992 6462
rect 7974 6462 7992 6480
rect 7974 6480 7992 6498
rect 7974 6498 7992 6516
rect 7974 6516 7992 6534
rect 7974 6534 7992 6552
rect 7974 6552 7992 6570
rect 7974 6570 7992 6588
rect 7974 6588 7992 6606
rect 7974 6606 7992 6624
rect 7974 6624 7992 6642
rect 7974 6642 7992 6660
rect 7974 6660 7992 6678
rect 7974 6678 7992 6696
rect 7974 6696 7992 6714
rect 7974 6714 7992 6732
rect 7974 6732 7992 6750
rect 7974 6750 7992 6768
rect 7974 6768 7992 6786
rect 7974 6786 7992 6804
rect 7974 6804 7992 6822
rect 7974 6822 7992 6840
rect 7974 6840 7992 6858
rect 7974 6858 7992 6876
rect 7974 6876 7992 6894
rect 7974 6894 7992 6912
rect 7974 6912 7992 6930
rect 7974 6930 7992 6948
rect 7974 6948 7992 6966
rect 7974 6966 7992 6984
rect 7974 6984 7992 7002
rect 7992 2394 8010 2412
rect 7992 2412 8010 2430
rect 7992 2430 8010 2448
rect 7992 2448 8010 2466
rect 7992 2466 8010 2484
rect 7992 2484 8010 2502
rect 7992 2502 8010 2520
rect 7992 2520 8010 2538
rect 7992 2538 8010 2556
rect 7992 2556 8010 2574
rect 7992 2574 8010 2592
rect 7992 2592 8010 2610
rect 7992 2610 8010 2628
rect 7992 2628 8010 2646
rect 7992 2646 8010 2664
rect 7992 2664 8010 2682
rect 7992 2682 8010 2700
rect 7992 2700 8010 2718
rect 7992 2718 8010 2736
rect 7992 2736 8010 2754
rect 7992 2754 8010 2772
rect 7992 2772 8010 2790
rect 7992 2790 8010 2808
rect 7992 2808 8010 2826
rect 7992 2826 8010 2844
rect 7992 2844 8010 2862
rect 7992 2862 8010 2880
rect 7992 2880 8010 2898
rect 7992 2898 8010 2916
rect 7992 2916 8010 2934
rect 7992 2934 8010 2952
rect 7992 2952 8010 2970
rect 7992 2970 8010 2988
rect 7992 2988 8010 3006
rect 7992 3006 8010 3024
rect 7992 3024 8010 3042
rect 7992 3042 8010 3060
rect 7992 3060 8010 3078
rect 7992 3078 8010 3096
rect 7992 3096 8010 3114
rect 7992 3114 8010 3132
rect 7992 3132 8010 3150
rect 7992 3150 8010 3168
rect 7992 3168 8010 3186
rect 7992 3186 8010 3204
rect 7992 3204 8010 3222
rect 7992 3222 8010 3240
rect 7992 3240 8010 3258
rect 7992 3258 8010 3276
rect 7992 3276 8010 3294
rect 7992 3294 8010 3312
rect 7992 3312 8010 3330
rect 7992 3330 8010 3348
rect 7992 3348 8010 3366
rect 7992 5256 8010 5274
rect 7992 5274 8010 5292
rect 7992 5292 8010 5310
rect 7992 5310 8010 5328
rect 7992 5328 8010 5346
rect 7992 5346 8010 5364
rect 7992 5364 8010 5382
rect 7992 5382 8010 5400
rect 7992 5400 8010 5418
rect 7992 5418 8010 5436
rect 7992 5436 8010 5454
rect 7992 5454 8010 5472
rect 7992 5472 8010 5490
rect 7992 5490 8010 5508
rect 7992 5508 8010 5526
rect 7992 5526 8010 5544
rect 7992 5544 8010 5562
rect 7992 5562 8010 5580
rect 7992 5580 8010 5598
rect 7992 5598 8010 5616
rect 7992 5616 8010 5634
rect 7992 5634 8010 5652
rect 7992 5652 8010 5670
rect 7992 5670 8010 5688
rect 7992 5688 8010 5706
rect 7992 5706 8010 5724
rect 7992 5724 8010 5742
rect 7992 5742 8010 5760
rect 7992 5760 8010 5778
rect 7992 5778 8010 5796
rect 7992 5796 8010 5814
rect 7992 5814 8010 5832
rect 7992 5832 8010 5850
rect 7992 5850 8010 5868
rect 7992 5868 8010 5886
rect 7992 5886 8010 5904
rect 7992 5904 8010 5922
rect 7992 5922 8010 5940
rect 7992 5940 8010 5958
rect 7992 5958 8010 5976
rect 7992 5976 8010 5994
rect 7992 5994 8010 6012
rect 7992 6012 8010 6030
rect 7992 6030 8010 6048
rect 7992 6048 8010 6066
rect 7992 6066 8010 6084
rect 7992 6084 8010 6102
rect 7992 6102 8010 6120
rect 7992 6120 8010 6138
rect 7992 6138 8010 6156
rect 7992 6156 8010 6174
rect 7992 6174 8010 6192
rect 7992 6192 8010 6210
rect 7992 6210 8010 6228
rect 7992 6228 8010 6246
rect 7992 6246 8010 6264
rect 7992 6264 8010 6282
rect 7992 6282 8010 6300
rect 7992 6300 8010 6318
rect 7992 6318 8010 6336
rect 7992 6336 8010 6354
rect 7992 6354 8010 6372
rect 7992 6372 8010 6390
rect 7992 6390 8010 6408
rect 7992 6408 8010 6426
rect 7992 6426 8010 6444
rect 7992 6444 8010 6462
rect 7992 6462 8010 6480
rect 7992 6480 8010 6498
rect 7992 6498 8010 6516
rect 7992 6516 8010 6534
rect 7992 6534 8010 6552
rect 7992 6552 8010 6570
rect 7992 6570 8010 6588
rect 7992 6588 8010 6606
rect 7992 6606 8010 6624
rect 7992 6624 8010 6642
rect 7992 6642 8010 6660
rect 7992 6660 8010 6678
rect 7992 6678 8010 6696
rect 7992 6696 8010 6714
rect 7992 6714 8010 6732
rect 7992 6732 8010 6750
rect 7992 6750 8010 6768
rect 7992 6768 8010 6786
rect 7992 6786 8010 6804
rect 7992 6804 8010 6822
rect 7992 6822 8010 6840
rect 7992 6840 8010 6858
rect 7992 6858 8010 6876
rect 7992 6876 8010 6894
rect 7992 6894 8010 6912
rect 7992 6912 8010 6930
rect 7992 6930 8010 6948
rect 7992 6948 8010 6966
rect 7992 6966 8010 6984
rect 7992 6984 8010 7002
rect 7992 7002 8010 7020
rect 8010 2412 8028 2430
rect 8010 2430 8028 2448
rect 8010 2448 8028 2466
rect 8010 2466 8028 2484
rect 8010 2484 8028 2502
rect 8010 2502 8028 2520
rect 8010 2520 8028 2538
rect 8010 2538 8028 2556
rect 8010 2556 8028 2574
rect 8010 2574 8028 2592
rect 8010 2592 8028 2610
rect 8010 2610 8028 2628
rect 8010 2628 8028 2646
rect 8010 2646 8028 2664
rect 8010 2664 8028 2682
rect 8010 2682 8028 2700
rect 8010 2700 8028 2718
rect 8010 2718 8028 2736
rect 8010 2736 8028 2754
rect 8010 2754 8028 2772
rect 8010 2772 8028 2790
rect 8010 2790 8028 2808
rect 8010 2808 8028 2826
rect 8010 2826 8028 2844
rect 8010 2844 8028 2862
rect 8010 2862 8028 2880
rect 8010 2880 8028 2898
rect 8010 2898 8028 2916
rect 8010 2916 8028 2934
rect 8010 2934 8028 2952
rect 8010 2952 8028 2970
rect 8010 2970 8028 2988
rect 8010 2988 8028 3006
rect 8010 3006 8028 3024
rect 8010 3024 8028 3042
rect 8010 3042 8028 3060
rect 8010 3060 8028 3078
rect 8010 3078 8028 3096
rect 8010 3096 8028 3114
rect 8010 3114 8028 3132
rect 8010 3132 8028 3150
rect 8010 3150 8028 3168
rect 8010 3168 8028 3186
rect 8010 3186 8028 3204
rect 8010 3204 8028 3222
rect 8010 3222 8028 3240
rect 8010 3240 8028 3258
rect 8010 3258 8028 3276
rect 8010 3276 8028 3294
rect 8010 3294 8028 3312
rect 8010 3312 8028 3330
rect 8010 3330 8028 3348
rect 8010 3348 8028 3366
rect 8010 5274 8028 5292
rect 8010 5292 8028 5310
rect 8010 5310 8028 5328
rect 8010 5328 8028 5346
rect 8010 5346 8028 5364
rect 8010 5364 8028 5382
rect 8010 5382 8028 5400
rect 8010 5400 8028 5418
rect 8010 5418 8028 5436
rect 8010 5436 8028 5454
rect 8010 5454 8028 5472
rect 8010 5472 8028 5490
rect 8010 5490 8028 5508
rect 8010 5508 8028 5526
rect 8010 5526 8028 5544
rect 8010 5544 8028 5562
rect 8010 5562 8028 5580
rect 8010 5580 8028 5598
rect 8010 5598 8028 5616
rect 8010 5616 8028 5634
rect 8010 5634 8028 5652
rect 8010 5652 8028 5670
rect 8010 5670 8028 5688
rect 8010 5688 8028 5706
rect 8010 5706 8028 5724
rect 8010 5724 8028 5742
rect 8010 5742 8028 5760
rect 8010 5760 8028 5778
rect 8010 5778 8028 5796
rect 8010 5796 8028 5814
rect 8010 5814 8028 5832
rect 8010 5832 8028 5850
rect 8010 5850 8028 5868
rect 8010 5868 8028 5886
rect 8010 5886 8028 5904
rect 8010 5904 8028 5922
rect 8010 5922 8028 5940
rect 8010 5940 8028 5958
rect 8010 5958 8028 5976
rect 8010 5976 8028 5994
rect 8010 5994 8028 6012
rect 8010 6012 8028 6030
rect 8010 6030 8028 6048
rect 8010 6048 8028 6066
rect 8010 6066 8028 6084
rect 8010 6084 8028 6102
rect 8010 6102 8028 6120
rect 8010 6120 8028 6138
rect 8010 6138 8028 6156
rect 8010 6156 8028 6174
rect 8010 6174 8028 6192
rect 8010 6192 8028 6210
rect 8010 6210 8028 6228
rect 8010 6228 8028 6246
rect 8010 6246 8028 6264
rect 8010 6264 8028 6282
rect 8010 6282 8028 6300
rect 8010 6300 8028 6318
rect 8010 6318 8028 6336
rect 8010 6336 8028 6354
rect 8010 6354 8028 6372
rect 8010 6372 8028 6390
rect 8010 6390 8028 6408
rect 8010 6408 8028 6426
rect 8010 6426 8028 6444
rect 8010 6444 8028 6462
rect 8010 6462 8028 6480
rect 8010 6480 8028 6498
rect 8010 6498 8028 6516
rect 8010 6516 8028 6534
rect 8010 6534 8028 6552
rect 8010 6552 8028 6570
rect 8010 6570 8028 6588
rect 8010 6588 8028 6606
rect 8010 6606 8028 6624
rect 8010 6624 8028 6642
rect 8010 6642 8028 6660
rect 8010 6660 8028 6678
rect 8010 6678 8028 6696
rect 8010 6696 8028 6714
rect 8010 6714 8028 6732
rect 8010 6732 8028 6750
rect 8010 6750 8028 6768
rect 8010 6768 8028 6786
rect 8010 6786 8028 6804
rect 8010 6804 8028 6822
rect 8010 6822 8028 6840
rect 8010 6840 8028 6858
rect 8010 6858 8028 6876
rect 8010 6876 8028 6894
rect 8010 6894 8028 6912
rect 8010 6912 8028 6930
rect 8010 6930 8028 6948
rect 8010 6948 8028 6966
rect 8010 6966 8028 6984
rect 8010 6984 8028 7002
rect 8010 7002 8028 7020
rect 8010 7020 8028 7038
rect 8028 2430 8046 2448
rect 8028 2448 8046 2466
rect 8028 2466 8046 2484
rect 8028 2484 8046 2502
rect 8028 2502 8046 2520
rect 8028 2520 8046 2538
rect 8028 2538 8046 2556
rect 8028 2556 8046 2574
rect 8028 2574 8046 2592
rect 8028 2592 8046 2610
rect 8028 2610 8046 2628
rect 8028 2628 8046 2646
rect 8028 2646 8046 2664
rect 8028 2664 8046 2682
rect 8028 2682 8046 2700
rect 8028 2700 8046 2718
rect 8028 2718 8046 2736
rect 8028 2736 8046 2754
rect 8028 2754 8046 2772
rect 8028 2772 8046 2790
rect 8028 2790 8046 2808
rect 8028 2808 8046 2826
rect 8028 2826 8046 2844
rect 8028 2844 8046 2862
rect 8028 2862 8046 2880
rect 8028 2880 8046 2898
rect 8028 2898 8046 2916
rect 8028 2916 8046 2934
rect 8028 2934 8046 2952
rect 8028 2952 8046 2970
rect 8028 2970 8046 2988
rect 8028 2988 8046 3006
rect 8028 3006 8046 3024
rect 8028 3024 8046 3042
rect 8028 3042 8046 3060
rect 8028 3060 8046 3078
rect 8028 3078 8046 3096
rect 8028 3096 8046 3114
rect 8028 3114 8046 3132
rect 8028 3132 8046 3150
rect 8028 3150 8046 3168
rect 8028 3168 8046 3186
rect 8028 3186 8046 3204
rect 8028 3204 8046 3222
rect 8028 3222 8046 3240
rect 8028 3240 8046 3258
rect 8028 3258 8046 3276
rect 8028 3276 8046 3294
rect 8028 3294 8046 3312
rect 8028 3312 8046 3330
rect 8028 3330 8046 3348
rect 8028 3348 8046 3366
rect 8028 5310 8046 5328
rect 8028 5328 8046 5346
rect 8028 5346 8046 5364
rect 8028 5364 8046 5382
rect 8028 5382 8046 5400
rect 8028 5400 8046 5418
rect 8028 5418 8046 5436
rect 8028 5436 8046 5454
rect 8028 5454 8046 5472
rect 8028 5472 8046 5490
rect 8028 5490 8046 5508
rect 8028 5508 8046 5526
rect 8028 5526 8046 5544
rect 8028 5544 8046 5562
rect 8028 5562 8046 5580
rect 8028 5580 8046 5598
rect 8028 5598 8046 5616
rect 8028 5616 8046 5634
rect 8028 5634 8046 5652
rect 8028 5652 8046 5670
rect 8028 5670 8046 5688
rect 8028 5688 8046 5706
rect 8028 5706 8046 5724
rect 8028 5724 8046 5742
rect 8028 5742 8046 5760
rect 8028 5760 8046 5778
rect 8028 5778 8046 5796
rect 8028 5796 8046 5814
rect 8028 5814 8046 5832
rect 8028 5832 8046 5850
rect 8028 5850 8046 5868
rect 8028 5868 8046 5886
rect 8028 5886 8046 5904
rect 8028 5904 8046 5922
rect 8028 5922 8046 5940
rect 8028 5940 8046 5958
rect 8028 5958 8046 5976
rect 8028 5976 8046 5994
rect 8028 5994 8046 6012
rect 8028 6012 8046 6030
rect 8028 6030 8046 6048
rect 8028 6048 8046 6066
rect 8028 6066 8046 6084
rect 8028 6084 8046 6102
rect 8028 6102 8046 6120
rect 8028 6120 8046 6138
rect 8028 6138 8046 6156
rect 8028 6156 8046 6174
rect 8028 6174 8046 6192
rect 8028 6192 8046 6210
rect 8028 6210 8046 6228
rect 8028 6228 8046 6246
rect 8028 6246 8046 6264
rect 8028 6264 8046 6282
rect 8028 6282 8046 6300
rect 8028 6300 8046 6318
rect 8028 6318 8046 6336
rect 8028 6336 8046 6354
rect 8028 6354 8046 6372
rect 8028 6372 8046 6390
rect 8028 6390 8046 6408
rect 8028 6408 8046 6426
rect 8028 6426 8046 6444
rect 8028 6444 8046 6462
rect 8028 6462 8046 6480
rect 8028 6480 8046 6498
rect 8028 6498 8046 6516
rect 8028 6516 8046 6534
rect 8028 6534 8046 6552
rect 8028 6552 8046 6570
rect 8028 6570 8046 6588
rect 8028 6588 8046 6606
rect 8028 6606 8046 6624
rect 8028 6624 8046 6642
rect 8028 6642 8046 6660
rect 8028 6660 8046 6678
rect 8028 6678 8046 6696
rect 8028 6696 8046 6714
rect 8028 6714 8046 6732
rect 8028 6732 8046 6750
rect 8028 6750 8046 6768
rect 8028 6768 8046 6786
rect 8028 6786 8046 6804
rect 8028 6804 8046 6822
rect 8028 6822 8046 6840
rect 8028 6840 8046 6858
rect 8028 6858 8046 6876
rect 8028 6876 8046 6894
rect 8028 6894 8046 6912
rect 8028 6912 8046 6930
rect 8028 6930 8046 6948
rect 8028 6948 8046 6966
rect 8028 6966 8046 6984
rect 8028 6984 8046 7002
rect 8028 7002 8046 7020
rect 8028 7020 8046 7038
rect 8046 2430 8064 2448
rect 8046 2448 8064 2466
rect 8046 2466 8064 2484
rect 8046 2484 8064 2502
rect 8046 2502 8064 2520
rect 8046 2520 8064 2538
rect 8046 2538 8064 2556
rect 8046 2556 8064 2574
rect 8046 2574 8064 2592
rect 8046 2592 8064 2610
rect 8046 2610 8064 2628
rect 8046 2628 8064 2646
rect 8046 2646 8064 2664
rect 8046 2664 8064 2682
rect 8046 2682 8064 2700
rect 8046 2700 8064 2718
rect 8046 2718 8064 2736
rect 8046 2736 8064 2754
rect 8046 2754 8064 2772
rect 8046 2772 8064 2790
rect 8046 2790 8064 2808
rect 8046 2808 8064 2826
rect 8046 2826 8064 2844
rect 8046 2844 8064 2862
rect 8046 2862 8064 2880
rect 8046 2880 8064 2898
rect 8046 2898 8064 2916
rect 8046 2916 8064 2934
rect 8046 2934 8064 2952
rect 8046 2952 8064 2970
rect 8046 2970 8064 2988
rect 8046 2988 8064 3006
rect 8046 3006 8064 3024
rect 8046 3024 8064 3042
rect 8046 3042 8064 3060
rect 8046 3060 8064 3078
rect 8046 3078 8064 3096
rect 8046 3096 8064 3114
rect 8046 3114 8064 3132
rect 8046 3132 8064 3150
rect 8046 3150 8064 3168
rect 8046 3168 8064 3186
rect 8046 3186 8064 3204
rect 8046 3204 8064 3222
rect 8046 3222 8064 3240
rect 8046 3240 8064 3258
rect 8046 3258 8064 3276
rect 8046 3276 8064 3294
rect 8046 3294 8064 3312
rect 8046 3312 8064 3330
rect 8046 3330 8064 3348
rect 8046 3348 8064 3366
rect 8046 3366 8064 3384
rect 8046 5328 8064 5346
rect 8046 5346 8064 5364
rect 8046 5364 8064 5382
rect 8046 5382 8064 5400
rect 8046 5400 8064 5418
rect 8046 5418 8064 5436
rect 8046 5436 8064 5454
rect 8046 5454 8064 5472
rect 8046 5472 8064 5490
rect 8046 5490 8064 5508
rect 8046 5508 8064 5526
rect 8046 5526 8064 5544
rect 8046 5544 8064 5562
rect 8046 5562 8064 5580
rect 8046 5580 8064 5598
rect 8046 5598 8064 5616
rect 8046 5616 8064 5634
rect 8046 5634 8064 5652
rect 8046 5652 8064 5670
rect 8046 5670 8064 5688
rect 8046 5688 8064 5706
rect 8046 5706 8064 5724
rect 8046 5724 8064 5742
rect 8046 5742 8064 5760
rect 8046 5760 8064 5778
rect 8046 5778 8064 5796
rect 8046 5796 8064 5814
rect 8046 5814 8064 5832
rect 8046 5832 8064 5850
rect 8046 5850 8064 5868
rect 8046 5868 8064 5886
rect 8046 5886 8064 5904
rect 8046 5904 8064 5922
rect 8046 5922 8064 5940
rect 8046 5940 8064 5958
rect 8046 5958 8064 5976
rect 8046 5976 8064 5994
rect 8046 5994 8064 6012
rect 8046 6012 8064 6030
rect 8046 6030 8064 6048
rect 8046 6048 8064 6066
rect 8046 6066 8064 6084
rect 8046 6084 8064 6102
rect 8046 6102 8064 6120
rect 8046 6120 8064 6138
rect 8046 6138 8064 6156
rect 8046 6156 8064 6174
rect 8046 6174 8064 6192
rect 8046 6192 8064 6210
rect 8046 6210 8064 6228
rect 8046 6228 8064 6246
rect 8046 6246 8064 6264
rect 8046 6264 8064 6282
rect 8046 6282 8064 6300
rect 8046 6300 8064 6318
rect 8046 6318 8064 6336
rect 8046 6336 8064 6354
rect 8046 6354 8064 6372
rect 8046 6372 8064 6390
rect 8046 6390 8064 6408
rect 8046 6408 8064 6426
rect 8046 6426 8064 6444
rect 8046 6444 8064 6462
rect 8046 6462 8064 6480
rect 8046 6480 8064 6498
rect 8046 6498 8064 6516
rect 8046 6516 8064 6534
rect 8046 6534 8064 6552
rect 8046 6552 8064 6570
rect 8046 6570 8064 6588
rect 8046 6588 8064 6606
rect 8046 6606 8064 6624
rect 8046 6624 8064 6642
rect 8046 6642 8064 6660
rect 8046 6660 8064 6678
rect 8046 6678 8064 6696
rect 8046 6696 8064 6714
rect 8046 6714 8064 6732
rect 8046 6732 8064 6750
rect 8046 6750 8064 6768
rect 8046 6768 8064 6786
rect 8046 6786 8064 6804
rect 8046 6804 8064 6822
rect 8046 6822 8064 6840
rect 8046 6840 8064 6858
rect 8046 6858 8064 6876
rect 8046 6876 8064 6894
rect 8046 6894 8064 6912
rect 8046 6912 8064 6930
rect 8046 6930 8064 6948
rect 8046 6948 8064 6966
rect 8046 6966 8064 6984
rect 8046 6984 8064 7002
rect 8046 7002 8064 7020
rect 8046 7020 8064 7038
rect 8046 7038 8064 7056
rect 8064 2448 8082 2466
rect 8064 2466 8082 2484
rect 8064 2484 8082 2502
rect 8064 2502 8082 2520
rect 8064 2520 8082 2538
rect 8064 2538 8082 2556
rect 8064 2556 8082 2574
rect 8064 2574 8082 2592
rect 8064 2592 8082 2610
rect 8064 2610 8082 2628
rect 8064 2628 8082 2646
rect 8064 2646 8082 2664
rect 8064 2664 8082 2682
rect 8064 2682 8082 2700
rect 8064 2700 8082 2718
rect 8064 2718 8082 2736
rect 8064 2736 8082 2754
rect 8064 2754 8082 2772
rect 8064 2772 8082 2790
rect 8064 2790 8082 2808
rect 8064 2808 8082 2826
rect 8064 2826 8082 2844
rect 8064 2844 8082 2862
rect 8064 2862 8082 2880
rect 8064 2880 8082 2898
rect 8064 2898 8082 2916
rect 8064 2916 8082 2934
rect 8064 2934 8082 2952
rect 8064 2952 8082 2970
rect 8064 2970 8082 2988
rect 8064 2988 8082 3006
rect 8064 3006 8082 3024
rect 8064 3024 8082 3042
rect 8064 3042 8082 3060
rect 8064 3060 8082 3078
rect 8064 3078 8082 3096
rect 8064 3096 8082 3114
rect 8064 3114 8082 3132
rect 8064 3132 8082 3150
rect 8064 3150 8082 3168
rect 8064 3168 8082 3186
rect 8064 3186 8082 3204
rect 8064 3204 8082 3222
rect 8064 3222 8082 3240
rect 8064 3240 8082 3258
rect 8064 3258 8082 3276
rect 8064 3276 8082 3294
rect 8064 3294 8082 3312
rect 8064 3312 8082 3330
rect 8064 3330 8082 3348
rect 8064 3348 8082 3366
rect 8064 3366 8082 3384
rect 8064 5346 8082 5364
rect 8064 5364 8082 5382
rect 8064 5382 8082 5400
rect 8064 5400 8082 5418
rect 8064 5418 8082 5436
rect 8064 5436 8082 5454
rect 8064 5454 8082 5472
rect 8064 5472 8082 5490
rect 8064 5490 8082 5508
rect 8064 5508 8082 5526
rect 8064 5526 8082 5544
rect 8064 5544 8082 5562
rect 8064 5562 8082 5580
rect 8064 5580 8082 5598
rect 8064 5598 8082 5616
rect 8064 5616 8082 5634
rect 8064 5634 8082 5652
rect 8064 5652 8082 5670
rect 8064 5670 8082 5688
rect 8064 5688 8082 5706
rect 8064 5706 8082 5724
rect 8064 5724 8082 5742
rect 8064 5742 8082 5760
rect 8064 5760 8082 5778
rect 8064 5778 8082 5796
rect 8064 5796 8082 5814
rect 8064 5814 8082 5832
rect 8064 5832 8082 5850
rect 8064 5850 8082 5868
rect 8064 5868 8082 5886
rect 8064 5886 8082 5904
rect 8064 5904 8082 5922
rect 8064 5922 8082 5940
rect 8064 5940 8082 5958
rect 8064 5958 8082 5976
rect 8064 5976 8082 5994
rect 8064 5994 8082 6012
rect 8064 6012 8082 6030
rect 8064 6030 8082 6048
rect 8064 6048 8082 6066
rect 8064 6066 8082 6084
rect 8064 6084 8082 6102
rect 8064 6102 8082 6120
rect 8064 6120 8082 6138
rect 8064 6138 8082 6156
rect 8064 6156 8082 6174
rect 8064 6174 8082 6192
rect 8064 6192 8082 6210
rect 8064 6210 8082 6228
rect 8064 6228 8082 6246
rect 8064 6246 8082 6264
rect 8064 6264 8082 6282
rect 8064 6282 8082 6300
rect 8064 6300 8082 6318
rect 8064 6318 8082 6336
rect 8064 6336 8082 6354
rect 8064 6354 8082 6372
rect 8064 6372 8082 6390
rect 8064 6390 8082 6408
rect 8064 6408 8082 6426
rect 8064 6426 8082 6444
rect 8064 6444 8082 6462
rect 8064 6462 8082 6480
rect 8064 6480 8082 6498
rect 8064 6498 8082 6516
rect 8064 6516 8082 6534
rect 8064 6534 8082 6552
rect 8064 6552 8082 6570
rect 8064 6570 8082 6588
rect 8064 6588 8082 6606
rect 8064 6606 8082 6624
rect 8064 6624 8082 6642
rect 8064 6642 8082 6660
rect 8064 6660 8082 6678
rect 8064 6678 8082 6696
rect 8064 6696 8082 6714
rect 8064 6714 8082 6732
rect 8064 6732 8082 6750
rect 8064 6750 8082 6768
rect 8064 6768 8082 6786
rect 8064 6786 8082 6804
rect 8064 6804 8082 6822
rect 8064 6822 8082 6840
rect 8064 6840 8082 6858
rect 8064 6858 8082 6876
rect 8064 6876 8082 6894
rect 8064 6894 8082 6912
rect 8064 6912 8082 6930
rect 8064 6930 8082 6948
rect 8064 6948 8082 6966
rect 8064 6966 8082 6984
rect 8064 6984 8082 7002
rect 8064 7002 8082 7020
rect 8064 7020 8082 7038
rect 8064 7038 8082 7056
rect 8064 7056 8082 7074
rect 8082 2466 8100 2484
rect 8082 2484 8100 2502
rect 8082 2502 8100 2520
rect 8082 2520 8100 2538
rect 8082 2538 8100 2556
rect 8082 2556 8100 2574
rect 8082 2574 8100 2592
rect 8082 2592 8100 2610
rect 8082 2610 8100 2628
rect 8082 2628 8100 2646
rect 8082 2646 8100 2664
rect 8082 2664 8100 2682
rect 8082 2682 8100 2700
rect 8082 2700 8100 2718
rect 8082 2718 8100 2736
rect 8082 2736 8100 2754
rect 8082 2754 8100 2772
rect 8082 2772 8100 2790
rect 8082 2790 8100 2808
rect 8082 2808 8100 2826
rect 8082 2826 8100 2844
rect 8082 2844 8100 2862
rect 8082 2862 8100 2880
rect 8082 2880 8100 2898
rect 8082 2898 8100 2916
rect 8082 2916 8100 2934
rect 8082 2934 8100 2952
rect 8082 2952 8100 2970
rect 8082 2970 8100 2988
rect 8082 2988 8100 3006
rect 8082 3006 8100 3024
rect 8082 3024 8100 3042
rect 8082 3042 8100 3060
rect 8082 3060 8100 3078
rect 8082 3078 8100 3096
rect 8082 3096 8100 3114
rect 8082 3114 8100 3132
rect 8082 3132 8100 3150
rect 8082 3150 8100 3168
rect 8082 3168 8100 3186
rect 8082 3186 8100 3204
rect 8082 3204 8100 3222
rect 8082 3222 8100 3240
rect 8082 3240 8100 3258
rect 8082 3258 8100 3276
rect 8082 3276 8100 3294
rect 8082 3294 8100 3312
rect 8082 3312 8100 3330
rect 8082 3330 8100 3348
rect 8082 3348 8100 3366
rect 8082 3366 8100 3384
rect 8082 5382 8100 5400
rect 8082 5400 8100 5418
rect 8082 5418 8100 5436
rect 8082 5436 8100 5454
rect 8082 5454 8100 5472
rect 8082 5472 8100 5490
rect 8082 5490 8100 5508
rect 8082 5508 8100 5526
rect 8082 5526 8100 5544
rect 8082 5544 8100 5562
rect 8082 5562 8100 5580
rect 8082 5580 8100 5598
rect 8082 5598 8100 5616
rect 8082 5616 8100 5634
rect 8082 5634 8100 5652
rect 8082 5652 8100 5670
rect 8082 5670 8100 5688
rect 8082 5688 8100 5706
rect 8082 5706 8100 5724
rect 8082 5724 8100 5742
rect 8082 5742 8100 5760
rect 8082 5760 8100 5778
rect 8082 5778 8100 5796
rect 8082 5796 8100 5814
rect 8082 5814 8100 5832
rect 8082 5832 8100 5850
rect 8082 5850 8100 5868
rect 8082 5868 8100 5886
rect 8082 5886 8100 5904
rect 8082 5904 8100 5922
rect 8082 5922 8100 5940
rect 8082 5940 8100 5958
rect 8082 5958 8100 5976
rect 8082 5976 8100 5994
rect 8082 5994 8100 6012
rect 8082 6012 8100 6030
rect 8082 6030 8100 6048
rect 8082 6048 8100 6066
rect 8082 6066 8100 6084
rect 8082 6084 8100 6102
rect 8082 6102 8100 6120
rect 8082 6120 8100 6138
rect 8082 6138 8100 6156
rect 8082 6156 8100 6174
rect 8082 6174 8100 6192
rect 8082 6192 8100 6210
rect 8082 6210 8100 6228
rect 8082 6228 8100 6246
rect 8082 6246 8100 6264
rect 8082 6264 8100 6282
rect 8082 6282 8100 6300
rect 8082 6300 8100 6318
rect 8082 6318 8100 6336
rect 8082 6336 8100 6354
rect 8082 6354 8100 6372
rect 8082 6372 8100 6390
rect 8082 6390 8100 6408
rect 8082 6408 8100 6426
rect 8082 6426 8100 6444
rect 8082 6444 8100 6462
rect 8082 6462 8100 6480
rect 8082 6480 8100 6498
rect 8082 6498 8100 6516
rect 8082 6516 8100 6534
rect 8082 6534 8100 6552
rect 8082 6552 8100 6570
rect 8082 6570 8100 6588
rect 8082 6588 8100 6606
rect 8082 6606 8100 6624
rect 8082 6624 8100 6642
rect 8082 6642 8100 6660
rect 8082 6660 8100 6678
rect 8082 6678 8100 6696
rect 8082 6696 8100 6714
rect 8082 6714 8100 6732
rect 8082 6732 8100 6750
rect 8082 6750 8100 6768
rect 8082 6768 8100 6786
rect 8082 6786 8100 6804
rect 8082 6804 8100 6822
rect 8082 6822 8100 6840
rect 8082 6840 8100 6858
rect 8082 6858 8100 6876
rect 8082 6876 8100 6894
rect 8082 6894 8100 6912
rect 8082 6912 8100 6930
rect 8082 6930 8100 6948
rect 8082 6948 8100 6966
rect 8082 6966 8100 6984
rect 8082 6984 8100 7002
rect 8082 7002 8100 7020
rect 8082 7020 8100 7038
rect 8082 7038 8100 7056
rect 8082 7056 8100 7074
rect 8100 2484 8118 2502
rect 8100 2502 8118 2520
rect 8100 2520 8118 2538
rect 8100 2538 8118 2556
rect 8100 2556 8118 2574
rect 8100 2574 8118 2592
rect 8100 2592 8118 2610
rect 8100 2610 8118 2628
rect 8100 2628 8118 2646
rect 8100 2646 8118 2664
rect 8100 2664 8118 2682
rect 8100 2682 8118 2700
rect 8100 2700 8118 2718
rect 8100 2718 8118 2736
rect 8100 2736 8118 2754
rect 8100 2754 8118 2772
rect 8100 2772 8118 2790
rect 8100 2790 8118 2808
rect 8100 2808 8118 2826
rect 8100 2826 8118 2844
rect 8100 2844 8118 2862
rect 8100 2862 8118 2880
rect 8100 2880 8118 2898
rect 8100 2898 8118 2916
rect 8100 2916 8118 2934
rect 8100 2934 8118 2952
rect 8100 2952 8118 2970
rect 8100 2970 8118 2988
rect 8100 2988 8118 3006
rect 8100 3006 8118 3024
rect 8100 3024 8118 3042
rect 8100 3042 8118 3060
rect 8100 3060 8118 3078
rect 8100 3078 8118 3096
rect 8100 3096 8118 3114
rect 8100 3114 8118 3132
rect 8100 3132 8118 3150
rect 8100 3150 8118 3168
rect 8100 3168 8118 3186
rect 8100 3186 8118 3204
rect 8100 3204 8118 3222
rect 8100 3222 8118 3240
rect 8100 3240 8118 3258
rect 8100 3258 8118 3276
rect 8100 3276 8118 3294
rect 8100 3294 8118 3312
rect 8100 3312 8118 3330
rect 8100 3330 8118 3348
rect 8100 3348 8118 3366
rect 8100 3366 8118 3384
rect 8100 5400 8118 5418
rect 8100 5418 8118 5436
rect 8100 5436 8118 5454
rect 8100 5454 8118 5472
rect 8100 5472 8118 5490
rect 8100 5490 8118 5508
rect 8100 5508 8118 5526
rect 8100 5526 8118 5544
rect 8100 5544 8118 5562
rect 8100 5562 8118 5580
rect 8100 5580 8118 5598
rect 8100 5598 8118 5616
rect 8100 5616 8118 5634
rect 8100 5634 8118 5652
rect 8100 5652 8118 5670
rect 8100 5670 8118 5688
rect 8100 5688 8118 5706
rect 8100 5706 8118 5724
rect 8100 5724 8118 5742
rect 8100 5742 8118 5760
rect 8100 5760 8118 5778
rect 8100 5778 8118 5796
rect 8100 5796 8118 5814
rect 8100 5814 8118 5832
rect 8100 5832 8118 5850
rect 8100 5850 8118 5868
rect 8100 5868 8118 5886
rect 8100 5886 8118 5904
rect 8100 5904 8118 5922
rect 8100 5922 8118 5940
rect 8100 5940 8118 5958
rect 8100 5958 8118 5976
rect 8100 5976 8118 5994
rect 8100 5994 8118 6012
rect 8100 6012 8118 6030
rect 8100 6030 8118 6048
rect 8100 6048 8118 6066
rect 8100 6066 8118 6084
rect 8100 6084 8118 6102
rect 8100 6102 8118 6120
rect 8100 6120 8118 6138
rect 8100 6138 8118 6156
rect 8100 6156 8118 6174
rect 8100 6174 8118 6192
rect 8100 6192 8118 6210
rect 8100 6210 8118 6228
rect 8100 6228 8118 6246
rect 8100 6246 8118 6264
rect 8100 6264 8118 6282
rect 8100 6282 8118 6300
rect 8100 6300 8118 6318
rect 8100 6318 8118 6336
rect 8100 6336 8118 6354
rect 8100 6354 8118 6372
rect 8100 6372 8118 6390
rect 8100 6390 8118 6408
rect 8100 6408 8118 6426
rect 8100 6426 8118 6444
rect 8100 6444 8118 6462
rect 8100 6462 8118 6480
rect 8100 6480 8118 6498
rect 8100 6498 8118 6516
rect 8100 6516 8118 6534
rect 8100 6534 8118 6552
rect 8100 6552 8118 6570
rect 8100 6570 8118 6588
rect 8100 6588 8118 6606
rect 8100 6606 8118 6624
rect 8100 6624 8118 6642
rect 8100 6642 8118 6660
rect 8100 6660 8118 6678
rect 8100 6678 8118 6696
rect 8100 6696 8118 6714
rect 8100 6714 8118 6732
rect 8100 6732 8118 6750
rect 8100 6750 8118 6768
rect 8100 6768 8118 6786
rect 8100 6786 8118 6804
rect 8100 6804 8118 6822
rect 8100 6822 8118 6840
rect 8100 6840 8118 6858
rect 8100 6858 8118 6876
rect 8100 6876 8118 6894
rect 8100 6894 8118 6912
rect 8100 6912 8118 6930
rect 8100 6930 8118 6948
rect 8100 6948 8118 6966
rect 8100 6966 8118 6984
rect 8100 6984 8118 7002
rect 8100 7002 8118 7020
rect 8100 7020 8118 7038
rect 8100 7038 8118 7056
rect 8100 7056 8118 7074
rect 8100 7074 8118 7092
rect 8118 2484 8136 2502
rect 8118 2502 8136 2520
rect 8118 2520 8136 2538
rect 8118 2538 8136 2556
rect 8118 2556 8136 2574
rect 8118 2574 8136 2592
rect 8118 2592 8136 2610
rect 8118 2610 8136 2628
rect 8118 2628 8136 2646
rect 8118 2646 8136 2664
rect 8118 2664 8136 2682
rect 8118 2682 8136 2700
rect 8118 2700 8136 2718
rect 8118 2718 8136 2736
rect 8118 2736 8136 2754
rect 8118 2754 8136 2772
rect 8118 2772 8136 2790
rect 8118 2790 8136 2808
rect 8118 2808 8136 2826
rect 8118 2826 8136 2844
rect 8118 2844 8136 2862
rect 8118 2862 8136 2880
rect 8118 2880 8136 2898
rect 8118 2898 8136 2916
rect 8118 2916 8136 2934
rect 8118 2934 8136 2952
rect 8118 2952 8136 2970
rect 8118 2970 8136 2988
rect 8118 2988 8136 3006
rect 8118 3006 8136 3024
rect 8118 3024 8136 3042
rect 8118 3042 8136 3060
rect 8118 3060 8136 3078
rect 8118 3078 8136 3096
rect 8118 3096 8136 3114
rect 8118 3114 8136 3132
rect 8118 3132 8136 3150
rect 8118 3150 8136 3168
rect 8118 3168 8136 3186
rect 8118 3186 8136 3204
rect 8118 3204 8136 3222
rect 8118 3222 8136 3240
rect 8118 3240 8136 3258
rect 8118 3258 8136 3276
rect 8118 3276 8136 3294
rect 8118 3294 8136 3312
rect 8118 3312 8136 3330
rect 8118 3330 8136 3348
rect 8118 3348 8136 3366
rect 8118 3366 8136 3384
rect 8118 3384 8136 3402
rect 8118 5418 8136 5436
rect 8118 5436 8136 5454
rect 8118 5454 8136 5472
rect 8118 5472 8136 5490
rect 8118 5490 8136 5508
rect 8118 5508 8136 5526
rect 8118 5526 8136 5544
rect 8118 5544 8136 5562
rect 8118 5562 8136 5580
rect 8118 5580 8136 5598
rect 8118 5598 8136 5616
rect 8118 5616 8136 5634
rect 8118 5634 8136 5652
rect 8118 5652 8136 5670
rect 8118 5670 8136 5688
rect 8118 5688 8136 5706
rect 8118 5706 8136 5724
rect 8118 5724 8136 5742
rect 8118 5742 8136 5760
rect 8118 5760 8136 5778
rect 8118 5778 8136 5796
rect 8118 5796 8136 5814
rect 8118 5814 8136 5832
rect 8118 5832 8136 5850
rect 8118 5850 8136 5868
rect 8118 5868 8136 5886
rect 8118 5886 8136 5904
rect 8118 5904 8136 5922
rect 8118 5922 8136 5940
rect 8118 5940 8136 5958
rect 8118 5958 8136 5976
rect 8118 5976 8136 5994
rect 8118 5994 8136 6012
rect 8118 6012 8136 6030
rect 8118 6030 8136 6048
rect 8118 6048 8136 6066
rect 8118 6066 8136 6084
rect 8118 6084 8136 6102
rect 8118 6102 8136 6120
rect 8118 6120 8136 6138
rect 8118 6138 8136 6156
rect 8118 6156 8136 6174
rect 8118 6174 8136 6192
rect 8118 6192 8136 6210
rect 8118 6210 8136 6228
rect 8118 6228 8136 6246
rect 8118 6246 8136 6264
rect 8118 6264 8136 6282
rect 8118 6282 8136 6300
rect 8118 6300 8136 6318
rect 8118 6318 8136 6336
rect 8118 6336 8136 6354
rect 8118 6354 8136 6372
rect 8118 6372 8136 6390
rect 8118 6390 8136 6408
rect 8118 6408 8136 6426
rect 8118 6426 8136 6444
rect 8118 6444 8136 6462
rect 8118 6462 8136 6480
rect 8118 6480 8136 6498
rect 8118 6498 8136 6516
rect 8118 6516 8136 6534
rect 8118 6534 8136 6552
rect 8118 6552 8136 6570
rect 8118 6570 8136 6588
rect 8118 6588 8136 6606
rect 8118 6606 8136 6624
rect 8118 6624 8136 6642
rect 8118 6642 8136 6660
rect 8118 6660 8136 6678
rect 8118 6678 8136 6696
rect 8118 6696 8136 6714
rect 8118 6714 8136 6732
rect 8118 6732 8136 6750
rect 8118 6750 8136 6768
rect 8118 6768 8136 6786
rect 8118 6786 8136 6804
rect 8118 6804 8136 6822
rect 8118 6822 8136 6840
rect 8118 6840 8136 6858
rect 8118 6858 8136 6876
rect 8118 6876 8136 6894
rect 8118 6894 8136 6912
rect 8118 6912 8136 6930
rect 8118 6930 8136 6948
rect 8118 6948 8136 6966
rect 8118 6966 8136 6984
rect 8118 6984 8136 7002
rect 8118 7002 8136 7020
rect 8118 7020 8136 7038
rect 8118 7038 8136 7056
rect 8118 7056 8136 7074
rect 8118 7074 8136 7092
rect 8118 7092 8136 7110
rect 8136 2502 8154 2520
rect 8136 2520 8154 2538
rect 8136 2538 8154 2556
rect 8136 2556 8154 2574
rect 8136 2574 8154 2592
rect 8136 2592 8154 2610
rect 8136 2610 8154 2628
rect 8136 2628 8154 2646
rect 8136 2646 8154 2664
rect 8136 2664 8154 2682
rect 8136 2682 8154 2700
rect 8136 2700 8154 2718
rect 8136 2718 8154 2736
rect 8136 2736 8154 2754
rect 8136 2754 8154 2772
rect 8136 2772 8154 2790
rect 8136 2790 8154 2808
rect 8136 2808 8154 2826
rect 8136 2826 8154 2844
rect 8136 2844 8154 2862
rect 8136 2862 8154 2880
rect 8136 2880 8154 2898
rect 8136 2898 8154 2916
rect 8136 2916 8154 2934
rect 8136 2934 8154 2952
rect 8136 2952 8154 2970
rect 8136 2970 8154 2988
rect 8136 2988 8154 3006
rect 8136 3006 8154 3024
rect 8136 3024 8154 3042
rect 8136 3042 8154 3060
rect 8136 3060 8154 3078
rect 8136 3078 8154 3096
rect 8136 3096 8154 3114
rect 8136 3114 8154 3132
rect 8136 3132 8154 3150
rect 8136 3150 8154 3168
rect 8136 3168 8154 3186
rect 8136 3186 8154 3204
rect 8136 3204 8154 3222
rect 8136 3222 8154 3240
rect 8136 3240 8154 3258
rect 8136 3258 8154 3276
rect 8136 3276 8154 3294
rect 8136 3294 8154 3312
rect 8136 3312 8154 3330
rect 8136 3330 8154 3348
rect 8136 3348 8154 3366
rect 8136 3366 8154 3384
rect 8136 3384 8154 3402
rect 8136 5436 8154 5454
rect 8136 5454 8154 5472
rect 8136 5472 8154 5490
rect 8136 5490 8154 5508
rect 8136 5508 8154 5526
rect 8136 5526 8154 5544
rect 8136 5544 8154 5562
rect 8136 5562 8154 5580
rect 8136 5580 8154 5598
rect 8136 5598 8154 5616
rect 8136 5616 8154 5634
rect 8136 5634 8154 5652
rect 8136 5652 8154 5670
rect 8136 5670 8154 5688
rect 8136 5688 8154 5706
rect 8136 5706 8154 5724
rect 8136 5724 8154 5742
rect 8136 5742 8154 5760
rect 8136 5760 8154 5778
rect 8136 5778 8154 5796
rect 8136 5796 8154 5814
rect 8136 5814 8154 5832
rect 8136 5832 8154 5850
rect 8136 5850 8154 5868
rect 8136 5868 8154 5886
rect 8136 5886 8154 5904
rect 8136 5904 8154 5922
rect 8136 5922 8154 5940
rect 8136 5940 8154 5958
rect 8136 5958 8154 5976
rect 8136 5976 8154 5994
rect 8136 5994 8154 6012
rect 8136 6012 8154 6030
rect 8136 6030 8154 6048
rect 8136 6048 8154 6066
rect 8136 6066 8154 6084
rect 8136 6084 8154 6102
rect 8136 6102 8154 6120
rect 8136 6120 8154 6138
rect 8136 6138 8154 6156
rect 8136 6156 8154 6174
rect 8136 6174 8154 6192
rect 8136 6192 8154 6210
rect 8136 6210 8154 6228
rect 8136 6228 8154 6246
rect 8136 6246 8154 6264
rect 8136 6264 8154 6282
rect 8136 6282 8154 6300
rect 8136 6300 8154 6318
rect 8136 6318 8154 6336
rect 8136 6336 8154 6354
rect 8136 6354 8154 6372
rect 8136 6372 8154 6390
rect 8136 6390 8154 6408
rect 8136 6408 8154 6426
rect 8136 6426 8154 6444
rect 8136 6444 8154 6462
rect 8136 6462 8154 6480
rect 8136 6480 8154 6498
rect 8136 6498 8154 6516
rect 8136 6516 8154 6534
rect 8136 6534 8154 6552
rect 8136 6552 8154 6570
rect 8136 6570 8154 6588
rect 8136 6588 8154 6606
rect 8136 6606 8154 6624
rect 8136 6624 8154 6642
rect 8136 6642 8154 6660
rect 8136 6660 8154 6678
rect 8136 6678 8154 6696
rect 8136 6696 8154 6714
rect 8136 6714 8154 6732
rect 8136 6732 8154 6750
rect 8136 6750 8154 6768
rect 8136 6768 8154 6786
rect 8136 6786 8154 6804
rect 8136 6804 8154 6822
rect 8136 6822 8154 6840
rect 8136 6840 8154 6858
rect 8136 6858 8154 6876
rect 8136 6876 8154 6894
rect 8136 6894 8154 6912
rect 8136 6912 8154 6930
rect 8136 6930 8154 6948
rect 8136 6948 8154 6966
rect 8136 6966 8154 6984
rect 8136 6984 8154 7002
rect 8136 7002 8154 7020
rect 8136 7020 8154 7038
rect 8136 7038 8154 7056
rect 8136 7056 8154 7074
rect 8136 7074 8154 7092
rect 8136 7092 8154 7110
rect 8136 7110 8154 7128
rect 8154 2520 8172 2538
rect 8154 2538 8172 2556
rect 8154 2556 8172 2574
rect 8154 2574 8172 2592
rect 8154 2592 8172 2610
rect 8154 2610 8172 2628
rect 8154 2628 8172 2646
rect 8154 2646 8172 2664
rect 8154 2664 8172 2682
rect 8154 2682 8172 2700
rect 8154 2700 8172 2718
rect 8154 2718 8172 2736
rect 8154 2736 8172 2754
rect 8154 2754 8172 2772
rect 8154 2772 8172 2790
rect 8154 2790 8172 2808
rect 8154 2808 8172 2826
rect 8154 2826 8172 2844
rect 8154 2844 8172 2862
rect 8154 2862 8172 2880
rect 8154 2880 8172 2898
rect 8154 2898 8172 2916
rect 8154 2916 8172 2934
rect 8154 2934 8172 2952
rect 8154 2952 8172 2970
rect 8154 2970 8172 2988
rect 8154 2988 8172 3006
rect 8154 3006 8172 3024
rect 8154 3024 8172 3042
rect 8154 3042 8172 3060
rect 8154 3060 8172 3078
rect 8154 3078 8172 3096
rect 8154 3096 8172 3114
rect 8154 3114 8172 3132
rect 8154 3132 8172 3150
rect 8154 3150 8172 3168
rect 8154 3168 8172 3186
rect 8154 3186 8172 3204
rect 8154 3204 8172 3222
rect 8154 3222 8172 3240
rect 8154 3240 8172 3258
rect 8154 3258 8172 3276
rect 8154 3276 8172 3294
rect 8154 3294 8172 3312
rect 8154 3312 8172 3330
rect 8154 3330 8172 3348
rect 8154 3348 8172 3366
rect 8154 3366 8172 3384
rect 8154 3384 8172 3402
rect 8154 5472 8172 5490
rect 8154 5490 8172 5508
rect 8154 5508 8172 5526
rect 8154 5526 8172 5544
rect 8154 5544 8172 5562
rect 8154 5562 8172 5580
rect 8154 5580 8172 5598
rect 8154 5598 8172 5616
rect 8154 5616 8172 5634
rect 8154 5634 8172 5652
rect 8154 5652 8172 5670
rect 8154 5670 8172 5688
rect 8154 5688 8172 5706
rect 8154 5706 8172 5724
rect 8154 5724 8172 5742
rect 8154 5742 8172 5760
rect 8154 5760 8172 5778
rect 8154 5778 8172 5796
rect 8154 5796 8172 5814
rect 8154 5814 8172 5832
rect 8154 5832 8172 5850
rect 8154 5850 8172 5868
rect 8154 5868 8172 5886
rect 8154 5886 8172 5904
rect 8154 5904 8172 5922
rect 8154 5922 8172 5940
rect 8154 5940 8172 5958
rect 8154 5958 8172 5976
rect 8154 5976 8172 5994
rect 8154 5994 8172 6012
rect 8154 6012 8172 6030
rect 8154 6030 8172 6048
rect 8154 6048 8172 6066
rect 8154 6066 8172 6084
rect 8154 6084 8172 6102
rect 8154 6102 8172 6120
rect 8154 6120 8172 6138
rect 8154 6138 8172 6156
rect 8154 6156 8172 6174
rect 8154 6174 8172 6192
rect 8154 6192 8172 6210
rect 8154 6210 8172 6228
rect 8154 6228 8172 6246
rect 8154 6246 8172 6264
rect 8154 6264 8172 6282
rect 8154 6282 8172 6300
rect 8154 6300 8172 6318
rect 8154 6318 8172 6336
rect 8154 6336 8172 6354
rect 8154 6354 8172 6372
rect 8154 6372 8172 6390
rect 8154 6390 8172 6408
rect 8154 6408 8172 6426
rect 8154 6426 8172 6444
rect 8154 6444 8172 6462
rect 8154 6462 8172 6480
rect 8154 6480 8172 6498
rect 8154 6498 8172 6516
rect 8154 6516 8172 6534
rect 8154 6534 8172 6552
rect 8154 6552 8172 6570
rect 8154 6570 8172 6588
rect 8154 6588 8172 6606
rect 8154 6606 8172 6624
rect 8154 6624 8172 6642
rect 8154 6642 8172 6660
rect 8154 6660 8172 6678
rect 8154 6678 8172 6696
rect 8154 6696 8172 6714
rect 8154 6714 8172 6732
rect 8154 6732 8172 6750
rect 8154 6750 8172 6768
rect 8154 6768 8172 6786
rect 8154 6786 8172 6804
rect 8154 6804 8172 6822
rect 8154 6822 8172 6840
rect 8154 6840 8172 6858
rect 8154 6858 8172 6876
rect 8154 6876 8172 6894
rect 8154 6894 8172 6912
rect 8154 6912 8172 6930
rect 8154 6930 8172 6948
rect 8154 6948 8172 6966
rect 8154 6966 8172 6984
rect 8154 6984 8172 7002
rect 8154 7002 8172 7020
rect 8154 7020 8172 7038
rect 8154 7038 8172 7056
rect 8154 7056 8172 7074
rect 8154 7074 8172 7092
rect 8154 7092 8172 7110
rect 8154 7110 8172 7128
rect 8172 2520 8190 2538
rect 8172 2538 8190 2556
rect 8172 2556 8190 2574
rect 8172 2574 8190 2592
rect 8172 2592 8190 2610
rect 8172 2610 8190 2628
rect 8172 2628 8190 2646
rect 8172 2646 8190 2664
rect 8172 2664 8190 2682
rect 8172 2682 8190 2700
rect 8172 2700 8190 2718
rect 8172 2718 8190 2736
rect 8172 2736 8190 2754
rect 8172 2754 8190 2772
rect 8172 2772 8190 2790
rect 8172 2790 8190 2808
rect 8172 2808 8190 2826
rect 8172 2826 8190 2844
rect 8172 2844 8190 2862
rect 8172 2862 8190 2880
rect 8172 2880 8190 2898
rect 8172 2898 8190 2916
rect 8172 2916 8190 2934
rect 8172 2934 8190 2952
rect 8172 2952 8190 2970
rect 8172 2970 8190 2988
rect 8172 2988 8190 3006
rect 8172 3006 8190 3024
rect 8172 3024 8190 3042
rect 8172 3042 8190 3060
rect 8172 3060 8190 3078
rect 8172 3078 8190 3096
rect 8172 3096 8190 3114
rect 8172 3114 8190 3132
rect 8172 3132 8190 3150
rect 8172 3150 8190 3168
rect 8172 3168 8190 3186
rect 8172 3186 8190 3204
rect 8172 3204 8190 3222
rect 8172 3222 8190 3240
rect 8172 3240 8190 3258
rect 8172 3258 8190 3276
rect 8172 3276 8190 3294
rect 8172 3294 8190 3312
rect 8172 3312 8190 3330
rect 8172 3330 8190 3348
rect 8172 3348 8190 3366
rect 8172 3366 8190 3384
rect 8172 3384 8190 3402
rect 8172 5490 8190 5508
rect 8172 5508 8190 5526
rect 8172 5526 8190 5544
rect 8172 5544 8190 5562
rect 8172 5562 8190 5580
rect 8172 5580 8190 5598
rect 8172 5598 8190 5616
rect 8172 5616 8190 5634
rect 8172 5634 8190 5652
rect 8172 5652 8190 5670
rect 8172 5670 8190 5688
rect 8172 5688 8190 5706
rect 8172 5706 8190 5724
rect 8172 5724 8190 5742
rect 8172 5742 8190 5760
rect 8172 5760 8190 5778
rect 8172 5778 8190 5796
rect 8172 5796 8190 5814
rect 8172 5814 8190 5832
rect 8172 5832 8190 5850
rect 8172 5850 8190 5868
rect 8172 5868 8190 5886
rect 8172 5886 8190 5904
rect 8172 5904 8190 5922
rect 8172 5922 8190 5940
rect 8172 5940 8190 5958
rect 8172 5958 8190 5976
rect 8172 5976 8190 5994
rect 8172 5994 8190 6012
rect 8172 6012 8190 6030
rect 8172 6030 8190 6048
rect 8172 6048 8190 6066
rect 8172 6066 8190 6084
rect 8172 6084 8190 6102
rect 8172 6102 8190 6120
rect 8172 6120 8190 6138
rect 8172 6138 8190 6156
rect 8172 6156 8190 6174
rect 8172 6174 8190 6192
rect 8172 6192 8190 6210
rect 8172 6210 8190 6228
rect 8172 6228 8190 6246
rect 8172 6246 8190 6264
rect 8172 6264 8190 6282
rect 8172 6282 8190 6300
rect 8172 6300 8190 6318
rect 8172 6318 8190 6336
rect 8172 6336 8190 6354
rect 8172 6354 8190 6372
rect 8172 6372 8190 6390
rect 8172 6390 8190 6408
rect 8172 6408 8190 6426
rect 8172 6426 8190 6444
rect 8172 6444 8190 6462
rect 8172 6462 8190 6480
rect 8172 6480 8190 6498
rect 8172 6498 8190 6516
rect 8172 6516 8190 6534
rect 8172 6534 8190 6552
rect 8172 6552 8190 6570
rect 8172 6570 8190 6588
rect 8172 6588 8190 6606
rect 8172 6606 8190 6624
rect 8172 6624 8190 6642
rect 8172 6642 8190 6660
rect 8172 6660 8190 6678
rect 8172 6678 8190 6696
rect 8172 6696 8190 6714
rect 8172 6714 8190 6732
rect 8172 6732 8190 6750
rect 8172 6750 8190 6768
rect 8172 6768 8190 6786
rect 8172 6786 8190 6804
rect 8172 6804 8190 6822
rect 8172 6822 8190 6840
rect 8172 6840 8190 6858
rect 8172 6858 8190 6876
rect 8172 6876 8190 6894
rect 8172 6894 8190 6912
rect 8172 6912 8190 6930
rect 8172 6930 8190 6948
rect 8172 6948 8190 6966
rect 8172 6966 8190 6984
rect 8172 6984 8190 7002
rect 8172 7002 8190 7020
rect 8172 7020 8190 7038
rect 8172 7038 8190 7056
rect 8172 7056 8190 7074
rect 8172 7074 8190 7092
rect 8172 7092 8190 7110
rect 8172 7110 8190 7128
rect 8172 7128 8190 7146
rect 8190 2538 8208 2556
rect 8190 2556 8208 2574
rect 8190 2574 8208 2592
rect 8190 2592 8208 2610
rect 8190 2610 8208 2628
rect 8190 2628 8208 2646
rect 8190 2646 8208 2664
rect 8190 2664 8208 2682
rect 8190 2682 8208 2700
rect 8190 2700 8208 2718
rect 8190 2718 8208 2736
rect 8190 2736 8208 2754
rect 8190 2754 8208 2772
rect 8190 2772 8208 2790
rect 8190 2790 8208 2808
rect 8190 2808 8208 2826
rect 8190 2826 8208 2844
rect 8190 2844 8208 2862
rect 8190 2862 8208 2880
rect 8190 2880 8208 2898
rect 8190 2898 8208 2916
rect 8190 2916 8208 2934
rect 8190 2934 8208 2952
rect 8190 2952 8208 2970
rect 8190 2970 8208 2988
rect 8190 2988 8208 3006
rect 8190 3006 8208 3024
rect 8190 3024 8208 3042
rect 8190 3042 8208 3060
rect 8190 3060 8208 3078
rect 8190 3078 8208 3096
rect 8190 3096 8208 3114
rect 8190 3114 8208 3132
rect 8190 3132 8208 3150
rect 8190 3150 8208 3168
rect 8190 3168 8208 3186
rect 8190 3186 8208 3204
rect 8190 3204 8208 3222
rect 8190 3222 8208 3240
rect 8190 3240 8208 3258
rect 8190 3258 8208 3276
rect 8190 3276 8208 3294
rect 8190 3294 8208 3312
rect 8190 3312 8208 3330
rect 8190 3330 8208 3348
rect 8190 3348 8208 3366
rect 8190 3366 8208 3384
rect 8190 3384 8208 3402
rect 8190 3402 8208 3420
rect 8190 5526 8208 5544
rect 8190 5544 8208 5562
rect 8190 5562 8208 5580
rect 8190 5580 8208 5598
rect 8190 5598 8208 5616
rect 8190 5616 8208 5634
rect 8190 5634 8208 5652
rect 8190 5652 8208 5670
rect 8190 5670 8208 5688
rect 8190 5688 8208 5706
rect 8190 5706 8208 5724
rect 8190 5724 8208 5742
rect 8190 5742 8208 5760
rect 8190 5760 8208 5778
rect 8190 5778 8208 5796
rect 8190 5796 8208 5814
rect 8190 5814 8208 5832
rect 8190 5832 8208 5850
rect 8190 5850 8208 5868
rect 8190 5868 8208 5886
rect 8190 5886 8208 5904
rect 8190 5904 8208 5922
rect 8190 5922 8208 5940
rect 8190 5940 8208 5958
rect 8190 5958 8208 5976
rect 8190 5976 8208 5994
rect 8190 5994 8208 6012
rect 8190 6012 8208 6030
rect 8190 6030 8208 6048
rect 8190 6048 8208 6066
rect 8190 6066 8208 6084
rect 8190 6084 8208 6102
rect 8190 6102 8208 6120
rect 8190 6120 8208 6138
rect 8190 6138 8208 6156
rect 8190 6156 8208 6174
rect 8190 6174 8208 6192
rect 8190 6192 8208 6210
rect 8190 6210 8208 6228
rect 8190 6228 8208 6246
rect 8190 6246 8208 6264
rect 8190 6264 8208 6282
rect 8190 6282 8208 6300
rect 8190 6300 8208 6318
rect 8190 6318 8208 6336
rect 8190 6336 8208 6354
rect 8190 6354 8208 6372
rect 8190 6372 8208 6390
rect 8190 6390 8208 6408
rect 8190 6408 8208 6426
rect 8190 6426 8208 6444
rect 8190 6444 8208 6462
rect 8190 6462 8208 6480
rect 8190 6480 8208 6498
rect 8190 6498 8208 6516
rect 8190 6516 8208 6534
rect 8190 6534 8208 6552
rect 8190 6552 8208 6570
rect 8190 6570 8208 6588
rect 8190 6588 8208 6606
rect 8190 6606 8208 6624
rect 8190 6624 8208 6642
rect 8190 6642 8208 6660
rect 8190 6660 8208 6678
rect 8190 6678 8208 6696
rect 8190 6696 8208 6714
rect 8190 6714 8208 6732
rect 8190 6732 8208 6750
rect 8190 6750 8208 6768
rect 8190 6768 8208 6786
rect 8190 6786 8208 6804
rect 8190 6804 8208 6822
rect 8190 6822 8208 6840
rect 8190 6840 8208 6858
rect 8190 6858 8208 6876
rect 8190 6876 8208 6894
rect 8190 6894 8208 6912
rect 8190 6912 8208 6930
rect 8190 6930 8208 6948
rect 8190 6948 8208 6966
rect 8190 6966 8208 6984
rect 8190 6984 8208 7002
rect 8190 7002 8208 7020
rect 8190 7020 8208 7038
rect 8190 7038 8208 7056
rect 8190 7056 8208 7074
rect 8190 7074 8208 7092
rect 8190 7092 8208 7110
rect 8190 7110 8208 7128
rect 8190 7128 8208 7146
rect 8190 7146 8208 7164
rect 8208 2556 8226 2574
rect 8208 2574 8226 2592
rect 8208 2592 8226 2610
rect 8208 2610 8226 2628
rect 8208 2628 8226 2646
rect 8208 2646 8226 2664
rect 8208 2664 8226 2682
rect 8208 2682 8226 2700
rect 8208 2700 8226 2718
rect 8208 2718 8226 2736
rect 8208 2736 8226 2754
rect 8208 2754 8226 2772
rect 8208 2772 8226 2790
rect 8208 2790 8226 2808
rect 8208 2808 8226 2826
rect 8208 2826 8226 2844
rect 8208 2844 8226 2862
rect 8208 2862 8226 2880
rect 8208 2880 8226 2898
rect 8208 2898 8226 2916
rect 8208 2916 8226 2934
rect 8208 2934 8226 2952
rect 8208 2952 8226 2970
rect 8208 2970 8226 2988
rect 8208 2988 8226 3006
rect 8208 3006 8226 3024
rect 8208 3024 8226 3042
rect 8208 3042 8226 3060
rect 8208 3060 8226 3078
rect 8208 3078 8226 3096
rect 8208 3096 8226 3114
rect 8208 3114 8226 3132
rect 8208 3132 8226 3150
rect 8208 3150 8226 3168
rect 8208 3168 8226 3186
rect 8208 3186 8226 3204
rect 8208 3204 8226 3222
rect 8208 3222 8226 3240
rect 8208 3240 8226 3258
rect 8208 3258 8226 3276
rect 8208 3276 8226 3294
rect 8208 3294 8226 3312
rect 8208 3312 8226 3330
rect 8208 3330 8226 3348
rect 8208 3348 8226 3366
rect 8208 3366 8226 3384
rect 8208 3384 8226 3402
rect 8208 3402 8226 3420
rect 8208 5544 8226 5562
rect 8208 5562 8226 5580
rect 8208 5580 8226 5598
rect 8208 5598 8226 5616
rect 8208 5616 8226 5634
rect 8208 5634 8226 5652
rect 8208 5652 8226 5670
rect 8208 5670 8226 5688
rect 8208 5688 8226 5706
rect 8208 5706 8226 5724
rect 8208 5724 8226 5742
rect 8208 5742 8226 5760
rect 8208 5760 8226 5778
rect 8208 5778 8226 5796
rect 8208 5796 8226 5814
rect 8208 5814 8226 5832
rect 8208 5832 8226 5850
rect 8208 5850 8226 5868
rect 8208 5868 8226 5886
rect 8208 5886 8226 5904
rect 8208 5904 8226 5922
rect 8208 5922 8226 5940
rect 8208 5940 8226 5958
rect 8208 5958 8226 5976
rect 8208 5976 8226 5994
rect 8208 5994 8226 6012
rect 8208 6012 8226 6030
rect 8208 6030 8226 6048
rect 8208 6048 8226 6066
rect 8208 6066 8226 6084
rect 8208 6084 8226 6102
rect 8208 6102 8226 6120
rect 8208 6120 8226 6138
rect 8208 6138 8226 6156
rect 8208 6156 8226 6174
rect 8208 6174 8226 6192
rect 8208 6192 8226 6210
rect 8208 6210 8226 6228
rect 8208 6228 8226 6246
rect 8208 6246 8226 6264
rect 8208 6264 8226 6282
rect 8208 6282 8226 6300
rect 8208 6300 8226 6318
rect 8208 6318 8226 6336
rect 8208 6336 8226 6354
rect 8208 6354 8226 6372
rect 8208 6372 8226 6390
rect 8208 6390 8226 6408
rect 8208 6408 8226 6426
rect 8208 6426 8226 6444
rect 8208 6444 8226 6462
rect 8208 6462 8226 6480
rect 8208 6480 8226 6498
rect 8208 6498 8226 6516
rect 8208 6516 8226 6534
rect 8208 6534 8226 6552
rect 8208 6552 8226 6570
rect 8208 6570 8226 6588
rect 8208 6588 8226 6606
rect 8208 6606 8226 6624
rect 8208 6624 8226 6642
rect 8208 6642 8226 6660
rect 8208 6660 8226 6678
rect 8208 6678 8226 6696
rect 8208 6696 8226 6714
rect 8208 6714 8226 6732
rect 8208 6732 8226 6750
rect 8208 6750 8226 6768
rect 8208 6768 8226 6786
rect 8208 6786 8226 6804
rect 8208 6804 8226 6822
rect 8208 6822 8226 6840
rect 8208 6840 8226 6858
rect 8208 6858 8226 6876
rect 8208 6876 8226 6894
rect 8208 6894 8226 6912
rect 8208 6912 8226 6930
rect 8208 6930 8226 6948
rect 8208 6948 8226 6966
rect 8208 6966 8226 6984
rect 8208 6984 8226 7002
rect 8208 7002 8226 7020
rect 8208 7020 8226 7038
rect 8208 7038 8226 7056
rect 8208 7056 8226 7074
rect 8208 7074 8226 7092
rect 8208 7092 8226 7110
rect 8208 7110 8226 7128
rect 8208 7128 8226 7146
rect 8208 7146 8226 7164
rect 8226 2574 8244 2592
rect 8226 2592 8244 2610
rect 8226 2610 8244 2628
rect 8226 2628 8244 2646
rect 8226 2646 8244 2664
rect 8226 2664 8244 2682
rect 8226 2682 8244 2700
rect 8226 2700 8244 2718
rect 8226 2718 8244 2736
rect 8226 2736 8244 2754
rect 8226 2754 8244 2772
rect 8226 2772 8244 2790
rect 8226 2790 8244 2808
rect 8226 2808 8244 2826
rect 8226 2826 8244 2844
rect 8226 2844 8244 2862
rect 8226 2862 8244 2880
rect 8226 2880 8244 2898
rect 8226 2898 8244 2916
rect 8226 2916 8244 2934
rect 8226 2934 8244 2952
rect 8226 2952 8244 2970
rect 8226 2970 8244 2988
rect 8226 2988 8244 3006
rect 8226 3006 8244 3024
rect 8226 3024 8244 3042
rect 8226 3042 8244 3060
rect 8226 3060 8244 3078
rect 8226 3078 8244 3096
rect 8226 3096 8244 3114
rect 8226 3114 8244 3132
rect 8226 3132 8244 3150
rect 8226 3150 8244 3168
rect 8226 3168 8244 3186
rect 8226 3186 8244 3204
rect 8226 3204 8244 3222
rect 8226 3222 8244 3240
rect 8226 3240 8244 3258
rect 8226 3258 8244 3276
rect 8226 3276 8244 3294
rect 8226 3294 8244 3312
rect 8226 3312 8244 3330
rect 8226 3330 8244 3348
rect 8226 3348 8244 3366
rect 8226 3366 8244 3384
rect 8226 3384 8244 3402
rect 8226 3402 8244 3420
rect 8226 5562 8244 5580
rect 8226 5580 8244 5598
rect 8226 5598 8244 5616
rect 8226 5616 8244 5634
rect 8226 5634 8244 5652
rect 8226 5652 8244 5670
rect 8226 5670 8244 5688
rect 8226 5688 8244 5706
rect 8226 5706 8244 5724
rect 8226 5724 8244 5742
rect 8226 5742 8244 5760
rect 8226 5760 8244 5778
rect 8226 5778 8244 5796
rect 8226 5796 8244 5814
rect 8226 5814 8244 5832
rect 8226 5832 8244 5850
rect 8226 5850 8244 5868
rect 8226 5868 8244 5886
rect 8226 5886 8244 5904
rect 8226 5904 8244 5922
rect 8226 5922 8244 5940
rect 8226 5940 8244 5958
rect 8226 5958 8244 5976
rect 8226 5976 8244 5994
rect 8226 5994 8244 6012
rect 8226 6012 8244 6030
rect 8226 6030 8244 6048
rect 8226 6048 8244 6066
rect 8226 6066 8244 6084
rect 8226 6084 8244 6102
rect 8226 6102 8244 6120
rect 8226 6120 8244 6138
rect 8226 6138 8244 6156
rect 8226 6156 8244 6174
rect 8226 6174 8244 6192
rect 8226 6192 8244 6210
rect 8226 6210 8244 6228
rect 8226 6228 8244 6246
rect 8226 6246 8244 6264
rect 8226 6264 8244 6282
rect 8226 6282 8244 6300
rect 8226 6300 8244 6318
rect 8226 6318 8244 6336
rect 8226 6336 8244 6354
rect 8226 6354 8244 6372
rect 8226 6372 8244 6390
rect 8226 6390 8244 6408
rect 8226 6408 8244 6426
rect 8226 6426 8244 6444
rect 8226 6444 8244 6462
rect 8226 6462 8244 6480
rect 8226 6480 8244 6498
rect 8226 6498 8244 6516
rect 8226 6516 8244 6534
rect 8226 6534 8244 6552
rect 8226 6552 8244 6570
rect 8226 6570 8244 6588
rect 8226 6588 8244 6606
rect 8226 6606 8244 6624
rect 8226 6624 8244 6642
rect 8226 6642 8244 6660
rect 8226 6660 8244 6678
rect 8226 6678 8244 6696
rect 8226 6696 8244 6714
rect 8226 6714 8244 6732
rect 8226 6732 8244 6750
rect 8226 6750 8244 6768
rect 8226 6768 8244 6786
rect 8226 6786 8244 6804
rect 8226 6804 8244 6822
rect 8226 6822 8244 6840
rect 8226 6840 8244 6858
rect 8226 6858 8244 6876
rect 8226 6876 8244 6894
rect 8226 6894 8244 6912
rect 8226 6912 8244 6930
rect 8226 6930 8244 6948
rect 8226 6948 8244 6966
rect 8226 6966 8244 6984
rect 8226 6984 8244 7002
rect 8226 7002 8244 7020
rect 8226 7020 8244 7038
rect 8226 7038 8244 7056
rect 8226 7056 8244 7074
rect 8226 7074 8244 7092
rect 8226 7092 8244 7110
rect 8226 7110 8244 7128
rect 8226 7128 8244 7146
rect 8226 7146 8244 7164
rect 8226 7164 8244 7182
rect 8244 2574 8262 2592
rect 8244 2592 8262 2610
rect 8244 2610 8262 2628
rect 8244 2628 8262 2646
rect 8244 2646 8262 2664
rect 8244 2664 8262 2682
rect 8244 2682 8262 2700
rect 8244 2700 8262 2718
rect 8244 2718 8262 2736
rect 8244 2736 8262 2754
rect 8244 2754 8262 2772
rect 8244 2772 8262 2790
rect 8244 2790 8262 2808
rect 8244 2808 8262 2826
rect 8244 2826 8262 2844
rect 8244 2844 8262 2862
rect 8244 2862 8262 2880
rect 8244 2880 8262 2898
rect 8244 2898 8262 2916
rect 8244 2916 8262 2934
rect 8244 2934 8262 2952
rect 8244 2952 8262 2970
rect 8244 2970 8262 2988
rect 8244 2988 8262 3006
rect 8244 3006 8262 3024
rect 8244 3024 8262 3042
rect 8244 3042 8262 3060
rect 8244 3060 8262 3078
rect 8244 3078 8262 3096
rect 8244 3096 8262 3114
rect 8244 3114 8262 3132
rect 8244 3132 8262 3150
rect 8244 3150 8262 3168
rect 8244 3168 8262 3186
rect 8244 3186 8262 3204
rect 8244 3204 8262 3222
rect 8244 3222 8262 3240
rect 8244 3240 8262 3258
rect 8244 3258 8262 3276
rect 8244 3276 8262 3294
rect 8244 3294 8262 3312
rect 8244 3312 8262 3330
rect 8244 3330 8262 3348
rect 8244 3348 8262 3366
rect 8244 3366 8262 3384
rect 8244 3384 8262 3402
rect 8244 3402 8262 3420
rect 8244 5598 8262 5616
rect 8244 5616 8262 5634
rect 8244 5634 8262 5652
rect 8244 5652 8262 5670
rect 8244 5670 8262 5688
rect 8244 5688 8262 5706
rect 8244 5706 8262 5724
rect 8244 5724 8262 5742
rect 8244 5742 8262 5760
rect 8244 5760 8262 5778
rect 8244 5778 8262 5796
rect 8244 5796 8262 5814
rect 8244 5814 8262 5832
rect 8244 5832 8262 5850
rect 8244 5850 8262 5868
rect 8244 5868 8262 5886
rect 8244 5886 8262 5904
rect 8244 5904 8262 5922
rect 8244 5922 8262 5940
rect 8244 5940 8262 5958
rect 8244 5958 8262 5976
rect 8244 5976 8262 5994
rect 8244 5994 8262 6012
rect 8244 6012 8262 6030
rect 8244 6030 8262 6048
rect 8244 6048 8262 6066
rect 8244 6066 8262 6084
rect 8244 6084 8262 6102
rect 8244 6102 8262 6120
rect 8244 6120 8262 6138
rect 8244 6138 8262 6156
rect 8244 6156 8262 6174
rect 8244 6174 8262 6192
rect 8244 6192 8262 6210
rect 8244 6210 8262 6228
rect 8244 6228 8262 6246
rect 8244 6246 8262 6264
rect 8244 6264 8262 6282
rect 8244 6282 8262 6300
rect 8244 6300 8262 6318
rect 8244 6318 8262 6336
rect 8244 6336 8262 6354
rect 8244 6354 8262 6372
rect 8244 6372 8262 6390
rect 8244 6390 8262 6408
rect 8244 6408 8262 6426
rect 8244 6426 8262 6444
rect 8244 6444 8262 6462
rect 8244 6462 8262 6480
rect 8244 6480 8262 6498
rect 8244 6498 8262 6516
rect 8244 6516 8262 6534
rect 8244 6534 8262 6552
rect 8244 6552 8262 6570
rect 8244 6570 8262 6588
rect 8244 6588 8262 6606
rect 8244 6606 8262 6624
rect 8244 6624 8262 6642
rect 8244 6642 8262 6660
rect 8244 6660 8262 6678
rect 8244 6678 8262 6696
rect 8244 6696 8262 6714
rect 8244 6714 8262 6732
rect 8244 6732 8262 6750
rect 8244 6750 8262 6768
rect 8244 6768 8262 6786
rect 8244 6786 8262 6804
rect 8244 6804 8262 6822
rect 8244 6822 8262 6840
rect 8244 6840 8262 6858
rect 8244 6858 8262 6876
rect 8244 6876 8262 6894
rect 8244 6894 8262 6912
rect 8244 6912 8262 6930
rect 8244 6930 8262 6948
rect 8244 6948 8262 6966
rect 8244 6966 8262 6984
rect 8244 6984 8262 7002
rect 8244 7002 8262 7020
rect 8244 7020 8262 7038
rect 8244 7038 8262 7056
rect 8244 7056 8262 7074
rect 8244 7074 8262 7092
rect 8244 7092 8262 7110
rect 8244 7110 8262 7128
rect 8244 7128 8262 7146
rect 8244 7146 8262 7164
rect 8244 7164 8262 7182
rect 8244 7182 8262 7200
rect 8262 2592 8280 2610
rect 8262 2610 8280 2628
rect 8262 2628 8280 2646
rect 8262 2646 8280 2664
rect 8262 2664 8280 2682
rect 8262 2682 8280 2700
rect 8262 2700 8280 2718
rect 8262 2718 8280 2736
rect 8262 2736 8280 2754
rect 8262 2754 8280 2772
rect 8262 2772 8280 2790
rect 8262 2790 8280 2808
rect 8262 2808 8280 2826
rect 8262 2826 8280 2844
rect 8262 2844 8280 2862
rect 8262 2862 8280 2880
rect 8262 2880 8280 2898
rect 8262 2898 8280 2916
rect 8262 2916 8280 2934
rect 8262 2934 8280 2952
rect 8262 2952 8280 2970
rect 8262 2970 8280 2988
rect 8262 2988 8280 3006
rect 8262 3006 8280 3024
rect 8262 3024 8280 3042
rect 8262 3042 8280 3060
rect 8262 3060 8280 3078
rect 8262 3078 8280 3096
rect 8262 3096 8280 3114
rect 8262 3114 8280 3132
rect 8262 3132 8280 3150
rect 8262 3150 8280 3168
rect 8262 3168 8280 3186
rect 8262 3186 8280 3204
rect 8262 3204 8280 3222
rect 8262 3222 8280 3240
rect 8262 3240 8280 3258
rect 8262 3258 8280 3276
rect 8262 3276 8280 3294
rect 8262 3294 8280 3312
rect 8262 3312 8280 3330
rect 8262 3330 8280 3348
rect 8262 3348 8280 3366
rect 8262 3366 8280 3384
rect 8262 3384 8280 3402
rect 8262 3402 8280 3420
rect 8262 3420 8280 3438
rect 8262 5616 8280 5634
rect 8262 5634 8280 5652
rect 8262 5652 8280 5670
rect 8262 5670 8280 5688
rect 8262 5688 8280 5706
rect 8262 5706 8280 5724
rect 8262 5724 8280 5742
rect 8262 5742 8280 5760
rect 8262 5760 8280 5778
rect 8262 5778 8280 5796
rect 8262 5796 8280 5814
rect 8262 5814 8280 5832
rect 8262 5832 8280 5850
rect 8262 5850 8280 5868
rect 8262 5868 8280 5886
rect 8262 5886 8280 5904
rect 8262 5904 8280 5922
rect 8262 5922 8280 5940
rect 8262 5940 8280 5958
rect 8262 5958 8280 5976
rect 8262 5976 8280 5994
rect 8262 5994 8280 6012
rect 8262 6012 8280 6030
rect 8262 6030 8280 6048
rect 8262 6048 8280 6066
rect 8262 6066 8280 6084
rect 8262 6084 8280 6102
rect 8262 6102 8280 6120
rect 8262 6120 8280 6138
rect 8262 6138 8280 6156
rect 8262 6156 8280 6174
rect 8262 6174 8280 6192
rect 8262 6192 8280 6210
rect 8262 6210 8280 6228
rect 8262 6228 8280 6246
rect 8262 6246 8280 6264
rect 8262 6264 8280 6282
rect 8262 6282 8280 6300
rect 8262 6300 8280 6318
rect 8262 6318 8280 6336
rect 8262 6336 8280 6354
rect 8262 6354 8280 6372
rect 8262 6372 8280 6390
rect 8262 6390 8280 6408
rect 8262 6408 8280 6426
rect 8262 6426 8280 6444
rect 8262 6444 8280 6462
rect 8262 6462 8280 6480
rect 8262 6480 8280 6498
rect 8262 6498 8280 6516
rect 8262 6516 8280 6534
rect 8262 6534 8280 6552
rect 8262 6552 8280 6570
rect 8262 6570 8280 6588
rect 8262 6588 8280 6606
rect 8262 6606 8280 6624
rect 8262 6624 8280 6642
rect 8262 6642 8280 6660
rect 8262 6660 8280 6678
rect 8262 6678 8280 6696
rect 8262 6696 8280 6714
rect 8262 6714 8280 6732
rect 8262 6732 8280 6750
rect 8262 6750 8280 6768
rect 8262 6768 8280 6786
rect 8262 6786 8280 6804
rect 8262 6804 8280 6822
rect 8262 6822 8280 6840
rect 8262 6840 8280 6858
rect 8262 6858 8280 6876
rect 8262 6876 8280 6894
rect 8262 6894 8280 6912
rect 8262 6912 8280 6930
rect 8262 6930 8280 6948
rect 8262 6948 8280 6966
rect 8262 6966 8280 6984
rect 8262 6984 8280 7002
rect 8262 7002 8280 7020
rect 8262 7020 8280 7038
rect 8262 7038 8280 7056
rect 8262 7056 8280 7074
rect 8262 7074 8280 7092
rect 8262 7092 8280 7110
rect 8262 7110 8280 7128
rect 8262 7128 8280 7146
rect 8262 7146 8280 7164
rect 8262 7164 8280 7182
rect 8262 7182 8280 7200
rect 8280 2610 8298 2628
rect 8280 2628 8298 2646
rect 8280 2646 8298 2664
rect 8280 2664 8298 2682
rect 8280 2682 8298 2700
rect 8280 2700 8298 2718
rect 8280 2718 8298 2736
rect 8280 2736 8298 2754
rect 8280 2754 8298 2772
rect 8280 2772 8298 2790
rect 8280 2790 8298 2808
rect 8280 2808 8298 2826
rect 8280 2826 8298 2844
rect 8280 2844 8298 2862
rect 8280 2862 8298 2880
rect 8280 2880 8298 2898
rect 8280 2898 8298 2916
rect 8280 2916 8298 2934
rect 8280 2934 8298 2952
rect 8280 2952 8298 2970
rect 8280 2970 8298 2988
rect 8280 2988 8298 3006
rect 8280 3006 8298 3024
rect 8280 3024 8298 3042
rect 8280 3042 8298 3060
rect 8280 3060 8298 3078
rect 8280 3078 8298 3096
rect 8280 3096 8298 3114
rect 8280 3114 8298 3132
rect 8280 3132 8298 3150
rect 8280 3150 8298 3168
rect 8280 3168 8298 3186
rect 8280 3186 8298 3204
rect 8280 3204 8298 3222
rect 8280 3222 8298 3240
rect 8280 3240 8298 3258
rect 8280 3258 8298 3276
rect 8280 3276 8298 3294
rect 8280 3294 8298 3312
rect 8280 3312 8298 3330
rect 8280 3330 8298 3348
rect 8280 3348 8298 3366
rect 8280 3366 8298 3384
rect 8280 3384 8298 3402
rect 8280 3402 8298 3420
rect 8280 3420 8298 3438
rect 8280 5652 8298 5670
rect 8280 5670 8298 5688
rect 8280 5688 8298 5706
rect 8280 5706 8298 5724
rect 8280 5724 8298 5742
rect 8280 5742 8298 5760
rect 8280 5760 8298 5778
rect 8280 5778 8298 5796
rect 8280 5796 8298 5814
rect 8280 5814 8298 5832
rect 8280 5832 8298 5850
rect 8280 5850 8298 5868
rect 8280 5868 8298 5886
rect 8280 5886 8298 5904
rect 8280 5904 8298 5922
rect 8280 5922 8298 5940
rect 8280 5940 8298 5958
rect 8280 5958 8298 5976
rect 8280 5976 8298 5994
rect 8280 5994 8298 6012
rect 8280 6012 8298 6030
rect 8280 6030 8298 6048
rect 8280 6048 8298 6066
rect 8280 6066 8298 6084
rect 8280 6084 8298 6102
rect 8280 6102 8298 6120
rect 8280 6120 8298 6138
rect 8280 6138 8298 6156
rect 8280 6156 8298 6174
rect 8280 6174 8298 6192
rect 8280 6192 8298 6210
rect 8280 6210 8298 6228
rect 8280 6228 8298 6246
rect 8280 6246 8298 6264
rect 8280 6264 8298 6282
rect 8280 6282 8298 6300
rect 8280 6300 8298 6318
rect 8280 6318 8298 6336
rect 8280 6336 8298 6354
rect 8280 6354 8298 6372
rect 8280 6372 8298 6390
rect 8280 6390 8298 6408
rect 8280 6408 8298 6426
rect 8280 6426 8298 6444
rect 8280 6444 8298 6462
rect 8280 6462 8298 6480
rect 8280 6480 8298 6498
rect 8280 6498 8298 6516
rect 8280 6516 8298 6534
rect 8280 6534 8298 6552
rect 8280 6552 8298 6570
rect 8280 6570 8298 6588
rect 8280 6588 8298 6606
rect 8280 6606 8298 6624
rect 8280 6624 8298 6642
rect 8280 6642 8298 6660
rect 8280 6660 8298 6678
rect 8280 6678 8298 6696
rect 8280 6696 8298 6714
rect 8280 6714 8298 6732
rect 8280 6732 8298 6750
rect 8280 6750 8298 6768
rect 8280 6768 8298 6786
rect 8280 6786 8298 6804
rect 8280 6804 8298 6822
rect 8280 6822 8298 6840
rect 8280 6840 8298 6858
rect 8280 6858 8298 6876
rect 8280 6876 8298 6894
rect 8280 6894 8298 6912
rect 8280 6912 8298 6930
rect 8280 6930 8298 6948
rect 8280 6948 8298 6966
rect 8280 6966 8298 6984
rect 8280 6984 8298 7002
rect 8280 7002 8298 7020
rect 8280 7020 8298 7038
rect 8280 7038 8298 7056
rect 8280 7056 8298 7074
rect 8280 7074 8298 7092
rect 8280 7092 8298 7110
rect 8280 7110 8298 7128
rect 8280 7128 8298 7146
rect 8280 7146 8298 7164
rect 8280 7164 8298 7182
rect 8280 7182 8298 7200
rect 8280 7200 8298 7218
rect 8298 2628 8316 2646
rect 8298 2646 8316 2664
rect 8298 2664 8316 2682
rect 8298 2682 8316 2700
rect 8298 2700 8316 2718
rect 8298 2718 8316 2736
rect 8298 2736 8316 2754
rect 8298 2754 8316 2772
rect 8298 2772 8316 2790
rect 8298 2790 8316 2808
rect 8298 2808 8316 2826
rect 8298 2826 8316 2844
rect 8298 2844 8316 2862
rect 8298 2862 8316 2880
rect 8298 2880 8316 2898
rect 8298 2898 8316 2916
rect 8298 2916 8316 2934
rect 8298 2934 8316 2952
rect 8298 2952 8316 2970
rect 8298 2970 8316 2988
rect 8298 2988 8316 3006
rect 8298 3006 8316 3024
rect 8298 3024 8316 3042
rect 8298 3042 8316 3060
rect 8298 3060 8316 3078
rect 8298 3078 8316 3096
rect 8298 3096 8316 3114
rect 8298 3114 8316 3132
rect 8298 3132 8316 3150
rect 8298 3150 8316 3168
rect 8298 3168 8316 3186
rect 8298 3186 8316 3204
rect 8298 3204 8316 3222
rect 8298 3222 8316 3240
rect 8298 3240 8316 3258
rect 8298 3258 8316 3276
rect 8298 3276 8316 3294
rect 8298 3294 8316 3312
rect 8298 3312 8316 3330
rect 8298 3330 8316 3348
rect 8298 3348 8316 3366
rect 8298 3366 8316 3384
rect 8298 3384 8316 3402
rect 8298 3402 8316 3420
rect 8298 3420 8316 3438
rect 8298 5670 8316 5688
rect 8298 5688 8316 5706
rect 8298 5706 8316 5724
rect 8298 5724 8316 5742
rect 8298 5742 8316 5760
rect 8298 5760 8316 5778
rect 8298 5778 8316 5796
rect 8298 5796 8316 5814
rect 8298 5814 8316 5832
rect 8298 5832 8316 5850
rect 8298 5850 8316 5868
rect 8298 5868 8316 5886
rect 8298 5886 8316 5904
rect 8298 5904 8316 5922
rect 8298 5922 8316 5940
rect 8298 5940 8316 5958
rect 8298 5958 8316 5976
rect 8298 5976 8316 5994
rect 8298 5994 8316 6012
rect 8298 6012 8316 6030
rect 8298 6030 8316 6048
rect 8298 6048 8316 6066
rect 8298 6066 8316 6084
rect 8298 6084 8316 6102
rect 8298 6102 8316 6120
rect 8298 6120 8316 6138
rect 8298 6138 8316 6156
rect 8298 6156 8316 6174
rect 8298 6174 8316 6192
rect 8298 6192 8316 6210
rect 8298 6210 8316 6228
rect 8298 6228 8316 6246
rect 8298 6246 8316 6264
rect 8298 6264 8316 6282
rect 8298 6282 8316 6300
rect 8298 6300 8316 6318
rect 8298 6318 8316 6336
rect 8298 6336 8316 6354
rect 8298 6354 8316 6372
rect 8298 6372 8316 6390
rect 8298 6390 8316 6408
rect 8298 6408 8316 6426
rect 8298 6426 8316 6444
rect 8298 6444 8316 6462
rect 8298 6462 8316 6480
rect 8298 6480 8316 6498
rect 8298 6498 8316 6516
rect 8298 6516 8316 6534
rect 8298 6534 8316 6552
rect 8298 6552 8316 6570
rect 8298 6570 8316 6588
rect 8298 6588 8316 6606
rect 8298 6606 8316 6624
rect 8298 6624 8316 6642
rect 8298 6642 8316 6660
rect 8298 6660 8316 6678
rect 8298 6678 8316 6696
rect 8298 6696 8316 6714
rect 8298 6714 8316 6732
rect 8298 6732 8316 6750
rect 8298 6750 8316 6768
rect 8298 6768 8316 6786
rect 8298 6786 8316 6804
rect 8298 6804 8316 6822
rect 8298 6822 8316 6840
rect 8298 6840 8316 6858
rect 8298 6858 8316 6876
rect 8298 6876 8316 6894
rect 8298 6894 8316 6912
rect 8298 6912 8316 6930
rect 8298 6930 8316 6948
rect 8298 6948 8316 6966
rect 8298 6966 8316 6984
rect 8298 6984 8316 7002
rect 8298 7002 8316 7020
rect 8298 7020 8316 7038
rect 8298 7038 8316 7056
rect 8298 7056 8316 7074
rect 8298 7074 8316 7092
rect 8298 7092 8316 7110
rect 8298 7110 8316 7128
rect 8298 7128 8316 7146
rect 8298 7146 8316 7164
rect 8298 7164 8316 7182
rect 8298 7182 8316 7200
rect 8298 7200 8316 7218
rect 8298 7218 8316 7236
rect 8316 2646 8334 2664
rect 8316 2664 8334 2682
rect 8316 2682 8334 2700
rect 8316 2700 8334 2718
rect 8316 2718 8334 2736
rect 8316 2736 8334 2754
rect 8316 2754 8334 2772
rect 8316 2772 8334 2790
rect 8316 2790 8334 2808
rect 8316 2808 8334 2826
rect 8316 2826 8334 2844
rect 8316 2844 8334 2862
rect 8316 2862 8334 2880
rect 8316 2880 8334 2898
rect 8316 2898 8334 2916
rect 8316 2916 8334 2934
rect 8316 2934 8334 2952
rect 8316 2952 8334 2970
rect 8316 2970 8334 2988
rect 8316 2988 8334 3006
rect 8316 3006 8334 3024
rect 8316 3024 8334 3042
rect 8316 3042 8334 3060
rect 8316 3060 8334 3078
rect 8316 3078 8334 3096
rect 8316 3096 8334 3114
rect 8316 3114 8334 3132
rect 8316 3132 8334 3150
rect 8316 3150 8334 3168
rect 8316 3168 8334 3186
rect 8316 3186 8334 3204
rect 8316 3204 8334 3222
rect 8316 3222 8334 3240
rect 8316 3240 8334 3258
rect 8316 3258 8334 3276
rect 8316 3276 8334 3294
rect 8316 3294 8334 3312
rect 8316 3312 8334 3330
rect 8316 3330 8334 3348
rect 8316 3348 8334 3366
rect 8316 3366 8334 3384
rect 8316 3384 8334 3402
rect 8316 3402 8334 3420
rect 8316 3420 8334 3438
rect 8316 5688 8334 5706
rect 8316 5706 8334 5724
rect 8316 5724 8334 5742
rect 8316 5742 8334 5760
rect 8316 5760 8334 5778
rect 8316 5778 8334 5796
rect 8316 5796 8334 5814
rect 8316 5814 8334 5832
rect 8316 5832 8334 5850
rect 8316 5850 8334 5868
rect 8316 5868 8334 5886
rect 8316 5886 8334 5904
rect 8316 5904 8334 5922
rect 8316 5922 8334 5940
rect 8316 5940 8334 5958
rect 8316 5958 8334 5976
rect 8316 5976 8334 5994
rect 8316 5994 8334 6012
rect 8316 6012 8334 6030
rect 8316 6030 8334 6048
rect 8316 6048 8334 6066
rect 8316 6066 8334 6084
rect 8316 6084 8334 6102
rect 8316 6102 8334 6120
rect 8316 6120 8334 6138
rect 8316 6138 8334 6156
rect 8316 6156 8334 6174
rect 8316 6174 8334 6192
rect 8316 6192 8334 6210
rect 8316 6210 8334 6228
rect 8316 6228 8334 6246
rect 8316 6246 8334 6264
rect 8316 6264 8334 6282
rect 8316 6282 8334 6300
rect 8316 6300 8334 6318
rect 8316 6318 8334 6336
rect 8316 6336 8334 6354
rect 8316 6354 8334 6372
rect 8316 6372 8334 6390
rect 8316 6390 8334 6408
rect 8316 6408 8334 6426
rect 8316 6426 8334 6444
rect 8316 6444 8334 6462
rect 8316 6462 8334 6480
rect 8316 6480 8334 6498
rect 8316 6498 8334 6516
rect 8316 6516 8334 6534
rect 8316 6534 8334 6552
rect 8316 6552 8334 6570
rect 8316 6570 8334 6588
rect 8316 6588 8334 6606
rect 8316 6606 8334 6624
rect 8316 6624 8334 6642
rect 8316 6642 8334 6660
rect 8316 6660 8334 6678
rect 8316 6678 8334 6696
rect 8316 6696 8334 6714
rect 8316 6714 8334 6732
rect 8316 6732 8334 6750
rect 8316 6750 8334 6768
rect 8316 6768 8334 6786
rect 8316 6786 8334 6804
rect 8316 6804 8334 6822
rect 8316 6822 8334 6840
rect 8316 6840 8334 6858
rect 8316 6858 8334 6876
rect 8316 6876 8334 6894
rect 8316 6894 8334 6912
rect 8316 6912 8334 6930
rect 8316 6930 8334 6948
rect 8316 6948 8334 6966
rect 8316 6966 8334 6984
rect 8316 6984 8334 7002
rect 8316 7002 8334 7020
rect 8316 7020 8334 7038
rect 8316 7038 8334 7056
rect 8316 7056 8334 7074
rect 8316 7074 8334 7092
rect 8316 7092 8334 7110
rect 8316 7110 8334 7128
rect 8316 7128 8334 7146
rect 8316 7146 8334 7164
rect 8316 7164 8334 7182
rect 8316 7182 8334 7200
rect 8316 7200 8334 7218
rect 8316 7218 8334 7236
rect 8334 2646 8352 2664
rect 8334 2664 8352 2682
rect 8334 2682 8352 2700
rect 8334 2700 8352 2718
rect 8334 2718 8352 2736
rect 8334 2736 8352 2754
rect 8334 2754 8352 2772
rect 8334 2772 8352 2790
rect 8334 2790 8352 2808
rect 8334 2808 8352 2826
rect 8334 2826 8352 2844
rect 8334 2844 8352 2862
rect 8334 2862 8352 2880
rect 8334 2880 8352 2898
rect 8334 2898 8352 2916
rect 8334 2916 8352 2934
rect 8334 2934 8352 2952
rect 8334 2952 8352 2970
rect 8334 2970 8352 2988
rect 8334 2988 8352 3006
rect 8334 3006 8352 3024
rect 8334 3024 8352 3042
rect 8334 3042 8352 3060
rect 8334 3060 8352 3078
rect 8334 3078 8352 3096
rect 8334 3096 8352 3114
rect 8334 3114 8352 3132
rect 8334 3132 8352 3150
rect 8334 3150 8352 3168
rect 8334 3168 8352 3186
rect 8334 3186 8352 3204
rect 8334 3204 8352 3222
rect 8334 3222 8352 3240
rect 8334 3240 8352 3258
rect 8334 3258 8352 3276
rect 8334 3276 8352 3294
rect 8334 3294 8352 3312
rect 8334 3312 8352 3330
rect 8334 3330 8352 3348
rect 8334 3348 8352 3366
rect 8334 3366 8352 3384
rect 8334 3384 8352 3402
rect 8334 3402 8352 3420
rect 8334 3420 8352 3438
rect 8334 3438 8352 3456
rect 8334 5724 8352 5742
rect 8334 5742 8352 5760
rect 8334 5760 8352 5778
rect 8334 5778 8352 5796
rect 8334 5796 8352 5814
rect 8334 5814 8352 5832
rect 8334 5832 8352 5850
rect 8334 5850 8352 5868
rect 8334 5868 8352 5886
rect 8334 5886 8352 5904
rect 8334 5904 8352 5922
rect 8334 5922 8352 5940
rect 8334 5940 8352 5958
rect 8334 5958 8352 5976
rect 8334 5976 8352 5994
rect 8334 5994 8352 6012
rect 8334 6012 8352 6030
rect 8334 6030 8352 6048
rect 8334 6048 8352 6066
rect 8334 6066 8352 6084
rect 8334 6084 8352 6102
rect 8334 6102 8352 6120
rect 8334 6120 8352 6138
rect 8334 6138 8352 6156
rect 8334 6156 8352 6174
rect 8334 6174 8352 6192
rect 8334 6192 8352 6210
rect 8334 6210 8352 6228
rect 8334 6228 8352 6246
rect 8334 6246 8352 6264
rect 8334 6264 8352 6282
rect 8334 6282 8352 6300
rect 8334 6300 8352 6318
rect 8334 6318 8352 6336
rect 8334 6336 8352 6354
rect 8334 6354 8352 6372
rect 8334 6372 8352 6390
rect 8334 6390 8352 6408
rect 8334 6408 8352 6426
rect 8334 6426 8352 6444
rect 8334 6444 8352 6462
rect 8334 6462 8352 6480
rect 8334 6480 8352 6498
rect 8334 6498 8352 6516
rect 8334 6516 8352 6534
rect 8334 6534 8352 6552
rect 8334 6552 8352 6570
rect 8334 6570 8352 6588
rect 8334 6588 8352 6606
rect 8334 6606 8352 6624
rect 8334 6624 8352 6642
rect 8334 6642 8352 6660
rect 8334 6660 8352 6678
rect 8334 6678 8352 6696
rect 8334 6696 8352 6714
rect 8334 6714 8352 6732
rect 8334 6732 8352 6750
rect 8334 6750 8352 6768
rect 8334 6768 8352 6786
rect 8334 6786 8352 6804
rect 8334 6804 8352 6822
rect 8334 6822 8352 6840
rect 8334 6840 8352 6858
rect 8334 6858 8352 6876
rect 8334 6876 8352 6894
rect 8334 6894 8352 6912
rect 8334 6912 8352 6930
rect 8334 6930 8352 6948
rect 8334 6948 8352 6966
rect 8334 6966 8352 6984
rect 8334 6984 8352 7002
rect 8334 7002 8352 7020
rect 8334 7020 8352 7038
rect 8334 7038 8352 7056
rect 8334 7056 8352 7074
rect 8334 7074 8352 7092
rect 8334 7092 8352 7110
rect 8334 7110 8352 7128
rect 8334 7128 8352 7146
rect 8334 7146 8352 7164
rect 8334 7164 8352 7182
rect 8334 7182 8352 7200
rect 8334 7200 8352 7218
rect 8334 7218 8352 7236
rect 8334 7236 8352 7254
rect 8352 2664 8370 2682
rect 8352 2682 8370 2700
rect 8352 2700 8370 2718
rect 8352 2718 8370 2736
rect 8352 2736 8370 2754
rect 8352 2754 8370 2772
rect 8352 2772 8370 2790
rect 8352 2790 8370 2808
rect 8352 2808 8370 2826
rect 8352 2826 8370 2844
rect 8352 2844 8370 2862
rect 8352 2862 8370 2880
rect 8352 2880 8370 2898
rect 8352 2898 8370 2916
rect 8352 2916 8370 2934
rect 8352 2934 8370 2952
rect 8352 2952 8370 2970
rect 8352 2970 8370 2988
rect 8352 2988 8370 3006
rect 8352 3006 8370 3024
rect 8352 3024 8370 3042
rect 8352 3042 8370 3060
rect 8352 3060 8370 3078
rect 8352 3078 8370 3096
rect 8352 3096 8370 3114
rect 8352 3114 8370 3132
rect 8352 3132 8370 3150
rect 8352 3150 8370 3168
rect 8352 3168 8370 3186
rect 8352 3186 8370 3204
rect 8352 3204 8370 3222
rect 8352 3222 8370 3240
rect 8352 3240 8370 3258
rect 8352 3258 8370 3276
rect 8352 3276 8370 3294
rect 8352 3294 8370 3312
rect 8352 3312 8370 3330
rect 8352 3330 8370 3348
rect 8352 3348 8370 3366
rect 8352 3366 8370 3384
rect 8352 3384 8370 3402
rect 8352 3402 8370 3420
rect 8352 3420 8370 3438
rect 8352 3438 8370 3456
rect 8352 5742 8370 5760
rect 8352 5760 8370 5778
rect 8352 5778 8370 5796
rect 8352 5796 8370 5814
rect 8352 5814 8370 5832
rect 8352 5832 8370 5850
rect 8352 5850 8370 5868
rect 8352 5868 8370 5886
rect 8352 5886 8370 5904
rect 8352 5904 8370 5922
rect 8352 5922 8370 5940
rect 8352 5940 8370 5958
rect 8352 5958 8370 5976
rect 8352 5976 8370 5994
rect 8352 5994 8370 6012
rect 8352 6012 8370 6030
rect 8352 6030 8370 6048
rect 8352 6048 8370 6066
rect 8352 6066 8370 6084
rect 8352 6084 8370 6102
rect 8352 6102 8370 6120
rect 8352 6120 8370 6138
rect 8352 6138 8370 6156
rect 8352 6156 8370 6174
rect 8352 6174 8370 6192
rect 8352 6192 8370 6210
rect 8352 6210 8370 6228
rect 8352 6228 8370 6246
rect 8352 6246 8370 6264
rect 8352 6264 8370 6282
rect 8352 6282 8370 6300
rect 8352 6300 8370 6318
rect 8352 6318 8370 6336
rect 8352 6336 8370 6354
rect 8352 6354 8370 6372
rect 8352 6372 8370 6390
rect 8352 6390 8370 6408
rect 8352 6408 8370 6426
rect 8352 6426 8370 6444
rect 8352 6444 8370 6462
rect 8352 6462 8370 6480
rect 8352 6480 8370 6498
rect 8352 6498 8370 6516
rect 8352 6516 8370 6534
rect 8352 6534 8370 6552
rect 8352 6552 8370 6570
rect 8352 6570 8370 6588
rect 8352 6588 8370 6606
rect 8352 6606 8370 6624
rect 8352 6624 8370 6642
rect 8352 6642 8370 6660
rect 8352 6660 8370 6678
rect 8352 6678 8370 6696
rect 8352 6696 8370 6714
rect 8352 6714 8370 6732
rect 8352 6732 8370 6750
rect 8352 6750 8370 6768
rect 8352 6768 8370 6786
rect 8352 6786 8370 6804
rect 8352 6804 8370 6822
rect 8352 6822 8370 6840
rect 8352 6840 8370 6858
rect 8352 6858 8370 6876
rect 8352 6876 8370 6894
rect 8352 6894 8370 6912
rect 8352 6912 8370 6930
rect 8352 6930 8370 6948
rect 8352 6948 8370 6966
rect 8352 6966 8370 6984
rect 8352 6984 8370 7002
rect 8352 7002 8370 7020
rect 8352 7020 8370 7038
rect 8352 7038 8370 7056
rect 8352 7056 8370 7074
rect 8352 7074 8370 7092
rect 8352 7092 8370 7110
rect 8352 7110 8370 7128
rect 8352 7128 8370 7146
rect 8352 7146 8370 7164
rect 8352 7164 8370 7182
rect 8352 7182 8370 7200
rect 8352 7200 8370 7218
rect 8352 7218 8370 7236
rect 8352 7236 8370 7254
rect 8352 7254 8370 7272
rect 8370 2682 8388 2700
rect 8370 2700 8388 2718
rect 8370 2718 8388 2736
rect 8370 2736 8388 2754
rect 8370 2754 8388 2772
rect 8370 2772 8388 2790
rect 8370 2790 8388 2808
rect 8370 2808 8388 2826
rect 8370 2826 8388 2844
rect 8370 2844 8388 2862
rect 8370 2862 8388 2880
rect 8370 2880 8388 2898
rect 8370 2898 8388 2916
rect 8370 2916 8388 2934
rect 8370 2934 8388 2952
rect 8370 2952 8388 2970
rect 8370 2970 8388 2988
rect 8370 2988 8388 3006
rect 8370 3006 8388 3024
rect 8370 3024 8388 3042
rect 8370 3042 8388 3060
rect 8370 3060 8388 3078
rect 8370 3078 8388 3096
rect 8370 3096 8388 3114
rect 8370 3114 8388 3132
rect 8370 3132 8388 3150
rect 8370 3150 8388 3168
rect 8370 3168 8388 3186
rect 8370 3186 8388 3204
rect 8370 3204 8388 3222
rect 8370 3222 8388 3240
rect 8370 3240 8388 3258
rect 8370 3258 8388 3276
rect 8370 3276 8388 3294
rect 8370 3294 8388 3312
rect 8370 3312 8388 3330
rect 8370 3330 8388 3348
rect 8370 3348 8388 3366
rect 8370 3366 8388 3384
rect 8370 3384 8388 3402
rect 8370 3402 8388 3420
rect 8370 3420 8388 3438
rect 8370 3438 8388 3456
rect 8370 5778 8388 5796
rect 8370 5796 8388 5814
rect 8370 5814 8388 5832
rect 8370 5832 8388 5850
rect 8370 5850 8388 5868
rect 8370 5868 8388 5886
rect 8370 5886 8388 5904
rect 8370 5904 8388 5922
rect 8370 5922 8388 5940
rect 8370 5940 8388 5958
rect 8370 5958 8388 5976
rect 8370 5976 8388 5994
rect 8370 5994 8388 6012
rect 8370 6012 8388 6030
rect 8370 6030 8388 6048
rect 8370 6048 8388 6066
rect 8370 6066 8388 6084
rect 8370 6084 8388 6102
rect 8370 6102 8388 6120
rect 8370 6120 8388 6138
rect 8370 6138 8388 6156
rect 8370 6156 8388 6174
rect 8370 6174 8388 6192
rect 8370 6192 8388 6210
rect 8370 6210 8388 6228
rect 8370 6228 8388 6246
rect 8370 6246 8388 6264
rect 8370 6264 8388 6282
rect 8370 6282 8388 6300
rect 8370 6300 8388 6318
rect 8370 6318 8388 6336
rect 8370 6336 8388 6354
rect 8370 6354 8388 6372
rect 8370 6372 8388 6390
rect 8370 6390 8388 6408
rect 8370 6408 8388 6426
rect 8370 6426 8388 6444
rect 8370 6444 8388 6462
rect 8370 6462 8388 6480
rect 8370 6480 8388 6498
rect 8370 6498 8388 6516
rect 8370 6516 8388 6534
rect 8370 6534 8388 6552
rect 8370 6552 8388 6570
rect 8370 6570 8388 6588
rect 8370 6588 8388 6606
rect 8370 6606 8388 6624
rect 8370 6624 8388 6642
rect 8370 6642 8388 6660
rect 8370 6660 8388 6678
rect 8370 6678 8388 6696
rect 8370 6696 8388 6714
rect 8370 6714 8388 6732
rect 8370 6732 8388 6750
rect 8370 6750 8388 6768
rect 8370 6768 8388 6786
rect 8370 6786 8388 6804
rect 8370 6804 8388 6822
rect 8370 6822 8388 6840
rect 8370 6840 8388 6858
rect 8370 6858 8388 6876
rect 8370 6876 8388 6894
rect 8370 6894 8388 6912
rect 8370 6912 8388 6930
rect 8370 6930 8388 6948
rect 8370 6948 8388 6966
rect 8370 6966 8388 6984
rect 8370 6984 8388 7002
rect 8370 7002 8388 7020
rect 8370 7020 8388 7038
rect 8370 7038 8388 7056
rect 8370 7056 8388 7074
rect 8370 7074 8388 7092
rect 8370 7092 8388 7110
rect 8370 7110 8388 7128
rect 8370 7128 8388 7146
rect 8370 7146 8388 7164
rect 8370 7164 8388 7182
rect 8370 7182 8388 7200
rect 8370 7200 8388 7218
rect 8370 7218 8388 7236
rect 8370 7236 8388 7254
rect 8370 7254 8388 7272
rect 8388 2700 8406 2718
rect 8388 2718 8406 2736
rect 8388 2736 8406 2754
rect 8388 2754 8406 2772
rect 8388 2772 8406 2790
rect 8388 2790 8406 2808
rect 8388 2808 8406 2826
rect 8388 2826 8406 2844
rect 8388 2844 8406 2862
rect 8388 2862 8406 2880
rect 8388 2880 8406 2898
rect 8388 2898 8406 2916
rect 8388 2916 8406 2934
rect 8388 2934 8406 2952
rect 8388 2952 8406 2970
rect 8388 2970 8406 2988
rect 8388 2988 8406 3006
rect 8388 3006 8406 3024
rect 8388 3024 8406 3042
rect 8388 3042 8406 3060
rect 8388 3060 8406 3078
rect 8388 3078 8406 3096
rect 8388 3096 8406 3114
rect 8388 3114 8406 3132
rect 8388 3132 8406 3150
rect 8388 3150 8406 3168
rect 8388 3168 8406 3186
rect 8388 3186 8406 3204
rect 8388 3204 8406 3222
rect 8388 3222 8406 3240
rect 8388 3240 8406 3258
rect 8388 3258 8406 3276
rect 8388 3276 8406 3294
rect 8388 3294 8406 3312
rect 8388 3312 8406 3330
rect 8388 3330 8406 3348
rect 8388 3348 8406 3366
rect 8388 3366 8406 3384
rect 8388 3384 8406 3402
rect 8388 3402 8406 3420
rect 8388 3420 8406 3438
rect 8388 3438 8406 3456
rect 8388 5796 8406 5814
rect 8388 5814 8406 5832
rect 8388 5832 8406 5850
rect 8388 5850 8406 5868
rect 8388 5868 8406 5886
rect 8388 5886 8406 5904
rect 8388 5904 8406 5922
rect 8388 5922 8406 5940
rect 8388 5940 8406 5958
rect 8388 5958 8406 5976
rect 8388 5976 8406 5994
rect 8388 5994 8406 6012
rect 8388 6012 8406 6030
rect 8388 6030 8406 6048
rect 8388 6048 8406 6066
rect 8388 6066 8406 6084
rect 8388 6084 8406 6102
rect 8388 6102 8406 6120
rect 8388 6120 8406 6138
rect 8388 6138 8406 6156
rect 8388 6156 8406 6174
rect 8388 6174 8406 6192
rect 8388 6192 8406 6210
rect 8388 6210 8406 6228
rect 8388 6228 8406 6246
rect 8388 6246 8406 6264
rect 8388 6264 8406 6282
rect 8388 6282 8406 6300
rect 8388 6300 8406 6318
rect 8388 6318 8406 6336
rect 8388 6336 8406 6354
rect 8388 6354 8406 6372
rect 8388 6372 8406 6390
rect 8388 6390 8406 6408
rect 8388 6408 8406 6426
rect 8388 6426 8406 6444
rect 8388 6444 8406 6462
rect 8388 6462 8406 6480
rect 8388 6480 8406 6498
rect 8388 6498 8406 6516
rect 8388 6516 8406 6534
rect 8388 6534 8406 6552
rect 8388 6552 8406 6570
rect 8388 6570 8406 6588
rect 8388 6588 8406 6606
rect 8388 6606 8406 6624
rect 8388 6624 8406 6642
rect 8388 6642 8406 6660
rect 8388 6660 8406 6678
rect 8388 6678 8406 6696
rect 8388 6696 8406 6714
rect 8388 6714 8406 6732
rect 8388 6732 8406 6750
rect 8388 6750 8406 6768
rect 8388 6768 8406 6786
rect 8388 6786 8406 6804
rect 8388 6804 8406 6822
rect 8388 6822 8406 6840
rect 8388 6840 8406 6858
rect 8388 6858 8406 6876
rect 8388 6876 8406 6894
rect 8388 6894 8406 6912
rect 8388 6912 8406 6930
rect 8388 6930 8406 6948
rect 8388 6948 8406 6966
rect 8388 6966 8406 6984
rect 8388 6984 8406 7002
rect 8388 7002 8406 7020
rect 8388 7020 8406 7038
rect 8388 7038 8406 7056
rect 8388 7056 8406 7074
rect 8388 7074 8406 7092
rect 8388 7092 8406 7110
rect 8388 7110 8406 7128
rect 8388 7128 8406 7146
rect 8388 7146 8406 7164
rect 8388 7164 8406 7182
rect 8388 7182 8406 7200
rect 8388 7200 8406 7218
rect 8388 7218 8406 7236
rect 8388 7236 8406 7254
rect 8388 7254 8406 7272
rect 8388 7272 8406 7290
rect 8406 2718 8424 2736
rect 8406 2736 8424 2754
rect 8406 2754 8424 2772
rect 8406 2772 8424 2790
rect 8406 2790 8424 2808
rect 8406 2808 8424 2826
rect 8406 2826 8424 2844
rect 8406 2844 8424 2862
rect 8406 2862 8424 2880
rect 8406 2880 8424 2898
rect 8406 2898 8424 2916
rect 8406 2916 8424 2934
rect 8406 2934 8424 2952
rect 8406 2952 8424 2970
rect 8406 2970 8424 2988
rect 8406 2988 8424 3006
rect 8406 3006 8424 3024
rect 8406 3024 8424 3042
rect 8406 3042 8424 3060
rect 8406 3060 8424 3078
rect 8406 3078 8424 3096
rect 8406 3096 8424 3114
rect 8406 3114 8424 3132
rect 8406 3132 8424 3150
rect 8406 3150 8424 3168
rect 8406 3168 8424 3186
rect 8406 3186 8424 3204
rect 8406 3204 8424 3222
rect 8406 3222 8424 3240
rect 8406 3240 8424 3258
rect 8406 3258 8424 3276
rect 8406 3276 8424 3294
rect 8406 3294 8424 3312
rect 8406 3312 8424 3330
rect 8406 3330 8424 3348
rect 8406 3348 8424 3366
rect 8406 3366 8424 3384
rect 8406 3384 8424 3402
rect 8406 3402 8424 3420
rect 8406 3420 8424 3438
rect 8406 3438 8424 3456
rect 8406 3456 8424 3474
rect 8406 5832 8424 5850
rect 8406 5850 8424 5868
rect 8406 5868 8424 5886
rect 8406 5886 8424 5904
rect 8406 5904 8424 5922
rect 8406 5922 8424 5940
rect 8406 5940 8424 5958
rect 8406 5958 8424 5976
rect 8406 5976 8424 5994
rect 8406 5994 8424 6012
rect 8406 6012 8424 6030
rect 8406 6030 8424 6048
rect 8406 6048 8424 6066
rect 8406 6066 8424 6084
rect 8406 6084 8424 6102
rect 8406 6102 8424 6120
rect 8406 6120 8424 6138
rect 8406 6138 8424 6156
rect 8406 6156 8424 6174
rect 8406 6174 8424 6192
rect 8406 6192 8424 6210
rect 8406 6210 8424 6228
rect 8406 6228 8424 6246
rect 8406 6246 8424 6264
rect 8406 6264 8424 6282
rect 8406 6282 8424 6300
rect 8406 6300 8424 6318
rect 8406 6318 8424 6336
rect 8406 6336 8424 6354
rect 8406 6354 8424 6372
rect 8406 6372 8424 6390
rect 8406 6390 8424 6408
rect 8406 6408 8424 6426
rect 8406 6426 8424 6444
rect 8406 6444 8424 6462
rect 8406 6462 8424 6480
rect 8406 6480 8424 6498
rect 8406 6498 8424 6516
rect 8406 6516 8424 6534
rect 8406 6534 8424 6552
rect 8406 6552 8424 6570
rect 8406 6570 8424 6588
rect 8406 6588 8424 6606
rect 8406 6606 8424 6624
rect 8406 6624 8424 6642
rect 8406 6642 8424 6660
rect 8406 6660 8424 6678
rect 8406 6678 8424 6696
rect 8406 6696 8424 6714
rect 8406 6714 8424 6732
rect 8406 6732 8424 6750
rect 8406 6750 8424 6768
rect 8406 6768 8424 6786
rect 8406 6786 8424 6804
rect 8406 6804 8424 6822
rect 8406 6822 8424 6840
rect 8406 6840 8424 6858
rect 8406 6858 8424 6876
rect 8406 6876 8424 6894
rect 8406 6894 8424 6912
rect 8406 6912 8424 6930
rect 8406 6930 8424 6948
rect 8406 6948 8424 6966
rect 8406 6966 8424 6984
rect 8406 6984 8424 7002
rect 8406 7002 8424 7020
rect 8406 7020 8424 7038
rect 8406 7038 8424 7056
rect 8406 7056 8424 7074
rect 8406 7074 8424 7092
rect 8406 7092 8424 7110
rect 8406 7110 8424 7128
rect 8406 7128 8424 7146
rect 8406 7146 8424 7164
rect 8406 7164 8424 7182
rect 8406 7182 8424 7200
rect 8406 7200 8424 7218
rect 8406 7218 8424 7236
rect 8406 7236 8424 7254
rect 8406 7254 8424 7272
rect 8406 7272 8424 7290
rect 8406 7290 8424 7308
rect 8424 2736 8442 2754
rect 8424 2754 8442 2772
rect 8424 2772 8442 2790
rect 8424 2790 8442 2808
rect 8424 2808 8442 2826
rect 8424 2826 8442 2844
rect 8424 2844 8442 2862
rect 8424 2862 8442 2880
rect 8424 2880 8442 2898
rect 8424 2898 8442 2916
rect 8424 2916 8442 2934
rect 8424 2934 8442 2952
rect 8424 2952 8442 2970
rect 8424 2970 8442 2988
rect 8424 2988 8442 3006
rect 8424 3006 8442 3024
rect 8424 3024 8442 3042
rect 8424 3042 8442 3060
rect 8424 3060 8442 3078
rect 8424 3078 8442 3096
rect 8424 3096 8442 3114
rect 8424 3114 8442 3132
rect 8424 3132 8442 3150
rect 8424 3150 8442 3168
rect 8424 3168 8442 3186
rect 8424 3186 8442 3204
rect 8424 3204 8442 3222
rect 8424 3222 8442 3240
rect 8424 3240 8442 3258
rect 8424 3258 8442 3276
rect 8424 3276 8442 3294
rect 8424 3294 8442 3312
rect 8424 3312 8442 3330
rect 8424 3330 8442 3348
rect 8424 3348 8442 3366
rect 8424 3366 8442 3384
rect 8424 3384 8442 3402
rect 8424 3402 8442 3420
rect 8424 3420 8442 3438
rect 8424 3438 8442 3456
rect 8424 3456 8442 3474
rect 8424 5868 8442 5886
rect 8424 5886 8442 5904
rect 8424 5904 8442 5922
rect 8424 5922 8442 5940
rect 8424 5940 8442 5958
rect 8424 5958 8442 5976
rect 8424 5976 8442 5994
rect 8424 5994 8442 6012
rect 8424 6012 8442 6030
rect 8424 6030 8442 6048
rect 8424 6048 8442 6066
rect 8424 6066 8442 6084
rect 8424 6084 8442 6102
rect 8424 6102 8442 6120
rect 8424 6120 8442 6138
rect 8424 6138 8442 6156
rect 8424 6156 8442 6174
rect 8424 6174 8442 6192
rect 8424 6192 8442 6210
rect 8424 6210 8442 6228
rect 8424 6228 8442 6246
rect 8424 6246 8442 6264
rect 8424 6264 8442 6282
rect 8424 6282 8442 6300
rect 8424 6300 8442 6318
rect 8424 6318 8442 6336
rect 8424 6336 8442 6354
rect 8424 6354 8442 6372
rect 8424 6372 8442 6390
rect 8424 6390 8442 6408
rect 8424 6408 8442 6426
rect 8424 6426 8442 6444
rect 8424 6444 8442 6462
rect 8424 6462 8442 6480
rect 8424 6480 8442 6498
rect 8424 6498 8442 6516
rect 8424 6516 8442 6534
rect 8424 6534 8442 6552
rect 8424 6552 8442 6570
rect 8424 6570 8442 6588
rect 8424 6588 8442 6606
rect 8424 6606 8442 6624
rect 8424 6624 8442 6642
rect 8424 6642 8442 6660
rect 8424 6660 8442 6678
rect 8424 6678 8442 6696
rect 8424 6696 8442 6714
rect 8424 6714 8442 6732
rect 8424 6732 8442 6750
rect 8424 6750 8442 6768
rect 8424 6768 8442 6786
rect 8424 6786 8442 6804
rect 8424 6804 8442 6822
rect 8424 6822 8442 6840
rect 8424 6840 8442 6858
rect 8424 6858 8442 6876
rect 8424 6876 8442 6894
rect 8424 6894 8442 6912
rect 8424 6912 8442 6930
rect 8424 6930 8442 6948
rect 8424 6948 8442 6966
rect 8424 6966 8442 6984
rect 8424 6984 8442 7002
rect 8424 7002 8442 7020
rect 8424 7020 8442 7038
rect 8424 7038 8442 7056
rect 8424 7056 8442 7074
rect 8424 7074 8442 7092
rect 8424 7092 8442 7110
rect 8424 7110 8442 7128
rect 8424 7128 8442 7146
rect 8424 7146 8442 7164
rect 8424 7164 8442 7182
rect 8424 7182 8442 7200
rect 8424 7200 8442 7218
rect 8424 7218 8442 7236
rect 8424 7236 8442 7254
rect 8424 7254 8442 7272
rect 8424 7272 8442 7290
rect 8424 7290 8442 7308
rect 8442 2736 8460 2754
rect 8442 2754 8460 2772
rect 8442 2772 8460 2790
rect 8442 2790 8460 2808
rect 8442 2808 8460 2826
rect 8442 2826 8460 2844
rect 8442 2844 8460 2862
rect 8442 2862 8460 2880
rect 8442 2880 8460 2898
rect 8442 2898 8460 2916
rect 8442 2916 8460 2934
rect 8442 2934 8460 2952
rect 8442 2952 8460 2970
rect 8442 2970 8460 2988
rect 8442 2988 8460 3006
rect 8442 3006 8460 3024
rect 8442 3024 8460 3042
rect 8442 3042 8460 3060
rect 8442 3060 8460 3078
rect 8442 3078 8460 3096
rect 8442 3096 8460 3114
rect 8442 3114 8460 3132
rect 8442 3132 8460 3150
rect 8442 3150 8460 3168
rect 8442 3168 8460 3186
rect 8442 3186 8460 3204
rect 8442 3204 8460 3222
rect 8442 3222 8460 3240
rect 8442 3240 8460 3258
rect 8442 3258 8460 3276
rect 8442 3276 8460 3294
rect 8442 3294 8460 3312
rect 8442 3312 8460 3330
rect 8442 3330 8460 3348
rect 8442 3348 8460 3366
rect 8442 3366 8460 3384
rect 8442 3384 8460 3402
rect 8442 3402 8460 3420
rect 8442 3420 8460 3438
rect 8442 3438 8460 3456
rect 8442 3456 8460 3474
rect 8442 5886 8460 5904
rect 8442 5904 8460 5922
rect 8442 5922 8460 5940
rect 8442 5940 8460 5958
rect 8442 5958 8460 5976
rect 8442 5976 8460 5994
rect 8442 5994 8460 6012
rect 8442 6012 8460 6030
rect 8442 6030 8460 6048
rect 8442 6048 8460 6066
rect 8442 6066 8460 6084
rect 8442 6084 8460 6102
rect 8442 6102 8460 6120
rect 8442 6120 8460 6138
rect 8442 6138 8460 6156
rect 8442 6156 8460 6174
rect 8442 6174 8460 6192
rect 8442 6192 8460 6210
rect 8442 6210 8460 6228
rect 8442 6228 8460 6246
rect 8442 6246 8460 6264
rect 8442 6264 8460 6282
rect 8442 6282 8460 6300
rect 8442 6300 8460 6318
rect 8442 6318 8460 6336
rect 8442 6336 8460 6354
rect 8442 6354 8460 6372
rect 8442 6372 8460 6390
rect 8442 6390 8460 6408
rect 8442 6408 8460 6426
rect 8442 6426 8460 6444
rect 8442 6444 8460 6462
rect 8442 6462 8460 6480
rect 8442 6480 8460 6498
rect 8442 6498 8460 6516
rect 8442 6516 8460 6534
rect 8442 6534 8460 6552
rect 8442 6552 8460 6570
rect 8442 6570 8460 6588
rect 8442 6588 8460 6606
rect 8442 6606 8460 6624
rect 8442 6624 8460 6642
rect 8442 6642 8460 6660
rect 8442 6660 8460 6678
rect 8442 6678 8460 6696
rect 8442 6696 8460 6714
rect 8442 6714 8460 6732
rect 8442 6732 8460 6750
rect 8442 6750 8460 6768
rect 8442 6768 8460 6786
rect 8442 6786 8460 6804
rect 8442 6804 8460 6822
rect 8442 6822 8460 6840
rect 8442 6840 8460 6858
rect 8442 6858 8460 6876
rect 8442 6876 8460 6894
rect 8442 6894 8460 6912
rect 8442 6912 8460 6930
rect 8442 6930 8460 6948
rect 8442 6948 8460 6966
rect 8442 6966 8460 6984
rect 8442 6984 8460 7002
rect 8442 7002 8460 7020
rect 8442 7020 8460 7038
rect 8442 7038 8460 7056
rect 8442 7056 8460 7074
rect 8442 7074 8460 7092
rect 8442 7092 8460 7110
rect 8442 7110 8460 7128
rect 8442 7128 8460 7146
rect 8442 7146 8460 7164
rect 8442 7164 8460 7182
rect 8442 7182 8460 7200
rect 8442 7200 8460 7218
rect 8442 7218 8460 7236
rect 8442 7236 8460 7254
rect 8442 7254 8460 7272
rect 8442 7272 8460 7290
rect 8442 7290 8460 7308
rect 8442 7308 8460 7326
rect 8460 2754 8478 2772
rect 8460 2772 8478 2790
rect 8460 2790 8478 2808
rect 8460 2808 8478 2826
rect 8460 2826 8478 2844
rect 8460 2844 8478 2862
rect 8460 2862 8478 2880
rect 8460 2880 8478 2898
rect 8460 2898 8478 2916
rect 8460 2916 8478 2934
rect 8460 2934 8478 2952
rect 8460 2952 8478 2970
rect 8460 2970 8478 2988
rect 8460 2988 8478 3006
rect 8460 3006 8478 3024
rect 8460 3024 8478 3042
rect 8460 3042 8478 3060
rect 8460 3060 8478 3078
rect 8460 3078 8478 3096
rect 8460 3096 8478 3114
rect 8460 3114 8478 3132
rect 8460 3132 8478 3150
rect 8460 3150 8478 3168
rect 8460 3168 8478 3186
rect 8460 3186 8478 3204
rect 8460 3204 8478 3222
rect 8460 3222 8478 3240
rect 8460 3240 8478 3258
rect 8460 3258 8478 3276
rect 8460 3276 8478 3294
rect 8460 3294 8478 3312
rect 8460 3312 8478 3330
rect 8460 3330 8478 3348
rect 8460 3348 8478 3366
rect 8460 3366 8478 3384
rect 8460 3384 8478 3402
rect 8460 3402 8478 3420
rect 8460 3420 8478 3438
rect 8460 3438 8478 3456
rect 8460 3456 8478 3474
rect 8460 5922 8478 5940
rect 8460 5940 8478 5958
rect 8460 5958 8478 5976
rect 8460 5976 8478 5994
rect 8460 5994 8478 6012
rect 8460 6012 8478 6030
rect 8460 6030 8478 6048
rect 8460 6048 8478 6066
rect 8460 6066 8478 6084
rect 8460 6084 8478 6102
rect 8460 6102 8478 6120
rect 8460 6120 8478 6138
rect 8460 6138 8478 6156
rect 8460 6156 8478 6174
rect 8460 6174 8478 6192
rect 8460 6192 8478 6210
rect 8460 6210 8478 6228
rect 8460 6228 8478 6246
rect 8460 6246 8478 6264
rect 8460 6264 8478 6282
rect 8460 6282 8478 6300
rect 8460 6300 8478 6318
rect 8460 6318 8478 6336
rect 8460 6336 8478 6354
rect 8460 6354 8478 6372
rect 8460 6372 8478 6390
rect 8460 6390 8478 6408
rect 8460 6408 8478 6426
rect 8460 6426 8478 6444
rect 8460 6444 8478 6462
rect 8460 6462 8478 6480
rect 8460 6480 8478 6498
rect 8460 6498 8478 6516
rect 8460 6516 8478 6534
rect 8460 6534 8478 6552
rect 8460 6552 8478 6570
rect 8460 6570 8478 6588
rect 8460 6588 8478 6606
rect 8460 6606 8478 6624
rect 8460 6624 8478 6642
rect 8460 6642 8478 6660
rect 8460 6660 8478 6678
rect 8460 6678 8478 6696
rect 8460 6696 8478 6714
rect 8460 6714 8478 6732
rect 8460 6732 8478 6750
rect 8460 6750 8478 6768
rect 8460 6768 8478 6786
rect 8460 6786 8478 6804
rect 8460 6804 8478 6822
rect 8460 6822 8478 6840
rect 8460 6840 8478 6858
rect 8460 6858 8478 6876
rect 8460 6876 8478 6894
rect 8460 6894 8478 6912
rect 8460 6912 8478 6930
rect 8460 6930 8478 6948
rect 8460 6948 8478 6966
rect 8460 6966 8478 6984
rect 8460 6984 8478 7002
rect 8460 7002 8478 7020
rect 8460 7020 8478 7038
rect 8460 7038 8478 7056
rect 8460 7056 8478 7074
rect 8460 7074 8478 7092
rect 8460 7092 8478 7110
rect 8460 7110 8478 7128
rect 8460 7128 8478 7146
rect 8460 7146 8478 7164
rect 8460 7164 8478 7182
rect 8460 7182 8478 7200
rect 8460 7200 8478 7218
rect 8460 7218 8478 7236
rect 8460 7236 8478 7254
rect 8460 7254 8478 7272
rect 8460 7272 8478 7290
rect 8460 7290 8478 7308
rect 8460 7308 8478 7326
rect 8460 7326 8478 7344
rect 8478 2772 8496 2790
rect 8478 2790 8496 2808
rect 8478 2808 8496 2826
rect 8478 2826 8496 2844
rect 8478 2844 8496 2862
rect 8478 2862 8496 2880
rect 8478 2880 8496 2898
rect 8478 2898 8496 2916
rect 8478 2916 8496 2934
rect 8478 2934 8496 2952
rect 8478 2952 8496 2970
rect 8478 2970 8496 2988
rect 8478 2988 8496 3006
rect 8478 3006 8496 3024
rect 8478 3024 8496 3042
rect 8478 3042 8496 3060
rect 8478 3060 8496 3078
rect 8478 3078 8496 3096
rect 8478 3096 8496 3114
rect 8478 3114 8496 3132
rect 8478 3132 8496 3150
rect 8478 3150 8496 3168
rect 8478 3168 8496 3186
rect 8478 3186 8496 3204
rect 8478 3204 8496 3222
rect 8478 3222 8496 3240
rect 8478 3240 8496 3258
rect 8478 3258 8496 3276
rect 8478 3276 8496 3294
rect 8478 3294 8496 3312
rect 8478 3312 8496 3330
rect 8478 3330 8496 3348
rect 8478 3348 8496 3366
rect 8478 3366 8496 3384
rect 8478 3384 8496 3402
rect 8478 3402 8496 3420
rect 8478 3420 8496 3438
rect 8478 3438 8496 3456
rect 8478 3456 8496 3474
rect 8478 3474 8496 3492
rect 8478 5958 8496 5976
rect 8478 5976 8496 5994
rect 8478 5994 8496 6012
rect 8478 6012 8496 6030
rect 8478 6030 8496 6048
rect 8478 6048 8496 6066
rect 8478 6066 8496 6084
rect 8478 6084 8496 6102
rect 8478 6102 8496 6120
rect 8478 6120 8496 6138
rect 8478 6138 8496 6156
rect 8478 6156 8496 6174
rect 8478 6174 8496 6192
rect 8478 6192 8496 6210
rect 8478 6210 8496 6228
rect 8478 6228 8496 6246
rect 8478 6246 8496 6264
rect 8478 6264 8496 6282
rect 8478 6282 8496 6300
rect 8478 6300 8496 6318
rect 8478 6318 8496 6336
rect 8478 6336 8496 6354
rect 8478 6354 8496 6372
rect 8478 6372 8496 6390
rect 8478 6390 8496 6408
rect 8478 6408 8496 6426
rect 8478 6426 8496 6444
rect 8478 6444 8496 6462
rect 8478 6462 8496 6480
rect 8478 6480 8496 6498
rect 8478 6498 8496 6516
rect 8478 6516 8496 6534
rect 8478 6534 8496 6552
rect 8478 6552 8496 6570
rect 8478 6570 8496 6588
rect 8478 6588 8496 6606
rect 8478 6606 8496 6624
rect 8478 6624 8496 6642
rect 8478 6642 8496 6660
rect 8478 6660 8496 6678
rect 8478 6678 8496 6696
rect 8478 6696 8496 6714
rect 8478 6714 8496 6732
rect 8478 6732 8496 6750
rect 8478 6750 8496 6768
rect 8478 6768 8496 6786
rect 8478 6786 8496 6804
rect 8478 6804 8496 6822
rect 8478 6822 8496 6840
rect 8478 6840 8496 6858
rect 8478 6858 8496 6876
rect 8478 6876 8496 6894
rect 8478 6894 8496 6912
rect 8478 6912 8496 6930
rect 8478 6930 8496 6948
rect 8478 6948 8496 6966
rect 8478 6966 8496 6984
rect 8478 6984 8496 7002
rect 8478 7002 8496 7020
rect 8478 7020 8496 7038
rect 8478 7038 8496 7056
rect 8478 7056 8496 7074
rect 8478 7074 8496 7092
rect 8478 7092 8496 7110
rect 8478 7110 8496 7128
rect 8478 7128 8496 7146
rect 8478 7146 8496 7164
rect 8478 7164 8496 7182
rect 8478 7182 8496 7200
rect 8478 7200 8496 7218
rect 8478 7218 8496 7236
rect 8478 7236 8496 7254
rect 8478 7254 8496 7272
rect 8478 7272 8496 7290
rect 8478 7290 8496 7308
rect 8478 7308 8496 7326
rect 8478 7326 8496 7344
rect 8496 2790 8514 2808
rect 8496 2808 8514 2826
rect 8496 2826 8514 2844
rect 8496 2844 8514 2862
rect 8496 2862 8514 2880
rect 8496 2880 8514 2898
rect 8496 2898 8514 2916
rect 8496 2916 8514 2934
rect 8496 2934 8514 2952
rect 8496 2952 8514 2970
rect 8496 2970 8514 2988
rect 8496 2988 8514 3006
rect 8496 3006 8514 3024
rect 8496 3024 8514 3042
rect 8496 3042 8514 3060
rect 8496 3060 8514 3078
rect 8496 3078 8514 3096
rect 8496 3096 8514 3114
rect 8496 3114 8514 3132
rect 8496 3132 8514 3150
rect 8496 3150 8514 3168
rect 8496 3168 8514 3186
rect 8496 3186 8514 3204
rect 8496 3204 8514 3222
rect 8496 3222 8514 3240
rect 8496 3240 8514 3258
rect 8496 3258 8514 3276
rect 8496 3276 8514 3294
rect 8496 3294 8514 3312
rect 8496 3312 8514 3330
rect 8496 3330 8514 3348
rect 8496 3348 8514 3366
rect 8496 3366 8514 3384
rect 8496 3384 8514 3402
rect 8496 3402 8514 3420
rect 8496 3420 8514 3438
rect 8496 3438 8514 3456
rect 8496 3456 8514 3474
rect 8496 3474 8514 3492
rect 8496 5976 8514 5994
rect 8496 5994 8514 6012
rect 8496 6012 8514 6030
rect 8496 6030 8514 6048
rect 8496 6048 8514 6066
rect 8496 6066 8514 6084
rect 8496 6084 8514 6102
rect 8496 6102 8514 6120
rect 8496 6120 8514 6138
rect 8496 6138 8514 6156
rect 8496 6156 8514 6174
rect 8496 6174 8514 6192
rect 8496 6192 8514 6210
rect 8496 6210 8514 6228
rect 8496 6228 8514 6246
rect 8496 6246 8514 6264
rect 8496 6264 8514 6282
rect 8496 6282 8514 6300
rect 8496 6300 8514 6318
rect 8496 6318 8514 6336
rect 8496 6336 8514 6354
rect 8496 6354 8514 6372
rect 8496 6372 8514 6390
rect 8496 6390 8514 6408
rect 8496 6408 8514 6426
rect 8496 6426 8514 6444
rect 8496 6444 8514 6462
rect 8496 6462 8514 6480
rect 8496 6480 8514 6498
rect 8496 6498 8514 6516
rect 8496 6516 8514 6534
rect 8496 6534 8514 6552
rect 8496 6552 8514 6570
rect 8496 6570 8514 6588
rect 8496 6588 8514 6606
rect 8496 6606 8514 6624
rect 8496 6624 8514 6642
rect 8496 6642 8514 6660
rect 8496 6660 8514 6678
rect 8496 6678 8514 6696
rect 8496 6696 8514 6714
rect 8496 6714 8514 6732
rect 8496 6732 8514 6750
rect 8496 6750 8514 6768
rect 8496 6768 8514 6786
rect 8496 6786 8514 6804
rect 8496 6804 8514 6822
rect 8496 6822 8514 6840
rect 8496 6840 8514 6858
rect 8496 6858 8514 6876
rect 8496 6876 8514 6894
rect 8496 6894 8514 6912
rect 8496 6912 8514 6930
rect 8496 6930 8514 6948
rect 8496 6948 8514 6966
rect 8496 6966 8514 6984
rect 8496 6984 8514 7002
rect 8496 7002 8514 7020
rect 8496 7020 8514 7038
rect 8496 7038 8514 7056
rect 8496 7056 8514 7074
rect 8496 7074 8514 7092
rect 8496 7092 8514 7110
rect 8496 7110 8514 7128
rect 8496 7128 8514 7146
rect 8496 7146 8514 7164
rect 8496 7164 8514 7182
rect 8496 7182 8514 7200
rect 8496 7200 8514 7218
rect 8496 7218 8514 7236
rect 8496 7236 8514 7254
rect 8496 7254 8514 7272
rect 8496 7272 8514 7290
rect 8496 7290 8514 7308
rect 8496 7308 8514 7326
rect 8496 7326 8514 7344
rect 8496 7344 8514 7362
rect 8514 2808 8532 2826
rect 8514 2826 8532 2844
rect 8514 2844 8532 2862
rect 8514 2862 8532 2880
rect 8514 2880 8532 2898
rect 8514 2898 8532 2916
rect 8514 2916 8532 2934
rect 8514 2934 8532 2952
rect 8514 2952 8532 2970
rect 8514 2970 8532 2988
rect 8514 2988 8532 3006
rect 8514 3006 8532 3024
rect 8514 3024 8532 3042
rect 8514 3042 8532 3060
rect 8514 3060 8532 3078
rect 8514 3078 8532 3096
rect 8514 3096 8532 3114
rect 8514 3114 8532 3132
rect 8514 3132 8532 3150
rect 8514 3150 8532 3168
rect 8514 3168 8532 3186
rect 8514 3186 8532 3204
rect 8514 3204 8532 3222
rect 8514 3222 8532 3240
rect 8514 3240 8532 3258
rect 8514 3258 8532 3276
rect 8514 3276 8532 3294
rect 8514 3294 8532 3312
rect 8514 3312 8532 3330
rect 8514 3330 8532 3348
rect 8514 3348 8532 3366
rect 8514 3366 8532 3384
rect 8514 3384 8532 3402
rect 8514 3402 8532 3420
rect 8514 3420 8532 3438
rect 8514 3438 8532 3456
rect 8514 3456 8532 3474
rect 8514 3474 8532 3492
rect 8514 6012 8532 6030
rect 8514 6030 8532 6048
rect 8514 6048 8532 6066
rect 8514 6066 8532 6084
rect 8514 6084 8532 6102
rect 8514 6102 8532 6120
rect 8514 6120 8532 6138
rect 8514 6138 8532 6156
rect 8514 6156 8532 6174
rect 8514 6174 8532 6192
rect 8514 6192 8532 6210
rect 8514 6210 8532 6228
rect 8514 6228 8532 6246
rect 8514 6246 8532 6264
rect 8514 6264 8532 6282
rect 8514 6282 8532 6300
rect 8514 6300 8532 6318
rect 8514 6318 8532 6336
rect 8514 6336 8532 6354
rect 8514 6354 8532 6372
rect 8514 6372 8532 6390
rect 8514 6390 8532 6408
rect 8514 6408 8532 6426
rect 8514 6426 8532 6444
rect 8514 6444 8532 6462
rect 8514 6462 8532 6480
rect 8514 6480 8532 6498
rect 8514 6498 8532 6516
rect 8514 6516 8532 6534
rect 8514 6534 8532 6552
rect 8514 6552 8532 6570
rect 8514 6570 8532 6588
rect 8514 6588 8532 6606
rect 8514 6606 8532 6624
rect 8514 6624 8532 6642
rect 8514 6642 8532 6660
rect 8514 6660 8532 6678
rect 8514 6678 8532 6696
rect 8514 6696 8532 6714
rect 8514 6714 8532 6732
rect 8514 6732 8532 6750
rect 8514 6750 8532 6768
rect 8514 6768 8532 6786
rect 8514 6786 8532 6804
rect 8514 6804 8532 6822
rect 8514 6822 8532 6840
rect 8514 6840 8532 6858
rect 8514 6858 8532 6876
rect 8514 6876 8532 6894
rect 8514 6894 8532 6912
rect 8514 6912 8532 6930
rect 8514 6930 8532 6948
rect 8514 6948 8532 6966
rect 8514 6966 8532 6984
rect 8514 6984 8532 7002
rect 8514 7002 8532 7020
rect 8514 7020 8532 7038
rect 8514 7038 8532 7056
rect 8514 7056 8532 7074
rect 8514 7074 8532 7092
rect 8514 7092 8532 7110
rect 8514 7110 8532 7128
rect 8514 7128 8532 7146
rect 8514 7146 8532 7164
rect 8514 7164 8532 7182
rect 8514 7182 8532 7200
rect 8514 7200 8532 7218
rect 8514 7218 8532 7236
rect 8514 7236 8532 7254
rect 8514 7254 8532 7272
rect 8514 7272 8532 7290
rect 8514 7290 8532 7308
rect 8514 7308 8532 7326
rect 8514 7326 8532 7344
rect 8514 7344 8532 7362
rect 8514 7362 8532 7380
rect 8532 2826 8550 2844
rect 8532 2844 8550 2862
rect 8532 2862 8550 2880
rect 8532 2880 8550 2898
rect 8532 2898 8550 2916
rect 8532 2916 8550 2934
rect 8532 2934 8550 2952
rect 8532 2952 8550 2970
rect 8532 2970 8550 2988
rect 8532 2988 8550 3006
rect 8532 3006 8550 3024
rect 8532 3024 8550 3042
rect 8532 3042 8550 3060
rect 8532 3060 8550 3078
rect 8532 3078 8550 3096
rect 8532 3096 8550 3114
rect 8532 3114 8550 3132
rect 8532 3132 8550 3150
rect 8532 3150 8550 3168
rect 8532 3168 8550 3186
rect 8532 3186 8550 3204
rect 8532 3204 8550 3222
rect 8532 3222 8550 3240
rect 8532 3240 8550 3258
rect 8532 3258 8550 3276
rect 8532 3276 8550 3294
rect 8532 3294 8550 3312
rect 8532 3312 8550 3330
rect 8532 3330 8550 3348
rect 8532 3348 8550 3366
rect 8532 3366 8550 3384
rect 8532 3384 8550 3402
rect 8532 3402 8550 3420
rect 8532 3420 8550 3438
rect 8532 3438 8550 3456
rect 8532 3456 8550 3474
rect 8532 3474 8550 3492
rect 8532 6048 8550 6066
rect 8532 6066 8550 6084
rect 8532 6084 8550 6102
rect 8532 6102 8550 6120
rect 8532 6120 8550 6138
rect 8532 6138 8550 6156
rect 8532 6156 8550 6174
rect 8532 6174 8550 6192
rect 8532 6192 8550 6210
rect 8532 6210 8550 6228
rect 8532 6228 8550 6246
rect 8532 6246 8550 6264
rect 8532 6264 8550 6282
rect 8532 6282 8550 6300
rect 8532 6300 8550 6318
rect 8532 6318 8550 6336
rect 8532 6336 8550 6354
rect 8532 6354 8550 6372
rect 8532 6372 8550 6390
rect 8532 6390 8550 6408
rect 8532 6408 8550 6426
rect 8532 6426 8550 6444
rect 8532 6444 8550 6462
rect 8532 6462 8550 6480
rect 8532 6480 8550 6498
rect 8532 6498 8550 6516
rect 8532 6516 8550 6534
rect 8532 6534 8550 6552
rect 8532 6552 8550 6570
rect 8532 6570 8550 6588
rect 8532 6588 8550 6606
rect 8532 6606 8550 6624
rect 8532 6624 8550 6642
rect 8532 6642 8550 6660
rect 8532 6660 8550 6678
rect 8532 6678 8550 6696
rect 8532 6696 8550 6714
rect 8532 6714 8550 6732
rect 8532 6732 8550 6750
rect 8532 6750 8550 6768
rect 8532 6768 8550 6786
rect 8532 6786 8550 6804
rect 8532 6804 8550 6822
rect 8532 6822 8550 6840
rect 8532 6840 8550 6858
rect 8532 6858 8550 6876
rect 8532 6876 8550 6894
rect 8532 6894 8550 6912
rect 8532 6912 8550 6930
rect 8532 6930 8550 6948
rect 8532 6948 8550 6966
rect 8532 6966 8550 6984
rect 8532 6984 8550 7002
rect 8532 7002 8550 7020
rect 8532 7020 8550 7038
rect 8532 7038 8550 7056
rect 8532 7056 8550 7074
rect 8532 7074 8550 7092
rect 8532 7092 8550 7110
rect 8532 7110 8550 7128
rect 8532 7128 8550 7146
rect 8532 7146 8550 7164
rect 8532 7164 8550 7182
rect 8532 7182 8550 7200
rect 8532 7200 8550 7218
rect 8532 7218 8550 7236
rect 8532 7236 8550 7254
rect 8532 7254 8550 7272
rect 8532 7272 8550 7290
rect 8532 7290 8550 7308
rect 8532 7308 8550 7326
rect 8532 7326 8550 7344
rect 8532 7344 8550 7362
rect 8532 7362 8550 7380
rect 8550 2844 8568 2862
rect 8550 2862 8568 2880
rect 8550 2880 8568 2898
rect 8550 2898 8568 2916
rect 8550 2916 8568 2934
rect 8550 2934 8568 2952
rect 8550 2952 8568 2970
rect 8550 2970 8568 2988
rect 8550 2988 8568 3006
rect 8550 3006 8568 3024
rect 8550 3024 8568 3042
rect 8550 3042 8568 3060
rect 8550 3060 8568 3078
rect 8550 3078 8568 3096
rect 8550 3096 8568 3114
rect 8550 3114 8568 3132
rect 8550 3132 8568 3150
rect 8550 3150 8568 3168
rect 8550 3168 8568 3186
rect 8550 3186 8568 3204
rect 8550 3204 8568 3222
rect 8550 3222 8568 3240
rect 8550 3240 8568 3258
rect 8550 3258 8568 3276
rect 8550 3276 8568 3294
rect 8550 3294 8568 3312
rect 8550 3312 8568 3330
rect 8550 3330 8568 3348
rect 8550 3348 8568 3366
rect 8550 3366 8568 3384
rect 8550 3384 8568 3402
rect 8550 3402 8568 3420
rect 8550 3420 8568 3438
rect 8550 3438 8568 3456
rect 8550 3456 8568 3474
rect 8550 3474 8568 3492
rect 8550 3492 8568 3510
rect 8550 6066 8568 6084
rect 8550 6084 8568 6102
rect 8550 6102 8568 6120
rect 8550 6120 8568 6138
rect 8550 6138 8568 6156
rect 8550 6156 8568 6174
rect 8550 6174 8568 6192
rect 8550 6192 8568 6210
rect 8550 6210 8568 6228
rect 8550 6228 8568 6246
rect 8550 6246 8568 6264
rect 8550 6264 8568 6282
rect 8550 6282 8568 6300
rect 8550 6300 8568 6318
rect 8550 6318 8568 6336
rect 8550 6336 8568 6354
rect 8550 6354 8568 6372
rect 8550 6372 8568 6390
rect 8550 6390 8568 6408
rect 8550 6408 8568 6426
rect 8550 6426 8568 6444
rect 8550 6444 8568 6462
rect 8550 6462 8568 6480
rect 8550 6480 8568 6498
rect 8550 6498 8568 6516
rect 8550 6516 8568 6534
rect 8550 6534 8568 6552
rect 8550 6552 8568 6570
rect 8550 6570 8568 6588
rect 8550 6588 8568 6606
rect 8550 6606 8568 6624
rect 8550 6624 8568 6642
rect 8550 6642 8568 6660
rect 8550 6660 8568 6678
rect 8550 6678 8568 6696
rect 8550 6696 8568 6714
rect 8550 6714 8568 6732
rect 8550 6732 8568 6750
rect 8550 6750 8568 6768
rect 8550 6768 8568 6786
rect 8550 6786 8568 6804
rect 8550 6804 8568 6822
rect 8550 6822 8568 6840
rect 8550 6840 8568 6858
rect 8550 6858 8568 6876
rect 8550 6876 8568 6894
rect 8550 6894 8568 6912
rect 8550 6912 8568 6930
rect 8550 6930 8568 6948
rect 8550 6948 8568 6966
rect 8550 6966 8568 6984
rect 8550 6984 8568 7002
rect 8550 7002 8568 7020
rect 8550 7020 8568 7038
rect 8550 7038 8568 7056
rect 8550 7056 8568 7074
rect 8550 7074 8568 7092
rect 8550 7092 8568 7110
rect 8550 7110 8568 7128
rect 8550 7128 8568 7146
rect 8550 7146 8568 7164
rect 8550 7164 8568 7182
rect 8550 7182 8568 7200
rect 8550 7200 8568 7218
rect 8550 7218 8568 7236
rect 8550 7236 8568 7254
rect 8550 7254 8568 7272
rect 8550 7272 8568 7290
rect 8550 7290 8568 7308
rect 8550 7308 8568 7326
rect 8550 7326 8568 7344
rect 8550 7344 8568 7362
rect 8550 7362 8568 7380
rect 8550 7380 8568 7398
rect 8568 2862 8586 2880
rect 8568 2880 8586 2898
rect 8568 2898 8586 2916
rect 8568 2916 8586 2934
rect 8568 2934 8586 2952
rect 8568 2952 8586 2970
rect 8568 2970 8586 2988
rect 8568 2988 8586 3006
rect 8568 3006 8586 3024
rect 8568 3024 8586 3042
rect 8568 3042 8586 3060
rect 8568 3060 8586 3078
rect 8568 3078 8586 3096
rect 8568 3096 8586 3114
rect 8568 3114 8586 3132
rect 8568 3132 8586 3150
rect 8568 3150 8586 3168
rect 8568 3168 8586 3186
rect 8568 3186 8586 3204
rect 8568 3204 8586 3222
rect 8568 3222 8586 3240
rect 8568 3240 8586 3258
rect 8568 3258 8586 3276
rect 8568 3276 8586 3294
rect 8568 3294 8586 3312
rect 8568 3312 8586 3330
rect 8568 3330 8586 3348
rect 8568 3348 8586 3366
rect 8568 3366 8586 3384
rect 8568 3384 8586 3402
rect 8568 3402 8586 3420
rect 8568 3420 8586 3438
rect 8568 3438 8586 3456
rect 8568 3456 8586 3474
rect 8568 3474 8586 3492
rect 8568 3492 8586 3510
rect 8568 6102 8586 6120
rect 8568 6120 8586 6138
rect 8568 6138 8586 6156
rect 8568 6156 8586 6174
rect 8568 6174 8586 6192
rect 8568 6192 8586 6210
rect 8568 6210 8586 6228
rect 8568 6228 8586 6246
rect 8568 6246 8586 6264
rect 8568 6264 8586 6282
rect 8568 6282 8586 6300
rect 8568 6300 8586 6318
rect 8568 6318 8586 6336
rect 8568 6336 8586 6354
rect 8568 6354 8586 6372
rect 8568 6372 8586 6390
rect 8568 6390 8586 6408
rect 8568 6408 8586 6426
rect 8568 6426 8586 6444
rect 8568 6444 8586 6462
rect 8568 6462 8586 6480
rect 8568 6480 8586 6498
rect 8568 6498 8586 6516
rect 8568 6516 8586 6534
rect 8568 6534 8586 6552
rect 8568 6552 8586 6570
rect 8568 6570 8586 6588
rect 8568 6588 8586 6606
rect 8568 6606 8586 6624
rect 8568 6624 8586 6642
rect 8568 6642 8586 6660
rect 8568 6660 8586 6678
rect 8568 6678 8586 6696
rect 8568 6696 8586 6714
rect 8568 6714 8586 6732
rect 8568 6732 8586 6750
rect 8568 6750 8586 6768
rect 8568 6768 8586 6786
rect 8568 6786 8586 6804
rect 8568 6804 8586 6822
rect 8568 6822 8586 6840
rect 8568 6840 8586 6858
rect 8568 6858 8586 6876
rect 8568 6876 8586 6894
rect 8568 6894 8586 6912
rect 8568 6912 8586 6930
rect 8568 6930 8586 6948
rect 8568 6948 8586 6966
rect 8568 6966 8586 6984
rect 8568 6984 8586 7002
rect 8568 7002 8586 7020
rect 8568 7020 8586 7038
rect 8568 7038 8586 7056
rect 8568 7056 8586 7074
rect 8568 7074 8586 7092
rect 8568 7092 8586 7110
rect 8568 7110 8586 7128
rect 8568 7128 8586 7146
rect 8568 7146 8586 7164
rect 8568 7164 8586 7182
rect 8568 7182 8586 7200
rect 8568 7200 8586 7218
rect 8568 7218 8586 7236
rect 8568 7236 8586 7254
rect 8568 7254 8586 7272
rect 8568 7272 8586 7290
rect 8568 7290 8586 7308
rect 8568 7308 8586 7326
rect 8568 7326 8586 7344
rect 8568 7344 8586 7362
rect 8568 7362 8586 7380
rect 8568 7380 8586 7398
rect 8586 2898 8604 2916
rect 8586 2916 8604 2934
rect 8586 2934 8604 2952
rect 8586 2952 8604 2970
rect 8586 2970 8604 2988
rect 8586 2988 8604 3006
rect 8586 3006 8604 3024
rect 8586 3024 8604 3042
rect 8586 3042 8604 3060
rect 8586 3060 8604 3078
rect 8586 3078 8604 3096
rect 8586 3096 8604 3114
rect 8586 3114 8604 3132
rect 8586 3132 8604 3150
rect 8586 3150 8604 3168
rect 8586 3168 8604 3186
rect 8586 3186 8604 3204
rect 8586 3204 8604 3222
rect 8586 3222 8604 3240
rect 8586 3240 8604 3258
rect 8586 3258 8604 3276
rect 8586 3276 8604 3294
rect 8586 3294 8604 3312
rect 8586 3312 8604 3330
rect 8586 3330 8604 3348
rect 8586 3348 8604 3366
rect 8586 3366 8604 3384
rect 8586 3384 8604 3402
rect 8586 3402 8604 3420
rect 8586 3420 8604 3438
rect 8586 3438 8604 3456
rect 8586 3456 8604 3474
rect 8586 3474 8604 3492
rect 8586 3492 8604 3510
rect 8586 6156 8604 6174
rect 8586 6174 8604 6192
rect 8586 6192 8604 6210
rect 8586 6210 8604 6228
rect 8586 6228 8604 6246
rect 8586 6246 8604 6264
rect 8586 6264 8604 6282
rect 8586 6282 8604 6300
rect 8586 6300 8604 6318
rect 8586 6318 8604 6336
rect 8586 6336 8604 6354
rect 8586 6354 8604 6372
rect 8586 6372 8604 6390
rect 8586 6390 8604 6408
rect 8586 6408 8604 6426
rect 8586 6426 8604 6444
rect 8586 6444 8604 6462
rect 8586 6462 8604 6480
rect 8586 6480 8604 6498
rect 8586 6498 8604 6516
rect 8586 6516 8604 6534
rect 8586 6534 8604 6552
rect 8586 6552 8604 6570
rect 8586 6570 8604 6588
rect 8586 6588 8604 6606
rect 8586 6606 8604 6624
rect 8586 6624 8604 6642
rect 8586 6642 8604 6660
rect 8586 6660 8604 6678
rect 8586 6678 8604 6696
rect 8586 6696 8604 6714
rect 8586 6714 8604 6732
rect 8586 6732 8604 6750
rect 8586 6750 8604 6768
rect 8586 6768 8604 6786
rect 8586 6786 8604 6804
rect 8586 6804 8604 6822
rect 8586 6822 8604 6840
rect 8586 6840 8604 6858
rect 8586 6858 8604 6876
rect 8586 6876 8604 6894
rect 8586 6894 8604 6912
rect 8586 6912 8604 6930
rect 8586 6930 8604 6948
rect 8586 6948 8604 6966
rect 8586 6966 8604 6984
rect 8586 6984 8604 7002
rect 8586 7002 8604 7020
rect 8586 7020 8604 7038
rect 8586 7038 8604 7056
rect 8586 7056 8604 7074
rect 8586 7074 8604 7092
rect 8586 7092 8604 7110
rect 8586 7110 8604 7128
rect 8586 7128 8604 7146
rect 8586 7146 8604 7164
rect 8586 7164 8604 7182
rect 8586 7182 8604 7200
rect 8586 7200 8604 7218
rect 8586 7218 8604 7236
rect 8586 7236 8604 7254
rect 8586 7254 8604 7272
rect 8586 7272 8604 7290
rect 8586 7290 8604 7308
rect 8586 7308 8604 7326
rect 8586 7326 8604 7344
rect 8586 7344 8604 7362
rect 8586 7362 8604 7380
rect 8586 7380 8604 7398
rect 8586 7398 8604 7416
rect 8604 2916 8622 2934
rect 8604 2934 8622 2952
rect 8604 2952 8622 2970
rect 8604 2970 8622 2988
rect 8604 2988 8622 3006
rect 8604 3006 8622 3024
rect 8604 3024 8622 3042
rect 8604 3042 8622 3060
rect 8604 3060 8622 3078
rect 8604 3078 8622 3096
rect 8604 3096 8622 3114
rect 8604 3114 8622 3132
rect 8604 3132 8622 3150
rect 8604 3150 8622 3168
rect 8604 3168 8622 3186
rect 8604 3186 8622 3204
rect 8604 3204 8622 3222
rect 8604 3222 8622 3240
rect 8604 3240 8622 3258
rect 8604 3258 8622 3276
rect 8604 3276 8622 3294
rect 8604 3294 8622 3312
rect 8604 3312 8622 3330
rect 8604 3330 8622 3348
rect 8604 3348 8622 3366
rect 8604 3366 8622 3384
rect 8604 3384 8622 3402
rect 8604 3402 8622 3420
rect 8604 3420 8622 3438
rect 8604 3438 8622 3456
rect 8604 3456 8622 3474
rect 8604 3474 8622 3492
rect 8604 3492 8622 3510
rect 8604 6192 8622 6210
rect 8604 6210 8622 6228
rect 8604 6228 8622 6246
rect 8604 6246 8622 6264
rect 8604 6264 8622 6282
rect 8604 6282 8622 6300
rect 8604 6300 8622 6318
rect 8604 6318 8622 6336
rect 8604 6336 8622 6354
rect 8604 6354 8622 6372
rect 8604 6372 8622 6390
rect 8604 6390 8622 6408
rect 8604 6408 8622 6426
rect 8604 6426 8622 6444
rect 8604 6444 8622 6462
rect 8604 6462 8622 6480
rect 8604 6480 8622 6498
rect 8604 6498 8622 6516
rect 8604 6516 8622 6534
rect 8604 6534 8622 6552
rect 8604 6552 8622 6570
rect 8604 6570 8622 6588
rect 8604 6588 8622 6606
rect 8604 6606 8622 6624
rect 8604 6624 8622 6642
rect 8604 6642 8622 6660
rect 8604 6660 8622 6678
rect 8604 6678 8622 6696
rect 8604 6696 8622 6714
rect 8604 6714 8622 6732
rect 8604 6732 8622 6750
rect 8604 6750 8622 6768
rect 8604 6768 8622 6786
rect 8604 6786 8622 6804
rect 8604 6804 8622 6822
rect 8604 6822 8622 6840
rect 8604 6840 8622 6858
rect 8604 6858 8622 6876
rect 8604 6876 8622 6894
rect 8604 6894 8622 6912
rect 8604 6912 8622 6930
rect 8604 6930 8622 6948
rect 8604 6948 8622 6966
rect 8604 6966 8622 6984
rect 8604 6984 8622 7002
rect 8604 7002 8622 7020
rect 8604 7020 8622 7038
rect 8604 7038 8622 7056
rect 8604 7056 8622 7074
rect 8604 7074 8622 7092
rect 8604 7092 8622 7110
rect 8604 7110 8622 7128
rect 8604 7128 8622 7146
rect 8604 7146 8622 7164
rect 8604 7164 8622 7182
rect 8604 7182 8622 7200
rect 8604 7200 8622 7218
rect 8604 7218 8622 7236
rect 8604 7236 8622 7254
rect 8604 7254 8622 7272
rect 8604 7272 8622 7290
rect 8604 7290 8622 7308
rect 8604 7308 8622 7326
rect 8604 7326 8622 7344
rect 8604 7344 8622 7362
rect 8604 7362 8622 7380
rect 8604 7380 8622 7398
rect 8604 7398 8622 7416
rect 8604 7416 8622 7434
rect 8622 2934 8640 2952
rect 8622 2952 8640 2970
rect 8622 2970 8640 2988
rect 8622 2988 8640 3006
rect 8622 3006 8640 3024
rect 8622 3024 8640 3042
rect 8622 3042 8640 3060
rect 8622 3060 8640 3078
rect 8622 3078 8640 3096
rect 8622 3096 8640 3114
rect 8622 3114 8640 3132
rect 8622 3132 8640 3150
rect 8622 3150 8640 3168
rect 8622 3168 8640 3186
rect 8622 3186 8640 3204
rect 8622 3204 8640 3222
rect 8622 3222 8640 3240
rect 8622 3240 8640 3258
rect 8622 3258 8640 3276
rect 8622 3276 8640 3294
rect 8622 3294 8640 3312
rect 8622 3312 8640 3330
rect 8622 3330 8640 3348
rect 8622 3348 8640 3366
rect 8622 3366 8640 3384
rect 8622 3384 8640 3402
rect 8622 3402 8640 3420
rect 8622 3420 8640 3438
rect 8622 3438 8640 3456
rect 8622 3456 8640 3474
rect 8622 3474 8640 3492
rect 8622 3492 8640 3510
rect 8622 3510 8640 3528
rect 8622 6228 8640 6246
rect 8622 6246 8640 6264
rect 8622 6264 8640 6282
rect 8622 6282 8640 6300
rect 8622 6300 8640 6318
rect 8622 6318 8640 6336
rect 8622 6336 8640 6354
rect 8622 6354 8640 6372
rect 8622 6372 8640 6390
rect 8622 6390 8640 6408
rect 8622 6408 8640 6426
rect 8622 6426 8640 6444
rect 8622 6444 8640 6462
rect 8622 6462 8640 6480
rect 8622 6480 8640 6498
rect 8622 6498 8640 6516
rect 8622 6516 8640 6534
rect 8622 6534 8640 6552
rect 8622 6552 8640 6570
rect 8622 6570 8640 6588
rect 8622 6588 8640 6606
rect 8622 6606 8640 6624
rect 8622 6624 8640 6642
rect 8622 6642 8640 6660
rect 8622 6660 8640 6678
rect 8622 6678 8640 6696
rect 8622 6696 8640 6714
rect 8622 6714 8640 6732
rect 8622 6732 8640 6750
rect 8622 6750 8640 6768
rect 8622 6768 8640 6786
rect 8622 6786 8640 6804
rect 8622 6804 8640 6822
rect 8622 6822 8640 6840
rect 8622 6840 8640 6858
rect 8622 6858 8640 6876
rect 8622 6876 8640 6894
rect 8622 6894 8640 6912
rect 8622 6912 8640 6930
rect 8622 6930 8640 6948
rect 8622 6948 8640 6966
rect 8622 6966 8640 6984
rect 8622 6984 8640 7002
rect 8622 7002 8640 7020
rect 8622 7020 8640 7038
rect 8622 7038 8640 7056
rect 8622 7056 8640 7074
rect 8622 7074 8640 7092
rect 8622 7092 8640 7110
rect 8622 7110 8640 7128
rect 8622 7128 8640 7146
rect 8622 7146 8640 7164
rect 8622 7164 8640 7182
rect 8622 7182 8640 7200
rect 8622 7200 8640 7218
rect 8622 7218 8640 7236
rect 8622 7236 8640 7254
rect 8622 7254 8640 7272
rect 8622 7272 8640 7290
rect 8622 7290 8640 7308
rect 8622 7308 8640 7326
rect 8622 7326 8640 7344
rect 8622 7344 8640 7362
rect 8622 7362 8640 7380
rect 8622 7380 8640 7398
rect 8622 7398 8640 7416
rect 8622 7416 8640 7434
rect 8640 2952 8658 2970
rect 8640 2970 8658 2988
rect 8640 2988 8658 3006
rect 8640 3006 8658 3024
rect 8640 3024 8658 3042
rect 8640 3042 8658 3060
rect 8640 3060 8658 3078
rect 8640 3078 8658 3096
rect 8640 3096 8658 3114
rect 8640 3114 8658 3132
rect 8640 3132 8658 3150
rect 8640 3150 8658 3168
rect 8640 3168 8658 3186
rect 8640 3186 8658 3204
rect 8640 3204 8658 3222
rect 8640 3222 8658 3240
rect 8640 3240 8658 3258
rect 8640 3258 8658 3276
rect 8640 3276 8658 3294
rect 8640 3294 8658 3312
rect 8640 3312 8658 3330
rect 8640 3330 8658 3348
rect 8640 3348 8658 3366
rect 8640 3366 8658 3384
rect 8640 3384 8658 3402
rect 8640 3402 8658 3420
rect 8640 3420 8658 3438
rect 8640 3438 8658 3456
rect 8640 3456 8658 3474
rect 8640 3474 8658 3492
rect 8640 3492 8658 3510
rect 8640 3510 8658 3528
rect 8640 6282 8658 6300
rect 8640 6300 8658 6318
rect 8640 6318 8658 6336
rect 8640 6336 8658 6354
rect 8640 6354 8658 6372
rect 8640 6372 8658 6390
rect 8640 6390 8658 6408
rect 8640 6408 8658 6426
rect 8640 6426 8658 6444
rect 8640 6444 8658 6462
rect 8640 6462 8658 6480
rect 8640 6480 8658 6498
rect 8640 6498 8658 6516
rect 8640 6516 8658 6534
rect 8640 6534 8658 6552
rect 8640 6552 8658 6570
rect 8640 6570 8658 6588
rect 8640 6588 8658 6606
rect 8640 6606 8658 6624
rect 8640 6624 8658 6642
rect 8640 6642 8658 6660
rect 8640 6660 8658 6678
rect 8640 6678 8658 6696
rect 8640 6696 8658 6714
rect 8640 6714 8658 6732
rect 8640 6732 8658 6750
rect 8640 6750 8658 6768
rect 8640 6768 8658 6786
rect 8640 6786 8658 6804
rect 8640 6804 8658 6822
rect 8640 6822 8658 6840
rect 8640 6840 8658 6858
rect 8640 6858 8658 6876
rect 8640 6876 8658 6894
rect 8640 6894 8658 6912
rect 8640 6912 8658 6930
rect 8640 6930 8658 6948
rect 8640 6948 8658 6966
rect 8640 6966 8658 6984
rect 8640 6984 8658 7002
rect 8640 7002 8658 7020
rect 8640 7020 8658 7038
rect 8640 7038 8658 7056
rect 8640 7056 8658 7074
rect 8640 7074 8658 7092
rect 8640 7092 8658 7110
rect 8640 7110 8658 7128
rect 8640 7128 8658 7146
rect 8640 7146 8658 7164
rect 8640 7164 8658 7182
rect 8640 7182 8658 7200
rect 8640 7200 8658 7218
rect 8640 7218 8658 7236
rect 8640 7236 8658 7254
rect 8640 7254 8658 7272
rect 8640 7272 8658 7290
rect 8640 7290 8658 7308
rect 8640 7308 8658 7326
rect 8640 7326 8658 7344
rect 8640 7344 8658 7362
rect 8640 7362 8658 7380
rect 8640 7380 8658 7398
rect 8640 7398 8658 7416
rect 8640 7416 8658 7434
rect 8640 7434 8658 7452
rect 8658 2970 8676 2988
rect 8658 2988 8676 3006
rect 8658 3006 8676 3024
rect 8658 3024 8676 3042
rect 8658 3042 8676 3060
rect 8658 3060 8676 3078
rect 8658 3078 8676 3096
rect 8658 3096 8676 3114
rect 8658 3114 8676 3132
rect 8658 3132 8676 3150
rect 8658 3150 8676 3168
rect 8658 3168 8676 3186
rect 8658 3186 8676 3204
rect 8658 3204 8676 3222
rect 8658 3222 8676 3240
rect 8658 3240 8676 3258
rect 8658 3258 8676 3276
rect 8658 3276 8676 3294
rect 8658 3294 8676 3312
rect 8658 3312 8676 3330
rect 8658 3330 8676 3348
rect 8658 3348 8676 3366
rect 8658 3366 8676 3384
rect 8658 3384 8676 3402
rect 8658 3402 8676 3420
rect 8658 3420 8676 3438
rect 8658 3438 8676 3456
rect 8658 3456 8676 3474
rect 8658 3474 8676 3492
rect 8658 3492 8676 3510
rect 8658 3510 8676 3528
rect 8658 6318 8676 6336
rect 8658 6336 8676 6354
rect 8658 6354 8676 6372
rect 8658 6372 8676 6390
rect 8658 6390 8676 6408
rect 8658 6408 8676 6426
rect 8658 6426 8676 6444
rect 8658 6444 8676 6462
rect 8658 6462 8676 6480
rect 8658 6480 8676 6498
rect 8658 6498 8676 6516
rect 8658 6516 8676 6534
rect 8658 6534 8676 6552
rect 8658 6552 8676 6570
rect 8658 6570 8676 6588
rect 8658 6588 8676 6606
rect 8658 6606 8676 6624
rect 8658 6624 8676 6642
rect 8658 6642 8676 6660
rect 8658 6660 8676 6678
rect 8658 6678 8676 6696
rect 8658 6696 8676 6714
rect 8658 6714 8676 6732
rect 8658 6732 8676 6750
rect 8658 6750 8676 6768
rect 8658 6768 8676 6786
rect 8658 6786 8676 6804
rect 8658 6804 8676 6822
rect 8658 6822 8676 6840
rect 8658 6840 8676 6858
rect 8658 6858 8676 6876
rect 8658 6876 8676 6894
rect 8658 6894 8676 6912
rect 8658 6912 8676 6930
rect 8658 6930 8676 6948
rect 8658 6948 8676 6966
rect 8658 6966 8676 6984
rect 8658 6984 8676 7002
rect 8658 7002 8676 7020
rect 8658 7020 8676 7038
rect 8658 7038 8676 7056
rect 8658 7056 8676 7074
rect 8658 7074 8676 7092
rect 8658 7092 8676 7110
rect 8658 7110 8676 7128
rect 8658 7128 8676 7146
rect 8658 7146 8676 7164
rect 8658 7164 8676 7182
rect 8658 7182 8676 7200
rect 8658 7200 8676 7218
rect 8658 7218 8676 7236
rect 8658 7236 8676 7254
rect 8658 7254 8676 7272
rect 8658 7272 8676 7290
rect 8658 7290 8676 7308
rect 8658 7308 8676 7326
rect 8658 7326 8676 7344
rect 8658 7344 8676 7362
rect 8658 7362 8676 7380
rect 8658 7380 8676 7398
rect 8658 7398 8676 7416
rect 8658 7416 8676 7434
rect 8658 7434 8676 7452
rect 8658 7452 8676 7470
rect 8676 3006 8694 3024
rect 8676 3024 8694 3042
rect 8676 3042 8694 3060
rect 8676 3060 8694 3078
rect 8676 3078 8694 3096
rect 8676 3096 8694 3114
rect 8676 3114 8694 3132
rect 8676 3132 8694 3150
rect 8676 3150 8694 3168
rect 8676 3168 8694 3186
rect 8676 3186 8694 3204
rect 8676 3204 8694 3222
rect 8676 3222 8694 3240
rect 8676 3240 8694 3258
rect 8676 3258 8694 3276
rect 8676 3276 8694 3294
rect 8676 3294 8694 3312
rect 8676 3312 8694 3330
rect 8676 3330 8694 3348
rect 8676 3348 8694 3366
rect 8676 3366 8694 3384
rect 8676 3384 8694 3402
rect 8676 3402 8694 3420
rect 8676 3420 8694 3438
rect 8676 3438 8694 3456
rect 8676 3456 8694 3474
rect 8676 3474 8694 3492
rect 8676 3492 8694 3510
rect 8676 3510 8694 3528
rect 8676 6354 8694 6372
rect 8676 6372 8694 6390
rect 8676 6390 8694 6408
rect 8676 6408 8694 6426
rect 8676 6426 8694 6444
rect 8676 6444 8694 6462
rect 8676 6462 8694 6480
rect 8676 6480 8694 6498
rect 8676 6498 8694 6516
rect 8676 6516 8694 6534
rect 8676 6534 8694 6552
rect 8676 6552 8694 6570
rect 8676 6570 8694 6588
rect 8676 6588 8694 6606
rect 8676 6606 8694 6624
rect 8676 6624 8694 6642
rect 8676 6642 8694 6660
rect 8676 6660 8694 6678
rect 8676 6678 8694 6696
rect 8676 6696 8694 6714
rect 8676 6714 8694 6732
rect 8676 6732 8694 6750
rect 8676 6750 8694 6768
rect 8676 6768 8694 6786
rect 8676 6786 8694 6804
rect 8676 6804 8694 6822
rect 8676 6822 8694 6840
rect 8676 6840 8694 6858
rect 8676 6858 8694 6876
rect 8676 6876 8694 6894
rect 8676 6894 8694 6912
rect 8676 6912 8694 6930
rect 8676 6930 8694 6948
rect 8676 6948 8694 6966
rect 8676 6966 8694 6984
rect 8676 6984 8694 7002
rect 8676 7002 8694 7020
rect 8676 7020 8694 7038
rect 8676 7038 8694 7056
rect 8676 7056 8694 7074
rect 8676 7074 8694 7092
rect 8676 7092 8694 7110
rect 8676 7110 8694 7128
rect 8676 7128 8694 7146
rect 8676 7146 8694 7164
rect 8676 7164 8694 7182
rect 8676 7182 8694 7200
rect 8676 7200 8694 7218
rect 8676 7218 8694 7236
rect 8676 7236 8694 7254
rect 8676 7254 8694 7272
rect 8676 7272 8694 7290
rect 8676 7290 8694 7308
rect 8676 7308 8694 7326
rect 8676 7326 8694 7344
rect 8676 7344 8694 7362
rect 8676 7362 8694 7380
rect 8676 7380 8694 7398
rect 8676 7398 8694 7416
rect 8676 7416 8694 7434
rect 8676 7434 8694 7452
rect 8676 7452 8694 7470
rect 8694 3024 8712 3042
rect 8694 3042 8712 3060
rect 8694 3060 8712 3078
rect 8694 3078 8712 3096
rect 8694 3096 8712 3114
rect 8694 3114 8712 3132
rect 8694 3132 8712 3150
rect 8694 3150 8712 3168
rect 8694 3168 8712 3186
rect 8694 3186 8712 3204
rect 8694 3204 8712 3222
rect 8694 3222 8712 3240
rect 8694 3240 8712 3258
rect 8694 3258 8712 3276
rect 8694 3276 8712 3294
rect 8694 3294 8712 3312
rect 8694 3312 8712 3330
rect 8694 3330 8712 3348
rect 8694 3348 8712 3366
rect 8694 3366 8712 3384
rect 8694 3384 8712 3402
rect 8694 3402 8712 3420
rect 8694 3420 8712 3438
rect 8694 3438 8712 3456
rect 8694 3456 8712 3474
rect 8694 3474 8712 3492
rect 8694 3492 8712 3510
rect 8694 3510 8712 3528
rect 8694 6426 8712 6444
rect 8694 6444 8712 6462
rect 8694 6462 8712 6480
rect 8694 6480 8712 6498
rect 8694 6498 8712 6516
rect 8694 6516 8712 6534
rect 8694 6534 8712 6552
rect 8694 6552 8712 6570
rect 8694 6570 8712 6588
rect 8694 6588 8712 6606
rect 8694 6606 8712 6624
rect 8694 6624 8712 6642
rect 8694 6642 8712 6660
rect 8694 6660 8712 6678
rect 8694 6678 8712 6696
rect 8694 6696 8712 6714
rect 8694 6714 8712 6732
rect 8694 6732 8712 6750
rect 8694 6750 8712 6768
rect 8694 6768 8712 6786
rect 8694 6786 8712 6804
rect 8694 6804 8712 6822
rect 8694 6822 8712 6840
rect 8694 6840 8712 6858
rect 8694 6858 8712 6876
rect 8694 6876 8712 6894
rect 8694 6894 8712 6912
rect 8694 6912 8712 6930
rect 8694 6930 8712 6948
rect 8694 6948 8712 6966
rect 8694 6966 8712 6984
rect 8694 6984 8712 7002
rect 8694 7002 8712 7020
rect 8694 7020 8712 7038
rect 8694 7038 8712 7056
rect 8694 7056 8712 7074
rect 8694 7074 8712 7092
rect 8694 7092 8712 7110
rect 8694 7110 8712 7128
rect 8694 7128 8712 7146
rect 8694 7146 8712 7164
rect 8694 7164 8712 7182
rect 8694 7182 8712 7200
rect 8694 7200 8712 7218
rect 8694 7218 8712 7236
rect 8694 7236 8712 7254
rect 8694 7254 8712 7272
rect 8694 7272 8712 7290
rect 8694 7290 8712 7308
rect 8694 7308 8712 7326
rect 8694 7326 8712 7344
rect 8694 7344 8712 7362
rect 8694 7362 8712 7380
rect 8694 7380 8712 7398
rect 8694 7398 8712 7416
rect 8694 7416 8712 7434
rect 8694 7434 8712 7452
rect 8694 7452 8712 7470
rect 8694 7470 8712 7488
rect 8712 3042 8730 3060
rect 8712 3060 8730 3078
rect 8712 3078 8730 3096
rect 8712 3096 8730 3114
rect 8712 3114 8730 3132
rect 8712 3132 8730 3150
rect 8712 3150 8730 3168
rect 8712 3168 8730 3186
rect 8712 3186 8730 3204
rect 8712 3204 8730 3222
rect 8712 3222 8730 3240
rect 8712 3240 8730 3258
rect 8712 3258 8730 3276
rect 8712 3276 8730 3294
rect 8712 3294 8730 3312
rect 8712 3312 8730 3330
rect 8712 3330 8730 3348
rect 8712 3348 8730 3366
rect 8712 3366 8730 3384
rect 8712 3384 8730 3402
rect 8712 3402 8730 3420
rect 8712 3420 8730 3438
rect 8712 3438 8730 3456
rect 8712 3456 8730 3474
rect 8712 3474 8730 3492
rect 8712 3492 8730 3510
rect 8712 3510 8730 3528
rect 8712 3528 8730 3546
rect 8712 6498 8730 6516
rect 8712 6516 8730 6534
rect 8712 6534 8730 6552
rect 8712 6552 8730 6570
rect 8712 6570 8730 6588
rect 8712 6588 8730 6606
rect 8712 6606 8730 6624
rect 8712 6624 8730 6642
rect 8712 6642 8730 6660
rect 8712 6660 8730 6678
rect 8712 6678 8730 6696
rect 8712 6696 8730 6714
rect 8712 6714 8730 6732
rect 8712 6732 8730 6750
rect 8712 6750 8730 6768
rect 8712 6768 8730 6786
rect 8712 6786 8730 6804
rect 8712 6804 8730 6822
rect 8712 6822 8730 6840
rect 8712 6840 8730 6858
rect 8712 6858 8730 6876
rect 8712 6876 8730 6894
rect 8712 6894 8730 6912
rect 8712 6912 8730 6930
rect 8712 6930 8730 6948
rect 8712 6948 8730 6966
rect 8712 6966 8730 6984
rect 8712 6984 8730 7002
rect 8712 7002 8730 7020
rect 8712 7020 8730 7038
rect 8712 7038 8730 7056
rect 8712 7056 8730 7074
rect 8712 7074 8730 7092
rect 8712 7092 8730 7110
rect 8712 7110 8730 7128
rect 8712 7128 8730 7146
rect 8712 7146 8730 7164
rect 8712 7164 8730 7182
rect 8712 7182 8730 7200
rect 8712 7200 8730 7218
rect 8712 7218 8730 7236
rect 8712 7236 8730 7254
rect 8712 7254 8730 7272
rect 8712 7272 8730 7290
rect 8712 7290 8730 7308
rect 8712 7308 8730 7326
rect 8712 7326 8730 7344
rect 8712 7344 8730 7362
rect 8712 7362 8730 7380
rect 8712 7380 8730 7398
rect 8712 7398 8730 7416
rect 8712 7416 8730 7434
rect 8712 7434 8730 7452
rect 8712 7452 8730 7470
rect 8712 7470 8730 7488
rect 8712 7488 8730 7506
rect 8730 3060 8748 3078
rect 8730 3078 8748 3096
rect 8730 3096 8748 3114
rect 8730 3114 8748 3132
rect 8730 3132 8748 3150
rect 8730 3150 8748 3168
rect 8730 3168 8748 3186
rect 8730 3186 8748 3204
rect 8730 3204 8748 3222
rect 8730 3222 8748 3240
rect 8730 3240 8748 3258
rect 8730 3258 8748 3276
rect 8730 3276 8748 3294
rect 8730 3294 8748 3312
rect 8730 3312 8748 3330
rect 8730 3330 8748 3348
rect 8730 3348 8748 3366
rect 8730 3366 8748 3384
rect 8730 3384 8748 3402
rect 8730 3402 8748 3420
rect 8730 3420 8748 3438
rect 8730 3438 8748 3456
rect 8730 3456 8748 3474
rect 8730 3474 8748 3492
rect 8730 3492 8748 3510
rect 8730 3510 8748 3528
rect 8730 3528 8748 3546
rect 8730 6570 8748 6588
rect 8730 6588 8748 6606
rect 8730 6606 8748 6624
rect 8730 6624 8748 6642
rect 8730 6642 8748 6660
rect 8730 6660 8748 6678
rect 8730 6678 8748 6696
rect 8730 6696 8748 6714
rect 8730 6714 8748 6732
rect 8730 6732 8748 6750
rect 8730 6750 8748 6768
rect 8730 6768 8748 6786
rect 8730 6786 8748 6804
rect 8730 6804 8748 6822
rect 8730 6822 8748 6840
rect 8730 6840 8748 6858
rect 8730 6858 8748 6876
rect 8730 6876 8748 6894
rect 8730 6894 8748 6912
rect 8730 6912 8748 6930
rect 8730 6930 8748 6948
rect 8730 6948 8748 6966
rect 8730 6966 8748 6984
rect 8730 6984 8748 7002
rect 8730 7002 8748 7020
rect 8730 7020 8748 7038
rect 8730 7038 8748 7056
rect 8730 7056 8748 7074
rect 8730 7074 8748 7092
rect 8730 7092 8748 7110
rect 8730 7110 8748 7128
rect 8730 7128 8748 7146
rect 8730 7146 8748 7164
rect 8730 7164 8748 7182
rect 8730 7182 8748 7200
rect 8730 7200 8748 7218
rect 8730 7218 8748 7236
rect 8730 7236 8748 7254
rect 8730 7254 8748 7272
rect 8730 7272 8748 7290
rect 8730 7290 8748 7308
rect 8730 7308 8748 7326
rect 8730 7326 8748 7344
rect 8730 7344 8748 7362
rect 8730 7362 8748 7380
rect 8730 7380 8748 7398
rect 8730 7398 8748 7416
rect 8730 7416 8748 7434
rect 8730 7434 8748 7452
rect 8730 7452 8748 7470
rect 8730 7470 8748 7488
rect 8730 7488 8748 7506
rect 8748 3096 8766 3114
rect 8748 3114 8766 3132
rect 8748 3132 8766 3150
rect 8748 3150 8766 3168
rect 8748 3168 8766 3186
rect 8748 3186 8766 3204
rect 8748 3204 8766 3222
rect 8748 3222 8766 3240
rect 8748 3240 8766 3258
rect 8748 3258 8766 3276
rect 8748 3276 8766 3294
rect 8748 3294 8766 3312
rect 8748 3312 8766 3330
rect 8748 3330 8766 3348
rect 8748 3348 8766 3366
rect 8748 3366 8766 3384
rect 8748 3384 8766 3402
rect 8748 3402 8766 3420
rect 8748 3420 8766 3438
rect 8748 3438 8766 3456
rect 8748 3456 8766 3474
rect 8748 3474 8766 3492
rect 8748 3492 8766 3510
rect 8748 3510 8766 3528
rect 8748 3528 8766 3546
rect 8748 6660 8766 6678
rect 8748 6678 8766 6696
rect 8748 6696 8766 6714
rect 8748 6714 8766 6732
rect 8748 6732 8766 6750
rect 8748 6750 8766 6768
rect 8748 6768 8766 6786
rect 8748 6786 8766 6804
rect 8748 6804 8766 6822
rect 8748 6822 8766 6840
rect 8748 6840 8766 6858
rect 8748 6858 8766 6876
rect 8748 6876 8766 6894
rect 8748 6894 8766 6912
rect 8748 6912 8766 6930
rect 8748 6930 8766 6948
rect 8748 6948 8766 6966
rect 8748 6966 8766 6984
rect 8748 6984 8766 7002
rect 8748 7002 8766 7020
rect 8748 7020 8766 7038
rect 8748 7038 8766 7056
rect 8748 7056 8766 7074
rect 8748 7074 8766 7092
rect 8748 7092 8766 7110
rect 8748 7110 8766 7128
rect 8748 7128 8766 7146
rect 8748 7146 8766 7164
rect 8748 7164 8766 7182
rect 8748 7182 8766 7200
rect 8748 7200 8766 7218
rect 8748 7218 8766 7236
rect 8748 7236 8766 7254
rect 8748 7254 8766 7272
rect 8748 7272 8766 7290
rect 8748 7290 8766 7308
rect 8748 7308 8766 7326
rect 8748 7326 8766 7344
rect 8748 7344 8766 7362
rect 8748 7362 8766 7380
rect 8748 7380 8766 7398
rect 8748 7398 8766 7416
rect 8748 7416 8766 7434
rect 8748 7434 8766 7452
rect 8748 7452 8766 7470
rect 8748 7470 8766 7488
rect 8748 7488 8766 7506
rect 8748 7506 8766 7524
rect 8766 3132 8784 3150
rect 8766 3150 8784 3168
rect 8766 3168 8784 3186
rect 8766 3186 8784 3204
rect 8766 3204 8784 3222
rect 8766 3222 8784 3240
rect 8766 3240 8784 3258
rect 8766 3258 8784 3276
rect 8766 3276 8784 3294
rect 8766 3294 8784 3312
rect 8766 3312 8784 3330
rect 8766 3330 8784 3348
rect 8766 3348 8784 3366
rect 8766 3366 8784 3384
rect 8766 3384 8784 3402
rect 8766 3402 8784 3420
rect 8766 3420 8784 3438
rect 8766 3438 8784 3456
rect 8766 3456 8784 3474
rect 8766 3474 8784 3492
rect 8766 3492 8784 3510
rect 8766 3510 8784 3528
rect 8766 3528 8784 3546
rect 8766 6804 8784 6822
rect 8766 6822 8784 6840
rect 8766 6840 8784 6858
rect 8766 6858 8784 6876
rect 8766 6876 8784 6894
rect 8766 6894 8784 6912
rect 8766 6912 8784 6930
rect 8766 6930 8784 6948
rect 8766 6948 8784 6966
rect 8766 6966 8784 6984
rect 8766 6984 8784 7002
rect 8766 7002 8784 7020
rect 8766 7020 8784 7038
rect 8766 7038 8784 7056
rect 8766 7056 8784 7074
rect 8766 7074 8784 7092
rect 8766 7092 8784 7110
rect 8766 7110 8784 7128
rect 8766 7128 8784 7146
rect 8766 7146 8784 7164
rect 8766 7164 8784 7182
rect 8766 7182 8784 7200
rect 8766 7200 8784 7218
rect 8766 7218 8784 7236
rect 8766 7236 8784 7254
rect 8766 7254 8784 7272
rect 8766 7272 8784 7290
rect 8766 7290 8784 7308
rect 8766 7308 8784 7326
rect 8766 7326 8784 7344
rect 8766 7344 8784 7362
rect 8766 7362 8784 7380
rect 8766 7380 8784 7398
rect 8766 7398 8784 7416
rect 8766 7416 8784 7434
rect 8766 7434 8784 7452
rect 8766 7452 8784 7470
rect 8766 7470 8784 7488
rect 8766 7488 8784 7506
rect 8766 7506 8784 7524
rect 8766 7524 8784 7542
rect 8784 3150 8802 3168
rect 8784 3168 8802 3186
rect 8784 3186 8802 3204
rect 8784 3204 8802 3222
rect 8784 3222 8802 3240
rect 8784 3240 8802 3258
rect 8784 3258 8802 3276
rect 8784 3276 8802 3294
rect 8784 3294 8802 3312
rect 8784 3312 8802 3330
rect 8784 3330 8802 3348
rect 8784 3348 8802 3366
rect 8784 3366 8802 3384
rect 8784 3384 8802 3402
rect 8784 3402 8802 3420
rect 8784 3420 8802 3438
rect 8784 3438 8802 3456
rect 8784 3456 8802 3474
rect 8784 3474 8802 3492
rect 8784 3492 8802 3510
rect 8784 3510 8802 3528
rect 8784 3528 8802 3546
rect 8784 3546 8802 3564
rect 8802 3186 8820 3204
rect 8802 3204 8820 3222
rect 8802 3222 8820 3240
rect 8802 3240 8820 3258
rect 8802 3258 8820 3276
rect 8802 3276 8820 3294
rect 8802 3294 8820 3312
rect 8802 3312 8820 3330
rect 8802 3330 8820 3348
rect 8802 3348 8820 3366
rect 8802 3366 8820 3384
rect 8802 3384 8820 3402
rect 8802 3402 8820 3420
rect 8802 3420 8820 3438
rect 8802 3438 8820 3456
rect 8802 3456 8820 3474
rect 8802 3474 8820 3492
rect 8802 3492 8820 3510
rect 8802 3510 8820 3528
rect 8802 3528 8820 3546
rect 8802 3546 8820 3564
rect 8820 3222 8838 3240
rect 8820 3240 8838 3258
rect 8820 3258 8838 3276
rect 8820 3276 8838 3294
rect 8820 3294 8838 3312
rect 8820 3312 8838 3330
rect 8820 3330 8838 3348
rect 8820 3348 8838 3366
rect 8820 3366 8838 3384
rect 8820 3384 8838 3402
rect 8820 3402 8838 3420
rect 8820 3420 8838 3438
rect 8820 3438 8838 3456
rect 8820 3456 8838 3474
rect 8820 3474 8838 3492
rect 8820 3492 8838 3510
rect 8820 3510 8838 3528
rect 8820 3528 8838 3546
rect 8820 3546 8838 3564
rect 8838 3258 8856 3276
rect 8838 3276 8856 3294
rect 8838 3294 8856 3312
rect 8838 3312 8856 3330
rect 8838 3330 8856 3348
rect 8838 3348 8856 3366
rect 8838 3366 8856 3384
rect 8838 3384 8856 3402
rect 8838 3402 8856 3420
rect 8838 3420 8856 3438
rect 8838 3438 8856 3456
rect 8838 3456 8856 3474
rect 8838 3474 8856 3492
rect 8838 3492 8856 3510
rect 8838 3510 8856 3528
rect 8838 3528 8856 3546
rect 8838 3546 8856 3564
rect 8856 3294 8874 3312
rect 8856 3312 8874 3330
rect 8856 3330 8874 3348
rect 8856 3348 8874 3366
rect 8856 3366 8874 3384
rect 8856 3384 8874 3402
rect 8856 3402 8874 3420
rect 8856 3420 8874 3438
rect 8856 3438 8874 3456
rect 8856 3456 8874 3474
rect 8856 3474 8874 3492
rect 8856 3492 8874 3510
rect 8856 3510 8874 3528
rect 8856 3528 8874 3546
rect 8856 3546 8874 3564
rect 8856 3564 8874 3582
rect 8874 3330 8892 3348
rect 8874 3348 8892 3366
rect 8874 3366 8892 3384
rect 8874 3384 8892 3402
rect 8874 3402 8892 3420
rect 8874 3420 8892 3438
rect 8874 3438 8892 3456
rect 8874 3456 8892 3474
rect 8874 3474 8892 3492
rect 8874 3492 8892 3510
rect 8874 3510 8892 3528
rect 8874 3528 8892 3546
rect 8874 3546 8892 3564
rect 8874 3564 8892 3582
rect 8892 3366 8910 3384
rect 8892 3384 8910 3402
rect 8892 3402 8910 3420
rect 8892 3420 8910 3438
rect 8892 3438 8910 3456
rect 8892 3456 8910 3474
rect 8892 3474 8910 3492
rect 8892 3492 8910 3510
rect 8892 3510 8910 3528
rect 8892 3528 8910 3546
rect 8892 3546 8910 3564
rect 8892 3564 8910 3582
rect 8910 3402 8928 3420
rect 8910 3420 8928 3438
rect 8910 3438 8928 3456
rect 8910 3456 8928 3474
rect 8910 3474 8928 3492
rect 8910 3492 8928 3510
rect 8910 3510 8928 3528
rect 8910 3528 8928 3546
rect 8910 3546 8928 3564
rect 8910 3564 8928 3582
rect 8928 3456 8946 3474
rect 8928 3474 8946 3492
rect 8928 3492 8946 3510
rect 8928 3510 8946 3528
rect 8928 3528 8946 3546
rect 8928 3546 8946 3564
rect 8928 3564 8946 3582
rect 8928 3582 8946 3600
rect 8946 3492 8964 3510
rect 8946 3510 8964 3528
rect 8946 3528 8964 3546
rect 8946 3546 8964 3564
rect 8946 3564 8964 3582
rect 8946 3582 8964 3600
rect 8964 3546 8982 3564
rect 8964 3564 8982 3582
rect 8964 3582 8982 3600
rect 8982 3582 9000 3600
<< properties >>
string FIXED_BBOX 0 0 9000 10566
<< end >>
