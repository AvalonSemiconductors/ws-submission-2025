VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin
  CLASS BLOCK ;
  FOREIGN tholin ;
  ORIGIN 0.000 0.000 ;
  SIZE 702.000 BY 583.200 ;
  OBS
      LAYER Metal1 ;
        RECT 6.000 4.800 695.400 577.800 ;
      LAYER Metal2 ;
        RECT 6.000 4.800 695.400 577.800 ;
      LAYER Metal3 ;
        RECT 6.000 4.800 695.400 577.800 ;
      LAYER Metal4 ;
        RECT 103.800 577.200 105.000 577.800 ;
        RECT 103.200 576.600 106.200 577.200 ;
        RECT 103.200 576.000 106.800 576.600 ;
        RECT 103.800 575.400 107.400 576.000 ;
        RECT 103.800 574.800 108.000 575.400 ;
        RECT 104.400 574.200 109.200 574.800 ;
        RECT 104.400 573.600 109.800 574.200 ;
        RECT 104.400 573.000 110.400 573.600 ;
        RECT 104.400 572.400 111.000 573.000 ;
        RECT 104.400 571.800 112.200 572.400 ;
        RECT 105.000 571.200 112.800 571.800 ;
        RECT 105.000 568.800 108.000 571.200 ;
        RECT 109.200 570.600 113.400 571.200 ;
        RECT 109.800 570.000 114.000 570.600 ;
        RECT 110.400 569.400 115.200 570.000 ;
        RECT 111.000 568.800 115.800 569.400 ;
        RECT 105.600 565.800 108.600 568.800 ;
        RECT 112.200 568.200 116.400 568.800 ;
        RECT 112.800 567.600 117.000 568.200 ;
        RECT 113.400 567.000 117.600 567.600 ;
        RECT 114.000 566.400 118.200 567.000 ;
        RECT 114.600 565.800 119.400 566.400 ;
        RECT 106.200 562.800 109.200 565.800 ;
        RECT 115.200 565.200 120.000 565.800 ;
        RECT 116.400 564.600 120.600 565.200 ;
        RECT 117.000 564.000 121.200 564.600 ;
        RECT 117.600 563.400 121.800 564.000 ;
        RECT 118.200 562.800 122.400 563.400 ;
        RECT 106.800 562.200 109.200 562.800 ;
        RECT 118.800 562.200 123.000 562.800 ;
        RECT 106.800 558.000 109.800 562.200 ;
        RECT 119.400 561.600 123.600 562.200 ;
        RECT 120.000 561.000 124.200 561.600 ;
        RECT 120.600 560.400 125.400 561.000 ;
        RECT 121.200 559.800 126.000 560.400 ;
        RECT 122.400 559.200 126.600 559.800 ;
        RECT 123.000 558.600 127.200 559.200 ;
        RECT 123.600 558.000 127.800 558.600 ;
        RECT 107.400 557.400 109.800 558.000 ;
        RECT 124.200 557.400 128.400 558.000 ;
        RECT 107.400 550.200 110.400 557.400 ;
        RECT 124.800 556.800 129.000 557.400 ;
        RECT 125.400 556.200 129.600 556.800 ;
        RECT 126.000 555.600 130.200 556.200 ;
        RECT 126.600 555.000 130.800 555.600 ;
        RECT 127.200 554.400 131.400 555.000 ;
        RECT 127.800 553.800 132.000 554.400 ;
        RECT 128.400 553.200 132.600 553.800 ;
        RECT 129.000 552.600 133.200 553.200 ;
        RECT 129.600 552.000 133.800 552.600 ;
        RECT 130.200 551.400 134.400 552.000 ;
        RECT 130.800 550.800 135.000 551.400 ;
        RECT 131.400 550.200 135.000 550.800 ;
        RECT 108.000 549.000 110.400 550.200 ;
        RECT 132.000 549.600 135.600 550.200 ;
        RECT 132.600 549.000 136.200 549.600 ;
        RECT 7.200 546.000 9.000 546.600 ;
        RECT 6.000 545.400 9.600 546.000 ;
        RECT 6.600 544.800 10.800 545.400 ;
        RECT 6.600 544.200 12.000 544.800 ;
        RECT 7.200 543.600 13.200 544.200 ;
        RECT 7.200 543.000 13.800 543.600 ;
        RECT 7.200 542.400 15.000 543.000 ;
        RECT 7.800 541.800 16.200 542.400 ;
        RECT 7.800 541.200 17.400 541.800 ;
        RECT 8.400 540.600 18.600 541.200 ;
        RECT 8.400 540.000 19.800 540.600 ;
        RECT 9.000 538.800 12.600 540.000 ;
        RECT 14.400 539.400 20.400 540.000 ;
        RECT 15.600 538.800 21.600 539.400 ;
        RECT 9.600 538.200 13.200 538.800 ;
        RECT 16.200 538.200 22.800 538.800 ;
        RECT 10.200 537.000 13.800 538.200 ;
        RECT 17.400 537.600 23.400 538.200 ;
        RECT 18.600 537.000 24.600 537.600 ;
        RECT 10.800 536.400 14.400 537.000 ;
        RECT 19.800 536.400 25.800 537.000 ;
        RECT 10.800 535.800 15.000 536.400 ;
        RECT 21.000 535.800 26.400 536.400 ;
        RECT 11.400 535.200 15.000 535.800 ;
        RECT 21.600 535.200 27.600 535.800 ;
        RECT 12.000 534.000 15.600 535.200 ;
        RECT 22.800 534.600 28.800 535.200 ;
        RECT 24.000 534.000 30.000 534.600 ;
        RECT 108.000 534.000 111.000 549.000 ;
        RECT 133.200 548.400 136.800 549.000 ;
        RECT 133.800 547.800 137.400 548.400 ;
        RECT 133.800 547.200 138.000 547.800 ;
        RECT 134.400 546.600 138.600 547.200 ;
        RECT 135.000 546.000 139.200 546.600 ;
        RECT 135.600 545.400 139.800 546.000 ;
        RECT 136.200 544.800 140.400 545.400 ;
        RECT 136.800 544.200 140.400 544.800 ;
        RECT 137.400 543.600 141.000 544.200 ;
        RECT 138.000 543.000 141.600 543.600 ;
        RECT 138.600 542.400 142.200 543.000 ;
        RECT 138.600 541.800 142.800 542.400 ;
        RECT 139.200 541.200 143.400 541.800 ;
        RECT 139.800 540.600 144.000 541.200 ;
        RECT 140.400 540.000 144.600 540.600 ;
        RECT 141.000 539.400 144.600 540.000 ;
        RECT 141.600 538.800 145.200 539.400 ;
        RECT 142.200 538.200 145.800 538.800 ;
        RECT 142.800 537.600 146.400 538.200 ;
        RECT 142.800 537.000 147.000 537.600 ;
        RECT 143.400 536.400 147.600 537.000 ;
        RECT 144.000 535.800 147.600 536.400 ;
        RECT 144.600 535.200 148.200 535.800 ;
        RECT 145.200 534.600 148.800 535.200 ;
        RECT 12.600 533.400 16.200 534.000 ;
        RECT 24.600 533.400 30.600 534.000 ;
        RECT 13.200 532.200 16.800 533.400 ;
        RECT 25.800 532.800 31.800 533.400 ;
        RECT 27.000 532.200 33.000 532.800 ;
        RECT 108.600 532.200 111.000 534.000 ;
        RECT 145.800 534.000 149.400 534.600 ;
        RECT 145.800 533.400 150.000 534.000 ;
        RECT 146.400 532.800 150.000 533.400 ;
        RECT 147.000 532.200 150.600 532.800 ;
        RECT 13.800 531.600 17.400 532.200 ;
        RECT 27.600 531.600 33.600 532.200 ;
        RECT 14.400 531.000 17.400 531.600 ;
        RECT 28.800 531.000 34.800 531.600 ;
        RECT 14.400 530.400 18.000 531.000 ;
        RECT 29.400 530.400 36.000 531.000 ;
        RECT 15.000 529.200 18.600 530.400 ;
        RECT 30.600 529.800 36.600 530.400 ;
        RECT 31.800 529.200 37.800 529.800 ;
        RECT 15.600 528.600 19.200 529.200 ;
        RECT 33.000 528.600 39.000 529.200 ;
        RECT 16.200 528.000 19.200 528.600 ;
        RECT 34.200 528.000 39.600 528.600 ;
        RECT 16.200 527.400 19.800 528.000 ;
        RECT 35.400 527.400 40.800 528.000 ;
        RECT 16.800 526.200 20.400 527.400 ;
        RECT 36.000 526.800 42.000 527.400 ;
        RECT 37.200 526.200 42.600 526.800 ;
        RECT 17.400 525.600 21.000 526.200 ;
        RECT 38.400 525.600 43.800 526.200 ;
        RECT 18.000 525.000 21.000 525.600 ;
        RECT 39.000 525.000 44.400 525.600 ;
        RECT 18.000 524.400 21.600 525.000 ;
        RECT 40.200 524.400 45.600 525.000 ;
        RECT 18.600 523.800 21.600 524.400 ;
        RECT 40.800 523.800 46.800 524.400 ;
        RECT 18.600 523.200 22.200 523.800 ;
        RECT 42.000 523.200 47.400 523.800 ;
        RECT 19.200 522.600 22.800 523.200 ;
        RECT 43.200 522.600 48.600 523.200 ;
        RECT 108.600 522.600 111.600 532.200 ;
        RECT 147.600 531.600 151.200 532.200 ;
        RECT 148.200 531.000 151.800 531.600 ;
        RECT 148.200 530.400 152.400 531.000 ;
        RECT 148.800 529.800 152.400 530.400 ;
        RECT 149.400 529.200 153.000 529.800 ;
        RECT 150.000 528.600 153.600 529.200 ;
        RECT 150.600 528.000 154.200 528.600 ;
        RECT 150.600 527.400 154.800 528.000 ;
        RECT 151.200 526.800 154.800 527.400 ;
        RECT 151.800 526.200 155.400 526.800 ;
        RECT 152.400 525.600 156.000 526.200 ;
        RECT 153.000 524.400 156.600 525.600 ;
        RECT 153.600 523.800 157.200 524.400 ;
        RECT 154.200 523.200 157.800 523.800 ;
        RECT 19.800 522.000 22.800 522.600 ;
        RECT 43.800 522.000 49.800 522.600 ;
        RECT 109.200 522.000 111.600 522.600 ;
        RECT 154.800 522.000 158.400 523.200 ;
        RECT 19.800 521.400 23.400 522.000 ;
        RECT 45.000 521.400 50.400 522.000 ;
        RECT 20.400 520.800 23.400 521.400 ;
        RECT 46.200 520.800 51.600 521.400 ;
        RECT 20.400 520.200 24.000 520.800 ;
        RECT 46.800 520.200 52.200 520.800 ;
        RECT 21.000 519.600 24.000 520.200 ;
        RECT 48.000 519.600 53.400 520.200 ;
        RECT 21.000 519.000 24.600 519.600 ;
        RECT 48.600 519.000 54.000 519.600 ;
        RECT 21.600 518.400 24.600 519.000 ;
        RECT 49.800 518.400 55.200 519.000 ;
        RECT 21.600 517.800 25.200 518.400 ;
        RECT 51.000 517.800 56.400 518.400 ;
        RECT 22.200 517.200 25.200 517.800 ;
        RECT 51.600 517.200 57.000 517.800 ;
        RECT 22.200 516.600 25.800 517.200 ;
        RECT 52.800 516.600 58.200 517.200 ;
        RECT 22.800 516.000 25.800 516.600 ;
        RECT 53.400 516.000 58.800 516.600 ;
        RECT 109.200 516.000 112.200 522.000 ;
        RECT 155.400 521.400 159.000 522.000 ;
        RECT 156.000 520.800 159.600 521.400 ;
        RECT 156.600 519.600 160.200 520.800 ;
        RECT 157.200 519.000 160.800 519.600 ;
        RECT 157.800 518.400 161.400 519.000 ;
        RECT 158.400 517.200 162.000 518.400 ;
        RECT 159.000 516.600 162.600 517.200 ;
        RECT 159.600 516.000 163.200 516.600 ;
        RECT 22.800 515.400 26.400 516.000 ;
        RECT 54.600 515.400 60.000 516.000 ;
        RECT 109.800 515.400 112.200 516.000 ;
        RECT 23.400 514.200 26.400 515.400 ;
        RECT 55.200 514.800 60.600 515.400 ;
        RECT 56.400 514.200 61.800 514.800 ;
        RECT 24.000 513.000 27.000 514.200 ;
        RECT 57.600 513.600 63.000 514.200 ;
        RECT 58.200 513.000 63.600 513.600 ;
        RECT 24.000 512.400 27.600 513.000 ;
        RECT 59.400 512.400 64.800 513.000 ;
        RECT 24.600 511.800 27.600 512.400 ;
        RECT 60.000 511.800 65.400 512.400 ;
        RECT 24.600 511.200 28.200 511.800 ;
        RECT 61.200 511.200 66.600 511.800 ;
        RECT 25.200 510.600 28.200 511.200 ;
        RECT 61.800 510.600 67.200 511.200 ;
        RECT 109.800 510.600 112.800 515.400 ;
        RECT 160.200 514.800 163.800 516.000 ;
        RECT 160.800 514.200 164.400 514.800 ;
        RECT 161.400 513.600 165.000 514.200 ;
        RECT 162.000 512.400 165.600 513.600 ;
        RECT 162.600 511.800 166.200 512.400 ;
        RECT 163.200 510.600 166.800 511.800 ;
        RECT 25.200 510.000 28.800 510.600 ;
        RECT 63.000 510.000 68.400 510.600 ;
        RECT 25.800 508.800 28.800 510.000 ;
        RECT 63.600 509.400 69.000 510.000 ;
        RECT 64.800 508.800 70.200 509.400 ;
        RECT 26.400 507.600 29.400 508.800 ;
        RECT 65.400 508.200 70.800 508.800 ;
        RECT 66.600 507.600 72.000 508.200 ;
        RECT 26.400 507.000 30.000 507.600 ;
        RECT 67.200 507.000 72.600 507.600 ;
        RECT 110.400 507.000 113.400 510.600 ;
        RECT 163.800 510.000 167.400 510.600 ;
        RECT 164.400 509.400 168.000 510.000 ;
        RECT 164.400 508.800 168.600 509.400 ;
        RECT 165.000 508.200 168.600 508.800 ;
        RECT 165.600 507.600 169.200 508.200 ;
        RECT 165.600 507.000 169.800 507.600 ;
        RECT 27.000 506.400 30.000 507.000 ;
        RECT 68.400 506.400 73.800 507.000 ;
        RECT 27.000 505.800 30.600 506.400 ;
        RECT 69.000 505.800 74.400 506.400 ;
        RECT 27.600 505.200 30.600 505.800 ;
        RECT 70.200 505.200 75.600 505.800 ;
        RECT 27.600 504.600 31.200 505.200 ;
        RECT 70.800 504.600 76.200 505.200 ;
        RECT 111.000 504.600 114.000 507.000 ;
        RECT 166.200 506.400 170.400 507.000 ;
        RECT 166.800 505.800 170.400 506.400 ;
        RECT 167.400 505.200 171.000 505.800 ;
        RECT 168.000 504.600 171.600 505.200 ;
        RECT 28.200 503.400 31.200 504.600 ;
        RECT 72.000 504.000 77.400 504.600 ;
        RECT 72.600 503.400 78.000 504.000 ;
        RECT 28.800 502.200 31.800 503.400 ;
        RECT 73.800 502.800 79.200 503.400 ;
        RECT 75.000 502.200 79.800 502.800 ;
        RECT 28.800 501.600 32.400 502.200 ;
        RECT 75.600 501.600 81.000 502.200 ;
        RECT 111.600 501.600 114.600 504.600 ;
        RECT 168.000 504.000 172.200 504.600 ;
        RECT 168.600 503.400 172.200 504.000 ;
        RECT 169.200 502.800 172.800 503.400 ;
        RECT 169.800 502.200 173.400 502.800 ;
        RECT 169.800 501.600 174.000 502.200 ;
        RECT 29.400 501.000 32.400 501.600 ;
        RECT 76.800 501.000 81.600 501.600 ;
        RECT 29.400 500.400 33.000 501.000 ;
        RECT 77.400 500.400 82.800 501.000 ;
        RECT 30.000 499.800 33.000 500.400 ;
        RECT 78.600 499.800 83.400 500.400 ;
        RECT 30.000 499.200 33.600 499.800 ;
        RECT 79.200 499.200 84.600 499.800 ;
        RECT 112.200 499.200 115.200 501.600 ;
        RECT 170.400 501.000 174.000 501.600 ;
        RECT 171.000 500.400 174.600 501.000 ;
        RECT 178.800 500.400 180.600 501.000 ;
        RECT 171.600 499.200 175.200 500.400 ;
        RECT 177.000 499.800 181.800 500.400 ;
        RECT 176.400 499.200 183.000 499.800 ;
        RECT 30.600 498.000 33.600 499.200 ;
        RECT 80.400 498.600 85.200 499.200 ;
        RECT 81.000 498.000 86.400 498.600 ;
        RECT 31.200 496.800 34.200 498.000 ;
        RECT 82.200 497.400 87.000 498.000 ;
        RECT 112.800 497.400 115.800 499.200 ;
        RECT 172.200 498.600 184.200 499.200 ;
        RECT 172.800 498.000 184.800 498.600 ;
        RECT 82.800 496.800 88.200 497.400 ;
        RECT 113.400 496.800 115.800 497.400 ;
        RECT 173.400 497.400 178.800 498.000 ;
        RECT 180.000 497.400 185.400 498.000 ;
        RECT 173.400 496.800 178.200 497.400 ;
        RECT 181.200 496.800 186.000 497.400 ;
        RECT 31.200 496.200 34.800 496.800 ;
        RECT 84.000 496.200 88.800 496.800 ;
        RECT 31.800 495.600 34.800 496.200 ;
        RECT 84.600 495.600 90.000 496.200 ;
        RECT 113.400 495.600 116.400 496.800 ;
        RECT 174.000 496.200 178.200 496.800 ;
        RECT 182.400 496.200 186.600 496.800 ;
        RECT 174.600 495.600 178.200 496.200 ;
        RECT 183.000 495.600 187.200 496.200 ;
        RECT 31.800 495.000 35.400 495.600 ;
        RECT 85.800 495.000 90.600 495.600 ;
        RECT 114.000 495.000 116.400 495.600 ;
        RECT 32.400 494.400 35.400 495.000 ;
        RECT 86.400 494.400 91.800 495.000 ;
        RECT 32.400 493.800 36.000 494.400 ;
        RECT 87.600 493.800 92.400 494.400 ;
        RECT 114.000 493.800 117.000 495.000 ;
        RECT 33.000 492.600 36.000 493.800 ;
        RECT 88.200 493.200 93.600 493.800 ;
        RECT 114.600 493.200 117.000 493.800 ;
        RECT 89.400 492.600 94.200 493.200 ;
        RECT 33.600 491.400 36.600 492.600 ;
        RECT 90.000 492.000 95.400 492.600 ;
        RECT 114.600 492.000 117.600 493.200 ;
        RECT 91.200 491.400 96.000 492.000 ;
        RECT 33.600 490.800 37.200 491.400 ;
        RECT 91.800 490.800 97.200 491.400 ;
        RECT 115.200 490.800 117.600 492.000 ;
        RECT 155.400 491.400 157.800 492.000 ;
        RECT 154.200 490.800 158.400 491.400 ;
        RECT 175.200 490.800 178.200 495.600 ;
        RECT 183.600 495.000 187.200 495.600 ;
        RECT 184.200 494.400 187.800 495.000 ;
        RECT 184.800 493.800 187.800 494.400 ;
        RECT 184.800 493.200 188.400 493.800 ;
        RECT 185.400 492.600 188.400 493.200 ;
        RECT 185.400 492.000 189.000 492.600 ;
        RECT 186.000 490.800 189.000 492.000 ;
        RECT 34.200 490.200 37.200 490.800 ;
        RECT 93.000 490.200 97.800 490.800 ;
        RECT 113.400 490.200 118.200 490.800 ;
        RECT 153.600 490.200 159.000 490.800 ;
        RECT 34.200 489.600 37.800 490.200 ;
        RECT 93.600 489.600 99.000 490.200 ;
        RECT 111.000 489.600 121.800 490.200 ;
        RECT 132.000 489.600 138.600 490.200 ;
        RECT 153.600 489.600 159.600 490.200 ;
        RECT 34.800 489.000 37.800 489.600 ;
        RECT 94.800 489.000 100.200 489.600 ;
        RECT 109.800 489.000 123.600 489.600 ;
        RECT 131.400 489.000 140.400 489.600 ;
        RECT 34.800 488.400 38.400 489.000 ;
        RECT 95.400 488.400 100.800 489.000 ;
        RECT 109.200 488.400 125.400 489.000 ;
        RECT 130.800 488.400 142.800 489.000 ;
        RECT 153.000 488.400 160.200 489.600 ;
        RECT 175.800 489.000 178.800 490.800 ;
        RECT 175.800 488.400 179.400 489.000 ;
        RECT 35.400 487.800 38.400 488.400 ;
        RECT 96.600 487.800 102.000 488.400 ;
        RECT 108.600 487.800 127.200 488.400 ;
        RECT 130.800 487.800 144.600 488.400 ;
        RECT 152.400 487.800 156.000 488.400 ;
        RECT 157.200 487.800 160.800 488.400 ;
        RECT 35.400 487.200 39.000 487.800 ;
        RECT 97.200 487.200 102.600 487.800 ;
        RECT 108.600 487.200 113.400 487.800 ;
        RECT 120.000 487.200 128.400 487.800 ;
        RECT 130.800 487.200 145.800 487.800 ;
        RECT 36.000 486.000 39.000 487.200 ;
        RECT 98.400 486.600 103.800 487.200 ;
        RECT 99.000 486.000 104.400 486.600 ;
        RECT 108.600 486.000 111.600 487.200 ;
        RECT 121.800 486.600 129.600 487.200 ;
        RECT 130.800 486.600 134.400 487.200 ;
        RECT 138.600 486.600 147.600 487.200 ;
        RECT 152.400 486.600 155.400 487.800 ;
        RECT 157.800 487.200 160.800 487.800 ;
        RECT 176.400 487.200 179.400 488.400 ;
        RECT 157.800 486.600 161.400 487.200 ;
        RECT 123.600 486.000 134.400 486.600 ;
        RECT 140.400 486.000 148.800 486.600 ;
        RECT 151.800 486.000 155.400 486.600 ;
        RECT 36.600 484.800 39.600 486.000 ;
        RECT 100.200 485.400 105.600 486.000 ;
        RECT 108.600 485.400 112.200 486.000 ;
        RECT 125.400 485.400 135.000 486.000 ;
        RECT 142.200 485.400 150.600 486.000 ;
        RECT 151.800 485.400 154.800 486.000 ;
        RECT 158.400 485.400 161.400 486.600 ;
        RECT 177.000 486.000 180.000 487.200 ;
        RECT 186.600 486.000 189.600 490.800 ;
        RECT 194.400 489.000 198.600 489.600 ;
        RECT 193.200 488.400 199.800 489.000 ;
        RECT 192.600 487.800 200.400 488.400 ;
        RECT 192.000 487.200 201.000 487.800 ;
        RECT 191.400 486.600 201.000 487.200 ;
        RECT 190.800 486.000 195.000 486.600 ;
        RECT 198.000 486.000 201.600 486.600 ;
        RECT 177.000 485.400 180.600 486.000 ;
        RECT 100.800 484.800 106.800 485.400 ;
        RECT 109.200 484.800 113.400 485.400 ;
        RECT 126.600 484.800 135.600 485.400 ;
        RECT 144.000 484.800 154.800 485.400 ;
        RECT 37.200 483.600 40.200 484.800 ;
        RECT 102.000 484.200 107.400 484.800 ;
        RECT 109.200 484.200 114.600 484.800 ;
        RECT 127.800 484.200 136.200 484.800 ;
        RECT 145.800 484.200 154.800 484.800 ;
        RECT 103.200 483.600 115.200 484.200 ;
        RECT 129.000 483.600 136.800 484.200 ;
        RECT 147.000 483.600 154.800 484.200 ;
        RECT 159.000 484.200 162.000 485.400 ;
        RECT 169.800 484.800 173.400 485.400 ;
        RECT 177.600 484.800 180.600 485.400 ;
        RECT 186.600 485.400 194.400 486.000 ;
        RECT 186.600 484.800 193.800 485.400 ;
        RECT 198.600 484.800 201.600 486.000 ;
        RECT 168.600 484.200 175.200 484.800 ;
        RECT 177.600 484.200 181.200 484.800 ;
        RECT 186.600 484.200 193.200 484.800 ;
        RECT 198.600 484.200 208.200 484.800 ;
        RECT 159.000 483.600 162.600 484.200 ;
        RECT 168.000 483.600 176.400 484.200 ;
        RECT 37.200 483.000 40.800 483.600 ;
        RECT 103.800 483.000 117.000 483.600 ;
        RECT 130.200 483.000 137.400 483.600 ;
        RECT 148.800 483.000 154.800 483.600 ;
        RECT 37.800 482.400 40.800 483.000 ;
        RECT 105.000 482.400 118.200 483.000 ;
        RECT 131.400 482.400 138.000 483.000 ;
        RECT 150.000 482.400 154.800 483.000 ;
        RECT 159.600 482.400 162.600 483.600 ;
        RECT 167.400 483.000 177.000 483.600 ;
        RECT 178.200 483.000 181.800 484.200 ;
        RECT 186.600 483.600 192.600 484.200 ;
        RECT 198.000 483.600 209.400 484.200 ;
        RECT 166.800 482.400 182.400 483.000 ;
        RECT 37.800 481.800 41.400 482.400 ;
        RECT 105.600 481.800 120.000 482.400 ;
        RECT 134.400 481.800 139.200 482.400 ;
        RECT 38.400 481.200 41.400 481.800 ;
        RECT 106.800 481.200 122.400 481.800 ;
        RECT 135.000 481.200 139.800 481.800 ;
        RECT 38.400 480.600 42.000 481.200 ;
        RECT 106.800 480.600 124.800 481.200 ;
        RECT 135.600 480.600 141.000 481.200 ;
        RECT 39.000 480.000 42.000 480.600 ;
        RECT 105.000 480.000 127.800 480.600 ;
        RECT 136.800 480.000 141.600 480.600 ;
        RECT 151.800 480.000 154.200 482.400 ;
        RECT 159.600 481.800 163.200 482.400 ;
        RECT 160.200 480.600 163.200 481.800 ;
        RECT 166.800 481.800 170.400 482.400 ;
        RECT 173.400 481.800 182.400 482.400 ;
        RECT 186.600 482.400 192.000 483.600 ;
        RECT 196.200 483.000 210.000 483.600 ;
        RECT 195.000 482.400 210.000 483.000 ;
        RECT 166.800 480.600 169.800 481.800 ;
        RECT 174.600 481.200 183.000 481.800 ;
        RECT 186.600 481.200 191.400 482.400 ;
        RECT 193.800 481.800 210.000 482.400 ;
        RECT 192.600 481.200 201.000 481.800 ;
        RECT 175.800 480.600 183.600 481.200 ;
        RECT 186.600 480.600 201.000 481.200 ;
        RECT 205.200 480.600 210.000 481.800 ;
        RECT 39.000 479.400 42.600 480.000 ;
        RECT 103.800 479.400 114.600 480.000 ;
        RECT 117.600 479.400 130.200 480.000 ;
        RECT 137.400 479.400 142.800 480.000 ;
        RECT 39.600 478.800 42.600 479.400 ;
        RECT 102.600 478.800 111.000 479.400 ;
        RECT 120.000 478.800 132.600 479.400 ;
        RECT 138.000 478.800 144.000 479.400 ;
        RECT 39.600 478.200 43.200 478.800 ;
        RECT 102.000 478.200 108.600 478.800 ;
        RECT 122.400 478.200 133.800 478.800 ;
        RECT 139.200 478.200 145.200 478.800 ;
        RECT 40.200 477.600 43.200 478.200 ;
        RECT 100.800 477.600 106.800 478.200 ;
        RECT 124.800 477.600 133.200 478.200 ;
        RECT 140.400 477.600 146.400 478.200 ;
        RECT 40.200 477.000 43.800 477.600 ;
        RECT 100.200 477.000 105.600 477.600 ;
        RECT 141.000 477.000 147.600 477.600 ;
        RECT 40.800 476.400 43.800 477.000 ;
        RECT 99.000 476.400 104.400 477.000 ;
        RECT 142.200 476.400 148.800 477.000 ;
        RECT 40.800 475.800 44.400 476.400 ;
        RECT 98.400 475.800 103.200 476.400 ;
        RECT 144.000 475.800 150.000 476.400 ;
        RECT 151.800 475.800 154.800 480.000 ;
        RECT 160.800 479.400 163.800 480.600 ;
        RECT 160.800 478.800 164.400 479.400 ;
        RECT 161.400 478.200 164.400 478.800 ;
        RECT 166.200 478.200 169.200 480.600 ;
        RECT 176.400 480.000 184.200 480.600 ;
        RECT 177.600 479.400 184.200 480.000 ;
        RECT 186.600 479.400 200.400 480.600 ;
        RECT 205.200 480.000 209.400 480.600 ;
        RECT 205.800 479.400 208.800 480.000 ;
        RECT 178.200 478.800 184.800 479.400 ;
        RECT 186.600 478.800 194.400 479.400 ;
        RECT 178.800 478.200 185.400 478.800 ;
        RECT 161.400 477.600 165.000 478.200 ;
        RECT 162.000 476.400 165.000 477.600 ;
        RECT 166.800 476.400 169.800 478.200 ;
        RECT 180.000 477.600 185.400 478.200 ;
        RECT 186.600 478.200 193.200 478.800 ;
        RECT 196.200 478.200 199.800 479.400 ;
        RECT 186.600 477.600 192.600 478.200 ;
        RECT 195.600 477.600 199.200 478.200 ;
        RECT 180.600 477.000 192.000 477.600 ;
        RECT 195.000 477.000 198.600 477.600 ;
        RECT 181.200 476.400 191.400 477.000 ;
        RECT 193.800 476.400 198.000 477.000 ;
        RECT 162.000 475.800 165.600 476.400 ;
        RECT 166.800 475.800 170.400 476.400 ;
        RECT 182.400 475.800 190.800 476.400 ;
        RECT 193.200 475.800 197.400 476.400 ;
        RECT 41.400 475.200 44.400 475.800 ;
        RECT 97.800 475.200 102.600 475.800 ;
        RECT 145.200 475.200 155.400 475.800 ;
        RECT 41.400 474.600 45.000 475.200 ;
        RECT 97.200 474.600 102.000 475.200 ;
        RECT 147.600 474.600 155.400 475.200 ;
        RECT 162.600 475.200 165.600 475.800 ;
        RECT 167.400 475.200 170.400 475.800 ;
        RECT 183.000 475.200 190.800 475.800 ;
        RECT 192.000 475.200 197.400 475.800 ;
        RECT 199.200 475.200 205.800 475.800 ;
        RECT 162.600 474.600 166.200 475.200 ;
        RECT 167.400 474.600 171.000 475.200 ;
        RECT 183.600 474.600 207.000 475.200 ;
        RECT 42.000 474.000 45.000 474.600 ;
        RECT 96.600 474.000 100.800 474.600 ;
        RECT 127.800 474.000 130.200 474.600 ;
        RECT 42.000 473.400 45.600 474.000 ;
        RECT 96.000 473.400 100.200 474.000 ;
        RECT 126.600 473.400 130.200 474.000 ;
        RECT 152.400 474.000 155.400 474.600 ;
        RECT 163.200 474.000 166.200 474.600 ;
        RECT 168.000 474.000 171.600 474.600 ;
        RECT 183.600 474.000 208.200 474.600 ;
        RECT 152.400 473.400 156.000 474.000 ;
        RECT 163.200 473.400 166.800 474.000 ;
        RECT 168.000 473.400 172.800 474.000 ;
        RECT 181.200 473.400 208.800 474.000 ;
        RECT 42.600 472.800 45.600 473.400 ;
        RECT 95.400 472.800 99.600 473.400 ;
        RECT 126.000 472.800 129.600 473.400 ;
        RECT 42.600 472.200 46.200 472.800 ;
        RECT 94.800 472.200 99.000 472.800 ;
        RECT 125.400 472.200 129.000 472.800 ;
        RECT 153.000 472.200 156.000 473.400 ;
        RECT 163.800 472.800 166.800 473.400 ;
        RECT 168.600 472.800 208.800 473.400 ;
        RECT 163.800 472.200 167.400 472.800 ;
        RECT 169.200 472.200 199.200 472.800 ;
        RECT 205.800 472.200 208.800 472.800 ;
        RECT 43.200 471.600 46.800 472.200 ;
        RECT 94.200 471.600 98.400 472.200 ;
        RECT 124.800 471.600 128.400 472.200 ;
        RECT 43.800 471.000 46.800 471.600 ;
        RECT 93.600 471.000 97.800 471.600 ;
        RECT 124.200 471.000 127.800 471.600 ;
        RECT 153.600 471.000 156.600 472.200 ;
        RECT 164.400 471.600 167.400 472.200 ;
        RECT 169.800 471.600 195.000 472.200 ;
        RECT 205.800 471.600 209.400 472.200 ;
        RECT 164.400 471.000 168.000 471.600 ;
        RECT 171.000 471.000 185.400 471.600 ;
        RECT 43.800 470.400 47.400 471.000 ;
        RECT 93.600 470.400 97.200 471.000 ;
        RECT 123.600 470.400 127.200 471.000 ;
        RECT 44.400 469.800 47.400 470.400 ;
        RECT 93.000 469.800 96.600 470.400 ;
        RECT 123.000 469.800 127.200 470.400 ;
        RECT 154.200 469.800 157.200 471.000 ;
        RECT 165.000 470.400 168.000 471.000 ;
        RECT 172.800 470.400 184.800 471.000 ;
        RECT 165.000 469.800 168.600 470.400 ;
        RECT 44.400 469.200 48.000 469.800 ;
        RECT 45.000 468.600 48.000 469.200 ;
        RECT 92.400 469.200 96.000 469.800 ;
        RECT 121.800 469.200 126.600 469.800 ;
        RECT 154.800 469.200 157.800 469.800 ;
        RECT 165.600 469.200 168.600 469.800 ;
        RECT 180.600 469.800 184.800 470.400 ;
        RECT 187.800 470.400 192.600 471.600 ;
        RECT 187.800 469.800 193.200 470.400 ;
        RECT 205.800 469.800 208.800 471.600 ;
        RECT 180.600 469.200 184.200 469.800 ;
        RECT 187.800 469.200 193.800 469.800 ;
        RECT 205.200 469.200 208.800 469.800 ;
        RECT 92.400 468.600 95.400 469.200 ;
        RECT 120.600 468.600 126.000 469.200 ;
        RECT 155.400 468.600 158.400 469.200 ;
        RECT 165.600 468.600 169.200 469.200 ;
        RECT 45.000 468.000 48.600 468.600 ;
        RECT 91.800 468.000 95.400 468.600 ;
        RECT 120.000 468.000 126.000 468.600 ;
        RECT 156.000 468.000 158.400 468.600 ;
        RECT 45.600 467.400 48.600 468.000 ;
        RECT 91.200 467.400 94.800 468.000 ;
        RECT 118.800 467.400 125.400 468.000 ;
        RECT 156.000 467.400 159.000 468.000 ;
        RECT 166.200 467.400 169.800 468.600 ;
        RECT 180.000 468.000 183.600 469.200 ;
        RECT 188.400 468.600 194.400 469.200 ;
        RECT 204.600 468.600 208.200 469.200 ;
        RECT 188.400 468.000 195.600 468.600 ;
        RECT 204.000 468.000 208.200 468.600 ;
        RECT 179.400 467.400 183.000 468.000 ;
        RECT 188.400 467.400 196.800 468.000 ;
        RECT 202.800 467.400 207.600 468.000 ;
        RECT 214.200 467.400 217.200 468.000 ;
        RECT 45.600 466.800 49.200 467.400 ;
        RECT 91.200 466.800 94.200 467.400 ;
        RECT 118.200 466.800 125.400 467.400 ;
        RECT 156.600 466.800 159.600 467.400 ;
        RECT 166.800 466.800 170.400 467.400 ;
        RECT 179.400 466.800 182.400 467.400 ;
        RECT 46.200 465.600 49.800 466.800 ;
        RECT 90.600 466.200 94.200 466.800 ;
        RECT 117.600 466.200 124.800 466.800 ;
        RECT 156.600 466.200 160.200 466.800 ;
        RECT 167.400 466.200 170.400 466.800 ;
        RECT 178.800 466.200 182.400 466.800 ;
        RECT 187.800 466.800 198.600 467.400 ;
        RECT 200.400 466.800 207.000 467.400 ;
        RECT 212.400 466.800 219.000 467.400 ;
        RECT 187.800 466.200 206.400 466.800 ;
        RECT 211.200 466.200 219.600 466.800 ;
        RECT 90.600 465.600 93.600 466.200 ;
        RECT 117.000 465.600 124.800 466.200 ;
        RECT 157.200 465.600 160.800 466.200 ;
        RECT 167.400 465.600 171.000 466.200 ;
        RECT 178.800 465.600 181.800 466.200 ;
        RECT 46.800 465.000 50.400 465.600 ;
        RECT 47.400 464.400 50.400 465.000 ;
        RECT 90.000 465.000 93.600 465.600 ;
        RECT 116.400 465.000 124.200 465.600 ;
        RECT 90.000 464.400 93.000 465.000 ;
        RECT 115.800 464.400 124.200 465.000 ;
        RECT 157.800 465.000 161.400 465.600 ;
        RECT 168.000 465.000 171.600 465.600 ;
        RECT 178.200 465.000 181.800 465.600 ;
        RECT 187.800 465.000 190.800 466.200 ;
        RECT 192.600 465.600 205.200 466.200 ;
        RECT 210.600 465.600 220.800 466.200 ;
        RECT 193.800 465.000 204.600 465.600 ;
        RECT 210.000 465.000 221.400 465.600 ;
        RECT 157.800 464.400 162.000 465.000 ;
        RECT 168.600 464.400 172.200 465.000 ;
        RECT 178.200 464.400 181.200 465.000 ;
        RECT 47.400 463.800 51.000 464.400 ;
        RECT 48.000 463.200 51.000 463.800 ;
        RECT 89.400 463.800 93.000 464.400 ;
        RECT 115.200 463.800 119.400 464.400 ;
        RECT 89.400 463.200 92.400 463.800 ;
        RECT 114.600 463.200 118.800 463.800 ;
        RECT 48.000 462.600 51.600 463.200 ;
        RECT 88.800 462.600 92.400 463.200 ;
        RECT 114.000 462.600 118.200 463.200 ;
        RECT 120.600 462.600 123.600 464.400 ;
        RECT 158.400 463.800 162.600 464.400 ;
        RECT 168.600 463.800 172.800 464.400 ;
        RECT 159.000 463.200 163.200 463.800 ;
        RECT 169.200 463.200 172.800 463.800 ;
        RECT 177.600 463.800 181.200 464.400 ;
        RECT 187.200 463.800 190.800 465.000 ;
        RECT 195.600 464.400 202.800 465.000 ;
        RECT 209.400 464.400 214.200 465.000 ;
        RECT 216.600 464.400 222.000 465.000 ;
        RECT 192.600 463.800 193.200 464.400 ;
        RECT 197.400 463.800 201.600 464.400 ;
        RECT 208.800 463.800 213.000 464.400 ;
        RECT 218.400 463.800 222.600 464.400 ;
        RECT 159.000 462.600 163.800 463.200 ;
        RECT 169.800 462.600 173.400 463.200 ;
        RECT 177.600 462.600 180.600 463.800 ;
        RECT 186.600 463.200 195.000 463.800 ;
        RECT 198.000 463.200 201.600 463.800 ;
        RECT 208.200 463.200 212.400 463.800 ;
        RECT 219.000 463.200 222.600 463.800 ;
        RECT 186.600 462.600 195.600 463.200 ;
        RECT 198.000 462.600 202.200 463.200 ;
        RECT 48.600 462.000 52.200 462.600 ;
        RECT 49.200 461.400 52.200 462.000 ;
        RECT 88.800 461.400 91.800 462.600 ;
        RECT 113.400 462.000 117.600 462.600 ;
        RECT 49.200 460.800 52.800 461.400 ;
        RECT 49.800 460.200 52.800 460.800 ;
        RECT 88.200 460.800 91.800 461.400 ;
        RECT 112.800 461.400 117.000 462.000 ;
        RECT 112.800 460.800 116.400 461.400 ;
        RECT 49.800 459.600 53.400 460.200 ;
        RECT 50.400 459.000 54.000 459.600 ;
        RECT 88.200 459.000 91.200 460.800 ;
        RECT 112.200 460.200 115.800 460.800 ;
        RECT 111.600 459.000 115.200 460.200 ;
        RECT 120.000 459.600 123.000 462.600 ;
        RECT 157.800 462.000 164.400 462.600 ;
        RECT 170.400 462.000 174.600 462.600 ;
        RECT 156.000 461.400 159.600 462.000 ;
        RECT 161.400 461.400 165.000 462.000 ;
        RECT 171.000 461.400 175.200 462.000 ;
        RECT 154.800 460.800 159.000 461.400 ;
        RECT 162.600 460.800 165.000 461.400 ;
        RECT 171.600 460.800 175.800 461.400 ;
        RECT 154.200 460.200 158.400 460.800 ;
        RECT 153.000 459.600 157.800 460.200 ;
        RECT 172.200 459.600 175.800 460.800 ;
        RECT 120.000 459.000 122.400 459.600 ;
        RECT 152.400 459.000 156.600 459.600 ;
        RECT 171.600 459.000 175.800 459.600 ;
        RECT 177.000 459.000 180.000 462.600 ;
        RECT 186.000 462.000 196.200 462.600 ;
        RECT 198.600 462.000 202.200 462.600 ;
        RECT 207.600 462.600 211.800 463.200 ;
        RECT 219.600 462.600 223.200 463.200 ;
        RECT 207.600 462.000 211.200 462.600 ;
        RECT 186.000 461.400 196.800 462.000 ;
        RECT 199.200 461.400 202.800 462.000 ;
        RECT 207.000 461.400 210.600 462.000 ;
        RECT 220.200 461.400 223.800 462.600 ;
        RECT 185.400 460.800 197.400 461.400 ;
        RECT 184.800 460.200 192.600 460.800 ;
        RECT 193.800 460.200 198.000 460.800 ;
        RECT 199.800 460.200 203.400 461.400 ;
        RECT 206.400 460.200 210.000 461.400 ;
        RECT 220.800 460.800 223.800 461.400 ;
        RECT 184.200 459.600 187.800 460.200 ;
        RECT 183.000 459.000 187.800 459.600 ;
        RECT 189.000 459.000 192.000 460.200 ;
        RECT 194.400 459.600 198.600 460.200 ;
        RECT 200.400 459.600 204.000 460.200 ;
        RECT 205.800 459.600 209.400 460.200 ;
        RECT 195.000 459.000 199.200 459.600 ;
        RECT 201.000 459.000 204.600 459.600 ;
        RECT 205.800 459.000 208.800 459.600 ;
        RECT 221.400 459.000 224.400 460.800 ;
        RECT 51.000 458.400 54.000 459.000 ;
        RECT 51.000 457.800 54.600 458.400 ;
        RECT 51.600 456.600 55.200 457.800 ;
        RECT 52.200 456.000 55.800 456.600 ;
        RECT 87.600 456.000 90.600 459.000 ;
        RECT 111.000 458.400 114.600 459.000 ;
        RECT 110.400 457.800 114.000 458.400 ;
        RECT 110.400 457.200 113.400 457.800 ;
        RECT 109.800 456.600 113.400 457.200 ;
        RECT 109.800 456.000 112.800 456.600 ;
        RECT 52.800 454.800 56.400 456.000 ;
        RECT 53.400 454.200 57.000 454.800 ;
        RECT 54.000 453.000 57.600 454.200 ;
        RECT 54.600 452.400 58.200 453.000 ;
        RECT 55.200 451.200 58.800 452.400 ;
        RECT 87.000 451.200 90.000 456.000 ;
        RECT 109.200 455.400 112.800 456.000 ;
        RECT 119.400 455.400 122.400 459.000 ;
        RECT 151.800 458.400 156.000 459.000 ;
        RECT 171.000 458.400 175.200 459.000 ;
        RECT 177.000 458.400 187.200 459.000 ;
        RECT 151.200 457.800 155.400 458.400 ;
        RECT 171.000 457.800 174.600 458.400 ;
        RECT 177.600 457.800 186.600 458.400 ;
        RECT 150.000 457.200 154.800 457.800 ;
        RECT 170.400 457.200 174.000 457.800 ;
        RECT 177.600 457.200 185.400 457.800 ;
        RECT 149.400 456.600 154.200 457.200 ;
        RECT 169.800 456.600 174.000 457.200 ;
        RECT 178.200 456.600 184.800 457.200 ;
        RECT 188.400 456.600 192.000 459.000 ;
        RECT 195.600 458.400 199.800 459.000 ;
        RECT 201.600 458.400 208.800 459.000 ;
        RECT 196.200 457.800 200.400 458.400 ;
        RECT 201.600 457.800 208.200 458.400 ;
        RECT 196.800 457.200 201.000 457.800 ;
        RECT 148.800 456.000 153.000 456.600 ;
        RECT 169.800 456.000 173.400 456.600 ;
        RECT 179.400 456.000 183.600 456.600 ;
        RECT 148.800 455.400 152.400 456.000 ;
        RECT 169.800 455.400 172.800 456.000 ;
        RECT 109.200 454.800 112.200 455.400 ;
        RECT 108.600 454.200 112.200 454.800 ;
        RECT 120.000 454.800 122.400 455.400 ;
        RECT 148.200 454.800 151.800 455.400 ;
        RECT 169.200 454.800 172.800 455.400 ;
        RECT 189.000 454.800 192.000 456.600 ;
        RECT 197.400 456.600 201.000 457.200 ;
        RECT 202.200 457.200 208.200 457.800 ;
        RECT 202.200 456.600 207.600 457.200 ;
        RECT 197.400 456.000 207.600 456.600 ;
        RECT 198.000 455.400 207.600 456.000 ;
        RECT 198.600 454.800 207.000 455.400 ;
        RECT 108.600 453.600 111.600 454.200 ;
        RECT 108.000 453.000 111.600 453.600 ;
        RECT 108.000 452.400 111.000 453.000 ;
        RECT 120.000 452.400 123.000 454.800 ;
        RECT 147.600 454.200 151.200 454.800 ;
        RECT 147.000 453.600 150.600 454.200 ;
        RECT 146.400 453.000 150.000 453.600 ;
        RECT 169.200 453.000 172.200 454.800 ;
        RECT 145.800 452.400 150.000 453.000 ;
        RECT 155.400 452.400 156.000 453.000 ;
        RECT 55.800 450.600 59.400 451.200 ;
        RECT 87.600 450.600 90.000 451.200 ;
        RECT 107.400 451.800 111.000 452.400 ;
        RECT 107.400 450.600 110.400 451.800 ;
        RECT 56.400 449.400 60.000 450.600 ;
        RECT 57.000 448.800 60.600 449.400 ;
        RECT 57.600 447.600 61.200 448.800 ;
        RECT 87.600 448.200 90.600 450.600 ;
        RECT 106.800 450.000 110.400 450.600 ;
        RECT 120.600 450.600 123.000 452.400 ;
        RECT 145.200 451.800 149.400 452.400 ;
        RECT 145.200 451.200 148.800 451.800 ;
        RECT 155.400 451.200 156.600 452.400 ;
        RECT 168.600 451.200 172.200 453.000 ;
        RECT 189.000 454.200 194.400 454.800 ;
        RECT 189.000 453.600 195.000 454.200 ;
        RECT 199.200 453.600 207.000 454.800 ;
        RECT 189.000 453.000 195.600 453.600 ;
        RECT 199.800 453.000 206.400 453.600 ;
        RECT 222.000 453.000 225.000 459.000 ;
        RECT 189.000 452.400 196.800 453.000 ;
        RECT 189.000 451.800 197.400 452.400 ;
        RECT 189.600 451.200 197.400 451.800 ;
        RECT 200.400 451.800 204.000 453.000 ;
        RECT 200.400 451.200 204.600 451.800 ;
        RECT 221.400 451.200 224.400 453.000 ;
        RECT 144.600 450.600 148.200 451.200 ;
        RECT 106.800 448.800 109.800 450.000 ;
        RECT 120.600 448.800 123.600 450.600 ;
        RECT 144.000 449.400 147.600 450.600 ;
        RECT 155.400 450.000 157.200 451.200 ;
        RECT 143.400 448.800 147.000 449.400 ;
        RECT 155.400 448.800 157.800 450.000 ;
        RECT 106.200 448.200 109.800 448.800 ;
        RECT 58.200 447.000 61.800 447.600 ;
        RECT 58.800 446.400 62.400 447.000 ;
        RECT 88.200 446.400 91.200 448.200 ;
        RECT 106.200 446.400 109.200 448.200 ;
        RECT 121.200 447.600 123.600 448.800 ;
        RECT 142.800 448.200 146.400 448.800 ;
        RECT 156.000 448.200 157.800 448.800 ;
        RECT 142.800 447.600 145.800 448.200 ;
        RECT 59.400 445.200 63.000 446.400 ;
        RECT 88.800 445.200 91.800 446.400 ;
        RECT 60.000 444.600 63.600 445.200 ;
        RECT 88.800 444.600 92.400 445.200 ;
        RECT 60.600 444.000 64.200 444.600 ;
        RECT 89.400 444.000 93.000 444.600 ;
        RECT 60.600 443.400 64.800 444.000 ;
        RECT 61.200 442.800 64.800 443.400 ;
        RECT 90.000 443.400 93.000 444.000 ;
        RECT 90.000 442.800 93.600 443.400 ;
        RECT 61.800 442.200 65.400 442.800 ;
        RECT 90.600 442.200 94.200 442.800 ;
        RECT 62.400 441.600 66.000 442.200 ;
        RECT 90.600 441.600 94.800 442.200 ;
        RECT 63.000 441.000 66.600 441.600 ;
        RECT 91.200 441.000 95.400 441.600 ;
        RECT 63.000 440.400 67.200 441.000 ;
        RECT 91.800 440.400 96.000 441.000 ;
        RECT 63.600 439.800 67.200 440.400 ;
        RECT 92.400 439.800 96.600 440.400 ;
        RECT 64.200 439.200 67.800 439.800 ;
        RECT 93.000 439.200 97.200 439.800 ;
        RECT 64.800 438.600 68.400 439.200 ;
        RECT 93.000 438.600 97.800 439.200 ;
        RECT 64.800 438.000 69.000 438.600 ;
        RECT 93.000 438.000 98.400 438.600 ;
        RECT 65.400 437.400 69.600 438.000 ;
        RECT 66.000 436.800 69.600 437.400 ;
        RECT 92.400 437.400 99.600 438.000 ;
        RECT 105.600 437.400 108.600 446.400 ;
        RECT 121.200 445.800 124.200 447.600 ;
        RECT 142.200 447.000 145.800 447.600 ;
        RECT 142.200 446.400 145.200 447.000 ;
        RECT 141.600 445.800 145.200 446.400 ;
        RECT 156.000 445.800 158.400 448.200 ;
        RECT 121.800 444.000 124.800 445.800 ;
        RECT 141.000 445.200 144.600 445.800 ;
        RECT 141.000 444.600 144.000 445.200 ;
        RECT 140.400 444.000 144.000 444.600 ;
        RECT 121.800 443.400 125.400 444.000 ;
        RECT 140.400 443.400 143.400 444.000 ;
        RECT 122.400 442.200 125.400 443.400 ;
        RECT 139.800 442.800 143.400 443.400 ;
        RECT 122.400 441.600 126.000 442.200 ;
        RECT 139.800 441.600 142.800 442.800 ;
        RECT 123.000 440.400 126.000 441.600 ;
        RECT 139.200 440.400 142.200 441.600 ;
        RECT 123.600 439.200 126.600 440.400 ;
        RECT 138.600 439.800 142.200 440.400 ;
        RECT 138.600 439.200 141.600 439.800 ;
        RECT 123.600 438.600 127.200 439.200 ;
        RECT 92.400 436.800 100.800 437.400 ;
        RECT 66.600 436.200 70.200 436.800 ;
        RECT 92.400 436.200 102.000 436.800 ;
        RECT 67.200 435.600 70.800 436.200 ;
        RECT 92.400 435.600 95.400 436.200 ;
        RECT 97.200 435.600 103.200 436.200 ;
        RECT 106.200 435.600 108.600 437.400 ;
        RECT 123.000 438.000 127.200 438.600 ;
        RECT 138.000 438.600 141.600 439.200 ;
        RECT 123.000 437.400 127.800 438.000 ;
        RECT 138.000 437.400 141.000 438.600 ;
        RECT 123.000 436.800 128.400 437.400 ;
        RECT 122.400 436.200 128.400 436.800 ;
        RECT 137.400 436.200 140.400 437.400 ;
        RECT 156.000 436.800 159.000 445.800 ;
        RECT 168.600 442.200 171.600 451.200 ;
        RECT 189.600 450.600 198.000 451.200 ;
        RECT 189.600 450.000 198.600 450.600 ;
        RECT 201.000 450.000 204.600 451.200 ;
        RECT 220.800 450.600 224.400 451.200 ;
        RECT 220.800 450.000 223.800 450.600 ;
        RECT 189.600 448.200 193.200 450.000 ;
        RECT 194.400 449.400 199.200 450.000 ;
        RECT 195.000 448.800 199.800 449.400 ;
        RECT 201.600 448.800 205.200 450.000 ;
        RECT 220.200 449.400 223.800 450.000 ;
        RECT 220.200 448.800 223.200 449.400 ;
        RECT 195.600 448.200 200.400 448.800 ;
        RECT 189.600 447.600 193.800 448.200 ;
        RECT 196.200 447.600 200.400 448.200 ;
        RECT 202.200 448.200 205.800 448.800 ;
        RECT 219.600 448.200 223.200 448.800 ;
        RECT 202.200 447.600 206.400 448.200 ;
        RECT 219.000 447.600 224.400 448.200 ;
        RECT 190.200 445.800 193.800 447.600 ;
        RECT 196.800 447.000 201.000 447.600 ;
        RECT 202.800 447.000 206.400 447.600 ;
        RECT 217.200 447.000 226.200 447.600 ;
        RECT 197.400 446.400 201.600 447.000 ;
        RECT 203.400 446.400 207.000 447.000 ;
        RECT 216.000 446.400 226.800 447.000 ;
        RECT 197.400 445.800 202.200 446.400 ;
        RECT 190.800 445.200 193.800 445.800 ;
        RECT 198.000 445.200 202.200 445.800 ;
        RECT 204.000 445.800 207.600 446.400 ;
        RECT 216.000 445.800 227.400 446.400 ;
        RECT 204.000 445.200 208.200 445.800 ;
        RECT 190.800 444.000 194.400 445.200 ;
        RECT 198.600 444.600 202.800 445.200 ;
        RECT 204.600 444.600 208.200 445.200 ;
        RECT 216.000 445.200 228.000 445.800 ;
        RECT 216.000 444.600 220.200 445.200 ;
        RECT 224.400 444.600 228.000 445.200 ;
        RECT 191.400 443.400 194.400 444.000 ;
        RECT 199.200 443.400 203.400 444.600 ;
        RECT 205.200 444.000 208.800 444.600 ;
        RECT 205.800 443.400 209.400 444.000 ;
        RECT 191.400 442.800 195.000 443.400 ;
        RECT 199.800 442.800 204.000 443.400 ;
        RECT 205.800 442.800 210.000 443.400 ;
        RECT 225.000 442.800 228.000 444.600 ;
        RECT 192.000 442.200 195.000 442.800 ;
        RECT 200.400 442.200 204.000 442.800 ;
        RECT 206.400 442.200 210.000 442.800 ;
        RECT 224.400 442.200 228.000 442.800 ;
        RECT 168.600 441.000 171.000 442.200 ;
        RECT 192.000 441.600 195.600 442.200 ;
        RECT 200.400 441.600 204.600 442.200 ;
        RECT 207.000 441.600 210.600 442.200 ;
        RECT 224.400 441.600 227.400 442.200 ;
        RECT 156.000 436.200 158.400 436.800 ;
        RECT 122.400 435.600 129.000 436.200 ;
        RECT 136.800 435.600 140.400 436.200 ;
        RECT 67.800 435.000 71.400 435.600 ;
        RECT 67.800 434.400 72.000 435.000 ;
        RECT 68.400 433.800 72.600 434.400 ;
        RECT 69.000 433.200 73.200 433.800 ;
        RECT 69.600 432.600 73.800 433.200 ;
        RECT 70.200 432.000 73.800 432.600 ;
        RECT 70.800 431.400 74.400 432.000 ;
        RECT 71.400 430.800 75.000 431.400 ;
        RECT 72.000 430.200 75.600 430.800 ;
        RECT 72.000 429.600 76.200 430.200 ;
        RECT 72.600 429.000 76.800 429.600 ;
        RECT 73.200 428.400 77.400 429.000 ;
        RECT 73.800 427.800 78.000 428.400 ;
        RECT 74.400 427.200 78.600 427.800 ;
        RECT 75.000 426.600 79.200 427.200 ;
        RECT 75.600 426.000 79.800 426.600 ;
        RECT 76.200 425.400 80.400 426.000 ;
        RECT 76.800 424.800 81.000 425.400 ;
        RECT 77.400 424.200 81.600 424.800 ;
        RECT 91.800 424.200 94.800 435.600 ;
        RECT 97.800 435.000 104.400 435.600 ;
        RECT 106.200 435.000 109.200 435.600 ;
        RECT 121.800 435.000 129.600 435.600 ;
        RECT 136.800 435.000 139.800 435.600 ;
        RECT 99.000 434.400 109.200 435.000 ;
        RECT 100.200 433.800 109.200 434.400 ;
        RECT 121.200 433.800 124.800 435.000 ;
        RECT 126.000 434.400 130.200 435.000 ;
        RECT 136.200 434.400 139.800 435.000 ;
        RECT 126.600 433.800 130.800 434.400 ;
        RECT 135.600 433.800 139.200 434.400 ;
        RECT 155.400 433.800 158.400 436.200 ;
        RECT 168.000 436.200 171.000 441.000 ;
        RECT 192.600 441.000 195.600 441.600 ;
        RECT 201.000 441.000 205.200 441.600 ;
        RECT 207.600 441.000 211.200 441.600 ;
        RECT 223.800 441.000 227.400 441.600 ;
        RECT 192.600 440.400 196.200 441.000 ;
        RECT 201.600 440.400 205.200 441.000 ;
        RECT 208.200 440.400 211.200 441.000 ;
        RECT 223.200 440.400 226.800 441.000 ;
        RECT 193.200 439.800 196.200 440.400 ;
        RECT 193.200 439.200 196.800 439.800 ;
        RECT 202.200 439.200 205.800 440.400 ;
        RECT 208.800 439.800 211.800 440.400 ;
        RECT 222.600 439.800 226.800 440.400 ;
        RECT 210.000 439.200 211.800 439.800 ;
        RECT 222.000 439.200 226.200 439.800 ;
        RECT 193.800 438.600 196.800 439.200 ;
        RECT 202.800 438.600 205.800 439.200 ;
        RECT 210.600 438.600 211.800 439.200 ;
        RECT 221.400 438.600 225.600 439.200 ;
        RECT 193.800 438.000 197.400 438.600 ;
        RECT 202.800 438.000 206.400 438.600 ;
        RECT 220.200 438.000 225.600 438.600 ;
        RECT 228.600 438.000 231.600 438.600 ;
        RECT 194.400 436.800 198.000 438.000 ;
        RECT 203.400 436.800 206.400 438.000 ;
        RECT 219.600 437.400 232.200 438.000 ;
        RECT 218.400 436.800 232.800 437.400 ;
        RECT 195.000 436.200 198.600 436.800 ;
        RECT 168.000 435.600 170.400 436.200 ;
        RECT 101.400 433.200 109.200 433.800 ;
        RECT 102.600 432.600 108.600 433.200 ;
        RECT 120.600 432.600 124.200 433.800 ;
        RECT 127.200 433.200 131.400 433.800 ;
        RECT 135.000 433.200 139.200 433.800 ;
        RECT 127.800 432.600 132.600 433.200 ;
        RECT 134.400 432.600 138.600 433.200 ;
        RECT 104.400 432.000 108.000 432.600 ;
        RECT 120.000 431.400 123.600 432.600 ;
        RECT 128.400 432.000 138.000 432.600 ;
        RECT 154.800 432.000 157.800 433.800 ;
        RECT 129.000 431.400 137.400 432.000 ;
        RECT 119.400 430.200 123.000 431.400 ;
        RECT 129.600 430.800 136.800 431.400 ;
        RECT 130.800 430.200 136.200 430.800 ;
        RECT 154.200 430.200 157.800 432.000 ;
        RECT 167.400 430.200 170.400 435.600 ;
        RECT 195.600 435.000 199.200 436.200 ;
        RECT 196.200 434.400 199.800 435.000 ;
        RECT 196.800 433.800 200.400 434.400 ;
        RECT 203.400 433.800 207.000 436.800 ;
        RECT 217.200 436.200 233.400 436.800 ;
        RECT 216.600 435.600 233.400 436.200 ;
        RECT 216.600 435.000 228.600 435.600 ;
        RECT 218.400 434.400 226.200 435.000 ;
        RECT 230.400 434.400 233.400 435.600 ;
        RECT 197.400 433.200 201.000 433.800 ;
        RECT 202.800 433.200 207.000 433.800 ;
        RECT 197.400 432.600 206.400 433.200 ;
        RECT 198.000 432.000 206.400 432.600 ;
        RECT 199.200 431.400 207.600 432.000 ;
        RECT 200.400 430.800 209.400 431.400 ;
        RECT 204.000 430.200 210.600 430.800 ;
        RECT 118.800 429.000 122.400 430.200 ;
        RECT 132.600 429.600 134.400 430.200 ;
        RECT 153.600 429.600 158.400 430.200 ;
        RECT 167.400 429.600 169.800 430.200 ;
        RECT 205.800 429.600 212.400 430.200 ;
        RECT 153.600 429.000 159.000 429.600 ;
        RECT 118.200 428.400 122.400 429.000 ;
        RECT 153.000 428.400 159.600 429.000 ;
        RECT 118.200 427.800 123.000 428.400 ;
        RECT 117.600 427.200 123.000 427.800 ;
        RECT 153.000 427.800 160.200 428.400 ;
        RECT 153.000 427.200 161.400 427.800 ;
        RECT 117.000 426.000 123.600 427.200 ;
        RECT 152.400 426.000 155.400 427.200 ;
        RECT 157.200 426.600 162.000 427.200 ;
        RECT 157.800 426.000 163.200 426.600 ;
        RECT 116.400 425.400 120.000 426.000 ;
        RECT 115.800 424.800 119.400 425.400 ;
        RECT 115.200 424.200 118.800 424.800 ;
        RECT 121.200 424.200 124.200 426.000 ;
        RECT 151.800 425.400 155.400 426.000 ;
        RECT 159.000 425.400 164.400 426.000 ;
        RECT 151.800 424.800 154.800 425.400 ;
        RECT 159.600 424.800 165.600 425.400 ;
        RECT 166.800 424.800 169.800 429.600 ;
        RECT 207.600 429.000 213.600 429.600 ;
        RECT 209.400 428.400 214.800 429.000 ;
        RECT 210.600 427.800 216.600 428.400 ;
        RECT 231.000 427.800 234.000 434.400 ;
        RECT 211.800 427.200 217.800 427.800 ;
        RECT 213.600 426.600 219.000 427.200 ;
        RECT 214.800 426.000 220.200 426.600 ;
        RECT 216.000 425.400 221.400 426.000 ;
        RECT 230.400 425.400 233.400 427.800 ;
        RECT 535.800 426.000 546.600 426.600 ;
        RECT 529.800 425.400 553.800 426.000 ;
        RECT 217.200 424.800 222.600 425.400 ;
        RECT 151.200 424.200 154.800 424.800 ;
        RECT 160.200 424.200 169.800 424.800 ;
        RECT 219.000 424.200 223.800 424.800 ;
        RECT 229.800 424.200 232.800 425.400 ;
        RECT 526.800 424.800 558.600 425.400 ;
        RECT 524.400 424.200 562.200 424.800 ;
        RECT 78.000 423.600 82.200 424.200 ;
        RECT 92.400 423.600 94.800 424.200 ;
        RECT 114.600 423.600 118.800 424.200 ;
        RECT 78.600 423.000 82.800 423.600 ;
        RECT 79.200 422.400 83.400 423.000 ;
        RECT 79.800 421.800 84.000 422.400 ;
        RECT 92.400 421.800 95.400 423.600 ;
        RECT 114.600 423.000 118.200 423.600 ;
        RECT 114.000 422.400 117.600 423.000 ;
        RECT 113.400 421.800 117.000 422.400 ;
        RECT 121.800 421.800 124.800 424.200 ;
        RECT 150.600 423.600 154.800 424.200 ;
        RECT 161.400 423.600 169.800 424.200 ;
        RECT 220.200 423.600 224.400 424.200 ;
        RECT 229.200 423.600 232.800 424.200 ;
        RECT 522.000 423.600 565.200 424.200 ;
        RECT 150.600 423.000 155.400 423.600 ;
        RECT 162.600 423.000 169.800 423.600 ;
        RECT 221.400 423.000 225.600 423.600 ;
        RECT 228.600 423.000 232.200 423.600 ;
        RECT 520.200 423.000 534.600 423.600 ;
        RECT 547.800 423.000 567.600 423.600 ;
        RECT 150.000 422.400 155.400 423.000 ;
        RECT 163.200 422.400 169.800 423.000 ;
        RECT 222.000 422.400 226.800 423.000 ;
        RECT 228.000 422.400 232.200 423.000 ;
        RECT 518.400 422.400 529.800 423.000 ;
        RECT 554.400 422.400 570.600 423.000 ;
        RECT 150.000 421.800 156.000 422.400 ;
        RECT 163.200 421.800 169.200 422.400 ;
        RECT 223.200 421.800 231.600 422.400 ;
        RECT 516.600 421.800 526.800 422.400 ;
        RECT 558.600 421.800 572.400 422.400 ;
        RECT 80.400 421.200 84.600 421.800 ;
        RECT 92.400 421.200 96.000 421.800 ;
        RECT 112.800 421.200 116.400 421.800 ;
        RECT 81.000 420.600 85.200 421.200 ;
        RECT 81.600 420.000 85.800 420.600 ;
        RECT 93.000 420.000 96.000 421.200 ;
        RECT 112.200 420.600 116.400 421.200 ;
        RECT 111.600 420.000 115.800 420.600 ;
        RECT 82.200 419.400 86.400 420.000 ;
        RECT 93.000 419.400 96.600 420.000 ;
        RECT 82.800 418.800 87.000 419.400 ;
        RECT 93.600 418.800 96.600 419.400 ;
        RECT 111.000 419.400 115.200 420.000 ;
        RECT 111.000 418.800 114.600 419.400 ;
        RECT 122.400 418.800 125.400 421.800 ;
        RECT 149.400 421.200 156.000 421.800 ;
        RECT 148.800 420.600 156.000 421.200 ;
        RECT 163.800 421.200 168.600 421.800 ;
        RECT 224.400 421.200 231.000 421.800 ;
        RECT 515.400 421.200 524.400 421.800 ;
        RECT 562.200 421.200 574.200 421.800 ;
        RECT 163.800 420.600 168.000 421.200 ;
        RECT 225.000 420.600 229.800 421.200 ;
        RECT 514.200 420.600 522.000 421.200 ;
        RECT 565.200 420.600 576.000 421.200 ;
        RECT 148.800 420.000 156.600 420.600 ;
        RECT 164.400 420.000 168.000 420.600 ;
        RECT 226.200 420.000 229.800 420.600 ;
        RECT 513.000 420.000 520.200 420.600 ;
        RECT 567.600 420.000 577.800 420.600 ;
        RECT 148.200 419.400 156.600 420.000 ;
        RECT 83.400 418.200 88.200 418.800 ;
        RECT 93.600 418.200 97.200 418.800 ;
        RECT 110.400 418.200 114.000 418.800 ;
        RECT 84.000 417.600 88.800 418.200 ;
        RECT 94.200 417.600 97.200 418.200 ;
        RECT 109.800 417.600 113.400 418.200 ;
        RECT 84.600 417.000 89.400 417.600 ;
        RECT 94.200 417.000 97.800 417.600 ;
        RECT 109.200 417.000 112.800 417.600 ;
        RECT 85.800 416.400 90.000 417.000 ;
        RECT 94.800 416.400 97.800 417.000 ;
        RECT 108.600 416.400 112.200 417.000 ;
        RECT 86.400 415.800 90.600 416.400 ;
        RECT 94.800 415.800 98.400 416.400 ;
        RECT 108.000 415.800 112.200 416.400 ;
        RECT 123.000 415.800 126.000 418.800 ;
        RECT 147.600 418.200 151.200 419.400 ;
        RECT 152.400 418.800 156.600 419.400 ;
        RECT 165.000 419.400 168.000 420.000 ;
        RECT 226.800 419.400 229.800 420.000 ;
        RECT 511.200 419.400 519.000 420.000 ;
        RECT 570.000 419.400 579.000 420.000 ;
        RECT 165.000 418.800 168.600 419.400 ;
        RECT 227.400 418.800 230.400 419.400 ;
        RECT 510.600 418.800 517.200 419.400 ;
        RECT 571.800 418.800 580.200 419.400 ;
        RECT 153.000 418.200 156.600 418.800 ;
        RECT 165.600 418.200 169.200 418.800 ;
        RECT 228.000 418.200 231.000 418.800 ;
        RECT 509.400 418.200 516.000 418.800 ;
        RECT 573.600 418.200 582.000 418.800 ;
        RECT 147.000 417.600 150.600 418.200 ;
        RECT 153.000 417.600 157.200 418.200 ;
        RECT 146.400 416.400 150.000 417.600 ;
        RECT 145.800 415.800 149.400 416.400 ;
        RECT 87.000 415.200 91.800 415.800 ;
        RECT 95.400 415.200 99.000 415.800 ;
        RECT 107.400 415.200 111.600 415.800 ;
        RECT 87.600 414.600 92.400 415.200 ;
        RECT 96.000 414.600 99.000 415.200 ;
        RECT 106.800 414.600 111.000 415.200 ;
        RECT 87.600 414.000 93.000 414.600 ;
        RECT 96.000 414.000 99.600 414.600 ;
        RECT 106.200 414.000 110.400 414.600 ;
        RECT 87.600 413.400 94.200 414.000 ;
        RECT 96.600 413.400 100.200 414.000 ;
        RECT 105.600 413.400 109.800 414.000 ;
        RECT 86.400 412.800 94.800 413.400 ;
        RECT 97.200 412.800 101.400 413.400 ;
        RECT 104.400 412.800 108.600 413.400 ;
        RECT 123.600 412.800 126.600 415.800 ;
        RECT 145.200 414.600 148.800 415.800 ;
        RECT 153.600 415.200 157.200 417.600 ;
        RECT 166.200 417.600 169.200 418.200 ;
        RECT 228.600 417.600 231.000 418.200 ;
        RECT 508.200 417.600 514.200 418.200 ;
        RECT 575.400 417.600 583.200 418.200 ;
        RECT 166.200 417.000 169.800 417.600 ;
        RECT 228.600 417.000 231.600 417.600 ;
        RECT 507.000 417.000 513.000 417.600 ;
        RECT 576.600 417.000 584.400 417.600 ;
        RECT 166.800 416.400 169.800 417.000 ;
        RECT 167.400 415.800 169.800 416.400 ;
        RECT 229.200 416.400 231.600 417.000 ;
        RECT 506.400 416.400 511.800 417.000 ;
        RECT 578.400 416.400 586.200 417.000 ;
        RECT 229.200 415.800 232.200 416.400 ;
        RECT 505.200 415.800 511.200 416.400 ;
        RECT 579.600 415.800 587.400 416.400 ;
        RECT 168.000 415.200 170.400 415.800 ;
        RECT 144.600 414.000 148.200 414.600 ;
        RECT 154.200 414.000 157.200 415.200 ;
        RECT 168.600 414.600 169.800 415.200 ;
        RECT 229.800 414.600 232.200 415.800 ;
        RECT 504.000 415.200 510.000 415.800 ;
        RECT 581.400 415.200 588.600 415.800 ;
        RECT 503.400 414.600 508.800 415.200 ;
        RECT 582.600 414.600 589.800 415.200 ;
        RECT 230.400 414.000 232.200 414.600 ;
        RECT 502.200 414.000 507.600 414.600 ;
        RECT 584.400 414.000 591.000 414.600 ;
        RECT 144.000 413.400 147.600 414.000 ;
        RECT 85.800 412.200 95.400 412.800 ;
        RECT 97.800 412.200 108.000 412.800 ;
        RECT 124.200 412.200 126.600 412.800 ;
        RECT 143.400 412.200 147.000 413.400 ;
        RECT 84.600 411.600 89.400 412.200 ;
        RECT 91.200 411.600 96.600 412.200 ;
        RECT 98.400 411.600 107.400 412.200 ;
        RECT 84.000 411.000 88.800 411.600 ;
        RECT 92.400 411.000 97.200 411.600 ;
        RECT 99.000 411.000 106.800 411.600 ;
        RECT 82.800 410.400 88.200 411.000 ;
        RECT 93.000 410.400 98.400 411.000 ;
        RECT 99.600 410.400 106.200 411.000 ;
        RECT 81.600 409.800 87.000 410.400 ;
        RECT 94.200 409.800 99.000 410.400 ;
        RECT 101.400 409.800 105.000 410.400 ;
        RECT 81.000 409.200 86.400 409.800 ;
        RECT 94.800 409.200 99.600 409.800 ;
        RECT 101.400 409.200 104.400 409.800 ;
        RECT 124.200 409.200 127.200 412.200 ;
        RECT 142.800 411.600 146.400 412.200 ;
        RECT 142.200 411.000 145.800 411.600 ;
        RECT 141.600 410.400 145.200 411.000 ;
        RECT 141.000 409.800 145.200 410.400 ;
        RECT 141.000 409.200 144.600 409.800 ;
        RECT 79.800 408.600 85.200 409.200 ;
        RECT 96.000 408.600 104.400 409.200 ;
        RECT 78.600 408.000 84.600 408.600 ;
        RECT 96.600 408.000 104.400 408.600 ;
        RECT 78.000 407.400 83.400 408.000 ;
        RECT 97.800 407.400 104.400 408.000 ;
        RECT 76.800 406.800 82.200 407.400 ;
        RECT 98.400 406.800 104.400 407.400 ;
        RECT 76.200 406.200 81.600 406.800 ;
        RECT 99.600 406.200 104.400 406.800 ;
        RECT 75.000 405.600 80.400 406.200 ;
        RECT 100.800 405.600 104.400 406.200 ;
        RECT 124.800 408.600 127.200 409.200 ;
        RECT 140.400 408.600 144.000 409.200 ;
        RECT 154.200 408.600 157.800 414.000 ;
        RECT 230.400 409.800 232.800 414.000 ;
        RECT 501.600 413.400 507.000 414.000 ;
        RECT 585.600 413.400 592.200 414.000 ;
        RECT 501.000 412.800 505.800 413.400 ;
        RECT 586.800 412.800 593.400 413.400 ;
        RECT 500.400 412.200 505.200 412.800 ;
        RECT 588.000 412.200 594.600 412.800 ;
        RECT 499.800 411.600 504.000 412.200 ;
        RECT 589.200 411.600 595.800 412.200 ;
        RECT 499.200 411.000 503.400 411.600 ;
        RECT 590.400 411.000 597.000 411.600 ;
        RECT 498.000 410.400 502.800 411.000 ;
        RECT 591.600 410.400 598.200 411.000 ;
        RECT 497.400 409.800 501.600 410.400 ;
        RECT 592.800 409.800 599.400 410.400 ;
        RECT 231.000 408.600 232.800 409.800 ;
        RECT 496.800 409.200 501.000 409.800 ;
        RECT 594.000 409.200 600.600 409.800 ;
        RECT 496.200 408.600 500.400 409.200 ;
        RECT 595.200 408.600 601.200 409.200 ;
        RECT 124.800 405.600 127.800 408.600 ;
        RECT 139.800 408.000 143.400 408.600 ;
        RECT 139.200 407.400 142.800 408.000 ;
        RECT 154.200 407.400 157.200 408.600 ;
        RECT 138.600 406.800 142.800 407.400 ;
        RECT 138.000 406.200 142.200 406.800 ;
        RECT 137.400 405.600 141.600 406.200 ;
        RECT 153.600 405.600 157.200 407.400 ;
        RECT 73.800 405.000 79.800 405.600 ;
        RECT 73.200 404.400 78.600 405.000 ;
        RECT 72.000 403.800 77.400 404.400 ;
        RECT 71.400 403.200 76.800 403.800 ;
        RECT 70.200 402.600 75.600 403.200 ;
        RECT 69.600 402.000 75.000 402.600 ;
        RECT 68.400 401.400 73.800 402.000 ;
        RECT 67.800 400.800 73.200 401.400 ;
        RECT 66.600 400.200 72.000 400.800 ;
        RECT 66.000 399.600 71.400 400.200 ;
        RECT 64.800 399.000 70.200 399.600 ;
        RECT 64.200 398.400 69.600 399.000 ;
        RECT 63.600 397.800 68.400 398.400 ;
        RECT 62.400 397.200 67.800 397.800 ;
        RECT 61.800 396.600 66.600 397.200 ;
        RECT 101.400 396.600 104.400 405.600 ;
        RECT 125.400 403.800 128.400 405.600 ;
        RECT 136.800 405.000 141.600 405.600 ;
        RECT 153.000 405.000 156.600 405.600 ;
        RECT 136.200 404.400 142.200 405.000 ;
        RECT 152.400 404.400 156.600 405.000 ;
        RECT 135.600 403.800 142.800 404.400 ;
        RECT 152.400 403.800 156.000 404.400 ;
        RECT 126.000 402.600 129.000 403.800 ;
        RECT 135.000 403.200 143.400 403.800 ;
        RECT 151.200 403.200 156.000 403.800 ;
        RECT 134.400 402.600 144.600 403.200 ;
        RECT 150.600 402.600 155.400 403.200 ;
        RECT 126.000 402.000 129.600 402.600 ;
        RECT 133.200 402.000 138.000 402.600 ;
        RECT 139.200 402.000 146.400 402.600 ;
        RECT 148.200 402.000 154.800 402.600 ;
        RECT 230.400 402.000 232.800 408.600 ;
        RECT 495.600 408.000 499.200 408.600 ;
        RECT 596.400 408.000 602.400 408.600 ;
        RECT 495.000 407.400 498.600 408.000 ;
        RECT 597.600 407.400 603.600 408.000 ;
        RECT 494.400 406.800 498.000 407.400 ;
        RECT 598.800 406.800 604.800 407.400 ;
        RECT 493.800 406.200 497.400 406.800 ;
        RECT 599.400 406.200 606.000 406.800 ;
        RECT 493.200 405.600 496.800 406.200 ;
        RECT 600.600 405.600 607.200 406.200 ;
        RECT 492.600 405.000 496.200 405.600 ;
        RECT 601.800 405.000 608.400 405.600 ;
        RECT 492.000 404.400 496.200 405.000 ;
        RECT 603.000 404.400 609.600 405.000 ;
        RECT 491.400 403.800 495.600 404.400 ;
        RECT 604.200 403.800 610.800 404.400 ;
        RECT 491.400 403.200 495.000 403.800 ;
        RECT 605.400 403.200 612.000 403.800 ;
        RECT 490.800 402.600 494.400 403.200 ;
        RECT 606.600 402.600 613.200 403.200 ;
        RECT 490.200 402.000 493.800 402.600 ;
        RECT 607.800 402.000 614.400 402.600 ;
        RECT 126.600 401.400 130.800 402.000 ;
        RECT 132.000 401.400 137.400 402.000 ;
        RECT 140.400 401.400 154.200 402.000 ;
        RECT 229.800 401.400 232.800 402.000 ;
        RECT 489.600 401.400 493.800 402.000 ;
        RECT 609.000 401.400 615.000 402.000 ;
        RECT 126.600 400.800 136.800 401.400 ;
        RECT 141.000 400.800 153.600 401.400 ;
        RECT 127.200 400.200 135.600 400.800 ;
        RECT 142.200 400.200 153.000 400.800 ;
        RECT 127.800 399.600 135.000 400.200 ;
        RECT 143.400 399.600 152.400 400.200 ;
        RECT 229.800 399.600 232.200 401.400 ;
        RECT 489.600 400.800 493.200 401.400 ;
        RECT 610.200 400.800 616.200 401.400 ;
        RECT 489.000 400.200 492.600 400.800 ;
        RECT 611.400 400.200 617.400 400.800 ;
        RECT 129.000 399.000 133.800 399.600 ;
        RECT 144.600 399.000 151.200 399.600 ;
        RECT 129.600 397.800 132.600 399.000 ;
        RECT 147.600 398.400 149.400 399.000 ;
        RECT 229.200 398.400 232.200 399.600 ;
        RECT 488.400 399.000 492.000 400.200 ;
        RECT 612.600 399.600 618.600 400.200 ;
        RECT 613.200 399.000 619.200 399.600 ;
        RECT 487.800 398.400 491.400 399.000 ;
        RECT 614.400 398.400 620.400 399.000 ;
        RECT 60.600 396.000 66.000 396.600 ;
        RECT 60.000 395.400 64.800 396.000 ;
        RECT 58.800 394.800 64.200 395.400 ;
        RECT 58.200 394.200 63.000 394.800 ;
        RECT 57.000 393.600 62.400 394.200 ;
        RECT 102.000 393.600 105.000 396.600 ;
        RECT 130.200 396.000 133.200 397.800 ;
        RECT 229.200 397.200 231.600 398.400 ;
        RECT 487.800 397.800 490.800 398.400 ;
        RECT 615.600 397.800 621.000 398.400 ;
        RECT 487.200 397.200 490.800 397.800 ;
        RECT 616.800 397.200 622.200 397.800 ;
        RECT 228.600 396.600 231.600 397.200 ;
        RECT 486.600 396.600 490.200 397.200 ;
        RECT 617.400 396.600 622.800 397.200 ;
        RECT 130.800 394.200 133.800 396.000 ;
        RECT 225.000 395.400 226.800 396.000 ;
        RECT 228.600 395.400 231.000 396.600 ;
        RECT 486.600 396.000 489.600 396.600 ;
        RECT 534.000 396.000 537.000 396.600 ;
        RECT 618.600 396.000 624.000 396.600 ;
        RECT 222.000 394.800 231.000 395.400 ;
        RECT 486.000 395.400 489.600 396.000 ;
        RECT 529.200 395.400 541.200 396.000 ;
        RECT 619.800 395.400 624.600 396.000 ;
        RECT 486.000 394.800 489.000 395.400 ;
        RECT 526.800 394.800 543.600 395.400 ;
        RECT 620.400 394.800 625.800 395.400 ;
        RECT 220.200 394.200 230.400 394.800 ;
        RECT 56.400 393.000 61.800 393.600 ;
        RECT 55.800 392.400 60.600 393.000 ;
        RECT 102.600 392.400 105.600 393.600 ;
        RECT 131.400 393.000 134.400 394.200 ;
        RECT 218.400 393.600 230.400 394.200 ;
        RECT 485.400 394.200 489.000 394.800 ;
        RECT 525.000 394.200 546.000 394.800 ;
        RECT 621.600 394.200 626.400 394.800 ;
        RECT 485.400 393.600 488.400 394.200 ;
        RECT 523.800 393.600 547.200 394.200 ;
        RECT 622.800 393.600 627.600 394.200 ;
        RECT 217.200 393.000 229.800 393.600 ;
        RECT 131.400 392.400 135.000 393.000 ;
        RECT 216.000 392.400 224.400 393.000 ;
        RECT 226.800 392.400 229.800 393.000 ;
        RECT 484.800 393.000 488.400 393.600 ;
        RECT 522.600 393.000 532.800 393.600 ;
        RECT 537.600 393.000 549.000 393.600 ;
        RECT 623.400 393.000 628.800 393.600 ;
        RECT 484.800 392.400 487.800 393.000 ;
        RECT 521.400 392.400 529.200 393.000 ;
        RECT 541.200 392.400 550.200 393.000 ;
        RECT 624.600 392.400 630.000 393.000 ;
        RECT 54.600 391.800 60.000 392.400 ;
        RECT 79.200 391.800 81.000 392.400 ;
        RECT 102.600 391.800 106.200 392.400 ;
        RECT 54.000 391.200 58.800 391.800 ;
        RECT 78.000 391.200 81.600 391.800 ;
        RECT 100.800 391.200 101.400 391.800 ;
        RECT 52.800 390.600 58.200 391.200 ;
        RECT 76.200 390.600 81.600 391.200 ;
        RECT 100.200 390.600 101.400 391.200 ;
        RECT 103.200 391.200 106.800 391.800 ;
        RECT 132.000 391.200 135.000 392.400 ;
        RECT 214.800 391.800 222.000 392.400 ;
        RECT 213.600 391.200 220.200 391.800 ;
        RECT 226.800 391.200 229.200 392.400 ;
        RECT 484.200 391.200 487.200 392.400 ;
        RECT 520.200 391.800 527.400 392.400 ;
        RECT 543.600 391.800 551.400 392.400 ;
        RECT 625.200 391.800 631.200 392.400 ;
        RECT 519.600 391.200 525.600 391.800 ;
        RECT 545.400 391.200 552.000 391.800 ;
        RECT 626.400 391.200 631.800 391.800 ;
        RECT 103.200 390.600 107.400 391.200 ;
        RECT 132.600 390.600 135.600 391.200 ;
        RECT 213.000 390.600 219.000 391.200 ;
        RECT 226.200 390.600 228.600 391.200 ;
        RECT 52.200 390.000 57.600 390.600 ;
        RECT 75.000 390.000 81.600 390.600 ;
        RECT 99.000 390.000 101.400 390.600 ;
        RECT 103.800 390.000 108.600 390.600 ;
        RECT 133.200 390.000 135.600 390.600 ;
        RECT 211.800 390.000 217.800 390.600 ;
        RECT 225.600 390.000 228.600 390.600 ;
        RECT 483.600 390.000 486.600 391.200 ;
        RECT 518.400 390.600 524.400 391.200 ;
        RECT 547.200 390.600 553.200 391.200 ;
        RECT 627.600 390.600 633.000 391.200 ;
        RECT 517.800 390.000 523.200 390.600 ;
        RECT 548.400 390.000 554.400 390.600 ;
        RECT 628.200 390.000 634.200 390.600 ;
        RECT 51.600 389.400 57.600 390.000 ;
        RECT 73.800 389.400 81.600 390.000 ;
        RECT 98.400 389.400 101.400 390.000 ;
        RECT 104.400 389.400 109.800 390.000 ;
        RECT 134.400 389.400 135.000 390.000 ;
        RECT 211.200 389.400 216.600 390.000 ;
        RECT 225.600 389.400 228.000 390.000 ;
        RECT 483.000 389.400 486.600 390.000 ;
        RECT 517.200 389.400 522.000 390.000 ;
        RECT 549.600 389.400 555.000 390.000 ;
        RECT 629.400 389.400 634.800 390.000 ;
        RECT 50.400 388.800 57.600 389.400 ;
        RECT 72.600 388.800 81.000 389.400 ;
        RECT 97.800 388.800 102.600 389.400 ;
        RECT 104.400 388.800 113.400 389.400 ;
        RECT 118.800 388.800 126.000 389.400 ;
        RECT 210.600 388.800 215.400 389.400 ;
        RECT 225.000 388.800 228.000 389.400 ;
        RECT 49.800 388.200 57.600 388.800 ;
        RECT 71.400 388.200 77.400 388.800 ;
        RECT 49.200 387.600 57.600 388.200 ;
        RECT 70.200 387.600 76.800 388.200 ;
        RECT 48.000 387.000 52.800 387.600 ;
        RECT 47.400 386.400 52.200 387.000 ;
        RECT 46.200 385.800 51.600 386.400 ;
        RECT 45.600 385.200 50.400 385.800 ;
        RECT 54.600 385.200 57.600 387.600 ;
        RECT 69.000 387.000 75.600 387.600 ;
        RECT 78.600 387.000 81.000 388.800 ;
        RECT 97.200 388.200 126.000 388.800 ;
        RECT 210.000 388.200 214.800 388.800 ;
        RECT 225.000 388.200 227.400 388.800 ;
        RECT 96.600 387.600 124.800 388.200 ;
        RECT 209.400 387.600 214.200 388.200 ;
        RECT 224.400 387.600 227.400 388.200 ;
        RECT 482.400 388.200 486.000 389.400 ;
        RECT 516.600 388.800 521.400 389.400 ;
        RECT 550.800 388.800 556.200 389.400 ;
        RECT 630.000 388.800 636.000 389.400 ;
        RECT 516.000 388.200 520.200 388.800 ;
        RECT 551.400 388.200 556.800 388.800 ;
        RECT 631.200 388.200 636.600 388.800 ;
        RECT 482.400 387.600 485.400 388.200 ;
        RECT 515.400 387.600 519.600 388.200 ;
        RECT 552.600 387.600 557.400 388.200 ;
        RECT 632.400 387.600 637.800 388.200 ;
        RECT 96.000 387.000 123.600 387.600 ;
        RECT 208.800 387.000 213.600 387.600 ;
        RECT 223.800 387.000 226.800 387.600 ;
        RECT 67.800 386.400 74.400 387.000 ;
        RECT 66.600 385.800 73.200 386.400 ;
        RECT 64.800 385.200 72.000 385.800 ;
        RECT 45.000 384.600 49.800 385.200 ;
        RECT 54.600 384.600 58.200 385.200 ;
        RECT 63.000 384.600 70.800 385.200 ;
        RECT 78.600 384.600 81.600 387.000 ;
        RECT 94.800 386.400 99.600 387.000 ;
        RECT 100.800 386.400 121.800 387.000 ;
        RECT 208.200 386.400 213.000 387.000 ;
        RECT 223.200 386.400 226.800 387.000 ;
        RECT 481.800 387.000 485.400 387.600 ;
        RECT 514.800 387.000 519.000 387.600 ;
        RECT 553.200 387.000 558.000 387.600 ;
        RECT 633.000 387.000 639.000 387.600 ;
        RECT 481.800 386.400 484.800 387.000 ;
        RECT 514.200 386.400 518.400 387.000 ;
        RECT 554.400 386.400 558.600 387.000 ;
        RECT 634.200 386.400 639.600 387.000 ;
        RECT 94.200 385.800 99.000 386.400 ;
        RECT 102.000 385.800 109.200 386.400 ;
        RECT 114.000 385.800 121.200 386.400 ;
        RECT 207.600 385.800 212.400 386.400 ;
        RECT 223.200 385.800 226.200 386.400 ;
        RECT 93.600 385.200 98.400 385.800 ;
        RECT 105.000 385.200 106.800 385.800 ;
        RECT 92.400 384.600 97.200 385.200 ;
        RECT 43.800 384.000 49.200 384.600 ;
        RECT 54.600 384.000 69.600 384.600 ;
        RECT 79.200 384.000 82.200 384.600 ;
        RECT 91.200 384.000 96.600 384.600 ;
        RECT 105.000 384.000 106.200 385.200 ;
        RECT 117.600 384.600 121.200 385.800 ;
        RECT 207.000 385.200 211.800 385.800 ;
        RECT 222.600 385.200 225.600 385.800 ;
        RECT 481.200 385.200 484.800 386.400 ;
        RECT 513.600 385.800 517.800 386.400 ;
        RECT 555.000 385.800 559.200 386.400 ;
        RECT 635.400 385.800 640.800 386.400 ;
        RECT 513.000 385.200 517.200 385.800 ;
        RECT 555.600 385.200 559.800 385.800 ;
        RECT 636.000 385.200 641.400 385.800 ;
        RECT 206.400 384.600 211.200 385.200 ;
        RECT 222.000 384.600 225.000 385.200 ;
        RECT 481.200 384.600 484.200 385.200 ;
        RECT 513.000 384.600 516.600 385.200 ;
        RECT 556.200 384.600 560.400 385.200 ;
        RECT 637.200 384.600 642.600 385.200 ;
        RECT 117.000 384.000 120.600 384.600 ;
        RECT 205.800 384.000 210.600 384.600 ;
        RECT 221.400 384.000 225.000 384.600 ;
        RECT 43.200 383.400 48.000 384.000 ;
        RECT 55.200 383.400 68.400 384.000 ;
        RECT 79.200 383.400 82.800 384.000 ;
        RECT 90.000 383.400 96.000 384.000 ;
        RECT 105.000 383.400 106.800 384.000 ;
        RECT 116.400 383.400 120.000 384.000 ;
        RECT 205.200 383.400 210.000 384.000 ;
        RECT 220.800 383.400 224.400 384.000 ;
        RECT 42.000 382.800 47.400 383.400 ;
        RECT 55.800 382.800 66.600 383.400 ;
        RECT 79.800 382.800 83.400 383.400 ;
        RECT 88.800 382.800 94.800 383.400 ;
        RECT 41.400 382.200 46.200 382.800 ;
        RECT 56.400 382.200 64.800 382.800 ;
        RECT 79.800 382.200 94.200 382.800 ;
        RECT 105.000 382.200 107.400 383.400 ;
        RECT 115.800 382.800 120.000 383.400 ;
        RECT 204.600 382.800 208.800 383.400 ;
        RECT 219.600 382.800 223.800 383.400 ;
        RECT 480.600 382.800 484.200 384.600 ;
        RECT 512.400 384.000 516.000 384.600 ;
        RECT 556.800 384.000 561.000 384.600 ;
        RECT 637.800 384.000 643.200 384.600 ;
        RECT 511.800 383.400 515.400 384.000 ;
        RECT 558.000 383.400 561.600 384.000 ;
        RECT 639.000 383.400 644.400 384.000 ;
        RECT 511.800 382.800 514.800 383.400 ;
        RECT 558.000 382.800 562.200 383.400 ;
        RECT 639.600 382.800 645.000 383.400 ;
        RECT 115.200 382.200 119.400 382.800 ;
        RECT 163.800 382.200 166.200 382.800 ;
        RECT 203.400 382.200 208.200 382.800 ;
        RECT 219.000 382.200 223.200 382.800 ;
        RECT 40.800 381.600 45.600 382.200 ;
        RECT 57.000 381.600 63.000 382.200 ;
        RECT 67.800 381.600 71.400 382.200 ;
        RECT 80.400 381.600 93.000 382.200 ;
        RECT 39.600 381.000 45.000 381.600 ;
        RECT 66.000 381.000 71.400 381.600 ;
        RECT 81.000 381.000 91.800 381.600 ;
        RECT 39.000 380.400 43.800 381.000 ;
        RECT 64.200 380.400 71.400 381.000 ;
        RECT 81.600 380.400 90.600 381.000 ;
        RECT 105.000 380.400 108.000 382.200 ;
        RECT 114.600 381.600 118.800 382.200 ;
        RECT 163.200 381.600 167.400 382.200 ;
        RECT 202.800 381.600 207.600 382.200 ;
        RECT 218.400 381.600 222.600 382.200 ;
        RECT 114.000 381.000 118.200 381.600 ;
        RECT 163.200 381.000 169.200 381.600 ;
        RECT 202.200 381.000 207.000 381.600 ;
        RECT 217.800 381.000 222.000 381.600 ;
        RECT 480.000 381.000 483.600 382.800 ;
        RECT 511.200 382.200 514.800 382.800 ;
        RECT 558.600 382.200 562.800 382.800 ;
        RECT 640.800 382.200 646.200 382.800 ;
        RECT 510.600 381.600 514.200 382.200 ;
        RECT 559.200 381.600 563.400 382.200 ;
        RECT 641.400 381.600 646.800 382.200 ;
        RECT 510.600 381.000 513.600 381.600 ;
        RECT 559.800 381.000 563.400 381.600 ;
        RECT 642.600 381.000 648.000 381.600 ;
        RECT 112.800 380.400 117.600 381.000 ;
        RECT 163.800 380.400 171.000 381.000 ;
        RECT 201.000 380.400 206.400 381.000 ;
        RECT 217.200 380.400 221.400 381.000 ;
        RECT 480.000 380.400 483.000 381.000 ;
        RECT 38.400 379.800 43.200 380.400 ;
        RECT 63.600 379.800 71.400 380.400 ;
        RECT 82.800 379.800 88.800 380.400 ;
        RECT 37.200 379.200 42.000 379.800 ;
        RECT 63.000 379.200 70.200 379.800 ;
        RECT 104.400 379.200 107.400 380.400 ;
        RECT 112.200 379.800 117.000 380.400 ;
        RECT 164.400 379.800 172.800 380.400 ;
        RECT 199.800 379.800 205.800 380.400 ;
        RECT 216.000 379.800 220.800 380.400 ;
        RECT 111.000 379.200 116.400 379.800 ;
        RECT 165.600 379.200 174.600 379.800 ;
        RECT 198.600 379.200 204.600 379.800 ;
        RECT 215.400 379.200 220.200 379.800 ;
        RECT 36.600 378.600 41.400 379.200 ;
        RECT 63.000 378.600 67.800 379.200 ;
        RECT 91.800 378.600 93.000 379.200 ;
        RECT 103.800 378.600 107.400 379.200 ;
        RECT 110.400 378.600 115.200 379.200 ;
        RECT 133.200 378.600 133.800 379.200 ;
        RECT 167.400 378.600 177.000 379.200 ;
        RECT 196.800 378.600 204.000 379.200 ;
        RECT 214.800 378.600 219.000 379.200 ;
        RECT 479.400 378.600 483.000 380.400 ;
        RECT 510.000 380.400 513.600 381.000 ;
        RECT 560.400 380.400 564.000 381.000 ;
        RECT 643.200 380.400 648.600 381.000 ;
        RECT 510.000 379.200 513.000 380.400 ;
        RECT 561.000 379.200 564.600 380.400 ;
        RECT 644.400 379.800 649.200 380.400 ;
        RECT 645.000 379.200 650.400 379.800 ;
        RECT 35.400 378.000 40.800 378.600 ;
        RECT 34.800 377.400 39.600 378.000 ;
        RECT 34.200 376.800 39.000 377.400 ;
        RECT 33.000 376.200 38.400 376.800 ;
        RECT 63.000 376.200 66.000 378.600 ;
        RECT 91.200 378.000 93.600 378.600 ;
        RECT 103.200 378.000 106.800 378.600 ;
        RECT 91.200 376.800 94.200 378.000 ;
        RECT 102.600 377.400 106.800 378.000 ;
        RECT 109.800 377.400 114.600 378.600 ;
        RECT 130.800 378.000 134.400 378.600 ;
        RECT 168.600 378.000 179.400 378.600 ;
        RECT 194.400 378.000 202.800 378.600 ;
        RECT 213.600 378.000 218.400 378.600 ;
        RECT 479.400 378.000 482.400 378.600 ;
        RECT 129.000 377.400 133.800 378.000 ;
        RECT 170.400 377.400 181.800 378.000 ;
        RECT 191.400 377.400 201.600 378.000 ;
        RECT 213.000 377.400 217.200 378.000 ;
        RECT 102.000 376.800 106.200 377.400 ;
        RECT 109.800 376.800 116.400 377.400 ;
        RECT 126.600 376.800 133.200 377.400 ;
        RECT 172.200 376.800 200.400 377.400 ;
        RECT 211.800 376.800 216.600 377.400 ;
        RECT 79.800 376.200 81.600 376.800 ;
        RECT 90.000 376.200 94.800 376.800 ;
        RECT 101.400 376.200 105.600 376.800 ;
        RECT 110.400 376.200 121.200 376.800 ;
        RECT 122.400 376.200 132.600 376.800 ;
        RECT 174.000 376.200 198.600 376.800 ;
        RECT 211.200 376.200 216.000 376.800 ;
        RECT 478.800 376.200 482.400 378.000 ;
        RECT 509.400 377.400 512.400 379.200 ;
        RECT 561.600 378.600 565.200 379.200 ;
        RECT 646.200 378.600 651.000 379.200 ;
        RECT 562.200 378.000 565.800 378.600 ;
        RECT 646.800 378.000 651.600 378.600 ;
        RECT 562.800 377.400 565.800 378.000 ;
        RECT 647.400 377.400 652.800 378.000 ;
        RECT 32.400 375.600 37.200 376.200 ;
        RECT 63.000 375.600 66.600 376.200 ;
        RECT 78.600 375.600 82.800 376.200 ;
        RECT 88.200 375.600 94.800 376.200 ;
        RECT 100.200 375.600 105.000 376.200 ;
        RECT 111.000 375.600 131.400 376.200 ;
        RECT 176.400 375.600 196.800 376.200 ;
        RECT 210.000 375.600 214.800 376.200 ;
        RECT 31.200 375.000 36.600 375.600 ;
        RECT 63.600 375.000 66.600 375.600 ;
        RECT 76.800 375.000 84.600 375.600 ;
        RECT 86.400 375.000 95.400 375.600 ;
        RECT 99.000 375.000 104.400 375.600 ;
        RECT 112.200 375.000 130.200 375.600 ;
        RECT 178.800 375.000 195.000 375.600 ;
        RECT 208.800 375.000 214.200 375.600 ;
        RECT 478.800 375.000 481.800 376.200 ;
        RECT 508.800 375.000 511.800 377.400 ;
        RECT 562.800 376.800 566.400 377.400 ;
        RECT 648.600 376.800 653.400 377.400 ;
        RECT 563.400 376.200 566.400 376.800 ;
        RECT 649.200 376.200 654.000 376.800 ;
        RECT 563.400 375.600 567.000 376.200 ;
        RECT 649.800 375.600 654.600 376.200 ;
        RECT 564.000 375.000 567.000 375.600 ;
        RECT 651.000 375.000 655.800 375.600 ;
        RECT 30.600 374.400 35.400 375.000 ;
        RECT 63.600 374.400 67.200 375.000 ;
        RECT 75.600 374.400 91.200 375.000 ;
        RECT 92.400 374.400 96.000 375.000 ;
        RECT 97.800 374.400 103.800 375.000 ;
        RECT 114.000 374.400 129.000 375.000 ;
        RECT 182.400 374.400 191.400 375.000 ;
        RECT 207.000 374.400 213.000 375.000 ;
        RECT 29.400 373.800 34.800 374.400 ;
        RECT 64.200 373.800 67.800 374.400 ;
        RECT 73.800 373.800 90.600 374.400 ;
        RECT 92.400 373.800 102.600 374.400 ;
        RECT 116.400 373.800 129.000 374.400 ;
        RECT 205.200 373.800 211.800 374.400 ;
        RECT 28.800 373.200 34.200 373.800 ;
        RECT 64.200 373.200 90.000 373.800 ;
        RECT 93.000 373.200 102.000 373.800 ;
        RECT 28.200 372.600 33.000 373.200 ;
        RECT 64.800 372.600 78.600 373.200 ;
        RECT 82.200 372.600 88.800 373.200 ;
        RECT 93.600 372.600 100.800 373.200 ;
        RECT 27.000 372.000 32.400 372.600 ;
        RECT 65.400 372.000 77.400 372.600 ;
        RECT 84.600 372.000 86.400 372.600 ;
        RECT 94.200 372.000 99.600 372.600 ;
        RECT 124.800 372.000 128.400 373.800 ;
        RECT 202.800 373.200 210.600 373.800 ;
        RECT 478.200 373.200 481.800 375.000 ;
        RECT 147.000 372.600 148.800 373.200 ;
        RECT 159.000 372.600 169.800 373.200 ;
        RECT 199.200 372.600 208.800 373.200 ;
        RECT 142.800 372.000 150.000 372.600 ;
        RECT 159.000 372.000 176.400 372.600 ;
        RECT 193.200 372.000 207.000 372.600 ;
        RECT 478.200 372.000 481.200 373.200 ;
        RECT 26.400 371.400 31.200 372.000 ;
        RECT 66.600 371.400 76.200 372.000 ;
        RECT 95.400 371.400 97.800 372.000 ;
        RECT 123.600 371.400 127.800 372.000 ;
        RECT 140.400 371.400 149.400 372.000 ;
        RECT 159.600 371.400 205.200 372.000 ;
        RECT 25.200 370.800 30.600 371.400 ;
        RECT 67.800 370.800 73.800 371.400 ;
        RECT 123.000 370.800 127.800 371.400 ;
        RECT 138.600 370.800 147.600 371.400 ;
        RECT 161.400 370.800 202.800 371.400 ;
        RECT 24.600 370.200 29.400 370.800 ;
        RECT 121.800 370.200 127.200 370.800 ;
        RECT 136.200 370.200 146.400 370.800 ;
        RECT 164.400 370.200 200.400 370.800 ;
        RECT 23.400 369.600 28.800 370.200 ;
        RECT 120.600 369.600 126.600 370.200 ;
        RECT 134.400 369.600 144.600 370.200 ;
        RECT 169.800 369.600 195.600 370.200 ;
        RECT 222.600 369.600 227.400 370.200 ;
        RECT 22.800 369.000 27.600 369.600 ;
        RECT 118.800 369.000 126.600 369.600 ;
        RECT 132.000 369.000 143.400 369.600 ;
        RECT 177.000 369.000 179.400 369.600 ;
        RECT 184.800 369.000 188.400 369.600 ;
        RECT 218.400 369.000 231.600 369.600 ;
        RECT 477.600 369.000 481.200 372.000 ;
        RECT 21.600 368.400 27.000 369.000 ;
        RECT 117.600 368.400 126.600 369.000 ;
        RECT 129.000 368.400 143.400 369.000 ;
        RECT 21.000 367.800 27.000 368.400 ;
        RECT 116.400 367.800 138.600 368.400 ;
        RECT 19.800 367.200 42.600 367.800 ;
        RECT 115.200 367.200 122.400 367.800 ;
        RECT 123.600 367.200 136.200 367.800 ;
        RECT 141.000 367.200 144.000 368.400 ;
        RECT 185.400 367.800 188.400 369.000 ;
        RECT 216.000 368.400 234.000 369.000 ;
        RECT 214.200 367.800 235.800 368.400 ;
        RECT 261.000 367.800 264.000 368.400 ;
        RECT 185.400 367.200 189.000 367.800 ;
        RECT 212.400 367.200 237.000 367.800 ;
        RECT 260.400 367.200 264.600 367.800 ;
        RECT 477.600 367.200 480.600 369.000 ;
        RECT 18.600 366.600 51.000 367.200 ;
        RECT 114.000 366.600 121.200 367.200 ;
        RECT 123.600 366.600 134.400 367.200 ;
        RECT 141.600 366.600 144.600 367.200 ;
        RECT 186.000 366.600 189.000 367.200 ;
        RECT 211.200 366.600 222.000 367.200 ;
        RECT 228.000 366.600 238.200 367.200 ;
        RECT 259.800 366.600 265.200 367.200 ;
        RECT 18.000 366.000 56.400 366.600 ;
        RECT 112.200 366.000 120.000 366.600 ;
        RECT 124.200 366.000 132.000 366.600 ;
        RECT 141.600 366.000 145.200 366.600 ;
        RECT 186.000 366.000 189.600 366.600 ;
        RECT 210.000 366.000 218.400 366.600 ;
        RECT 231.600 366.000 239.400 366.600 ;
        RECT 259.800 366.000 265.800 366.600 ;
        RECT 17.400 365.400 60.000 366.000 ;
        RECT 111.000 365.400 118.800 366.000 ;
        RECT 125.400 365.400 129.000 366.000 ;
        RECT 142.200 365.400 145.200 366.000 ;
        RECT 186.600 365.400 189.600 366.000 ;
        RECT 208.800 365.400 216.000 366.000 ;
        RECT 233.400 365.400 240.600 366.000 ;
        RECT 259.800 365.400 266.400 366.000 ;
        RECT 17.400 364.800 63.600 365.400 ;
        RECT 109.200 364.800 117.600 365.400 ;
        RECT 142.200 364.800 145.800 365.400 ;
        RECT 186.600 364.800 190.200 365.400 ;
        RECT 207.600 364.800 214.200 365.400 ;
        RECT 235.200 364.800 241.200 365.400 ;
        RECT 259.200 364.800 266.400 365.400 ;
        RECT 43.800 364.200 66.600 364.800 ;
        RECT 108.000 364.200 115.800 364.800 ;
        RECT 51.600 363.600 69.600 364.200 ;
        RECT 106.200 363.600 114.600 364.200 ;
        RECT 142.800 363.600 145.800 364.800 ;
        RECT 187.200 364.200 190.800 364.800 ;
        RECT 206.400 364.200 213.000 364.800 ;
        RECT 236.400 364.200 242.400 364.800 ;
        RECT 187.200 363.600 192.000 364.200 ;
        RECT 205.200 363.600 211.800 364.200 ;
        RECT 237.600 363.600 243.000 364.200 ;
        RECT 56.400 363.000 73.200 363.600 ;
        RECT 103.800 363.000 113.400 363.600 ;
        RECT 60.600 362.400 76.200 363.000 ;
        RECT 102.000 362.400 112.200 363.000 ;
        RECT 143.400 362.400 146.400 363.600 ;
        RECT 187.800 363.000 192.600 363.600 ;
        RECT 204.000 363.000 210.600 363.600 ;
        RECT 238.800 363.000 243.600 363.600 ;
        RECT 188.400 362.400 193.800 363.000 ;
        RECT 202.800 362.400 209.400 363.000 ;
        RECT 239.400 362.400 244.200 363.000 ;
        RECT 259.200 362.400 262.200 364.800 ;
        RECT 263.400 364.200 267.000 364.800 ;
        RECT 264.000 363.600 267.600 364.200 ;
        RECT 264.600 363.000 267.600 363.600 ;
        RECT 477.000 363.600 480.600 367.200 ;
        RECT 508.200 367.200 511.200 375.000 ;
        RECT 564.000 374.400 567.600 375.000 ;
        RECT 651.600 374.400 656.400 375.000 ;
        RECT 564.600 373.800 567.600 374.400 ;
        RECT 652.200 373.800 657.000 374.400 ;
        RECT 564.600 373.200 568.200 373.800 ;
        RECT 652.800 373.200 657.600 373.800 ;
        RECT 565.200 372.600 568.200 373.200 ;
        RECT 654.000 372.600 658.200 373.200 ;
        RECT 565.200 372.000 568.800 372.600 ;
        RECT 654.600 372.000 658.800 372.600 ;
        RECT 565.800 371.400 568.800 372.000 ;
        RECT 655.200 371.400 660.000 372.000 ;
        RECT 565.800 370.800 569.400 371.400 ;
        RECT 655.800 370.800 660.600 371.400 ;
        RECT 566.400 369.600 569.400 370.800 ;
        RECT 656.400 370.200 661.200 370.800 ;
        RECT 657.600 369.600 661.800 370.200 ;
        RECT 566.400 369.000 570.000 369.600 ;
        RECT 658.200 369.000 662.400 369.600 ;
        RECT 567.000 367.800 570.000 369.000 ;
        RECT 658.800 368.400 663.000 369.000 ;
        RECT 659.400 367.800 663.600 368.400 ;
        RECT 508.200 366.000 510.600 367.200 ;
        RECT 567.600 366.000 570.600 367.800 ;
        RECT 660.000 367.200 664.200 367.800 ;
        RECT 660.600 366.600 664.800 367.200 ;
        RECT 661.200 366.000 665.400 366.600 ;
        RECT 264.600 362.400 268.200 363.000 ;
        RECT 63.600 361.800 79.200 362.400 ;
        RECT 99.600 361.800 110.400 362.400 ;
        RECT 143.400 361.800 147.000 362.400 ;
        RECT 189.000 361.800 195.600 362.400 ;
        RECT 201.600 361.800 208.200 362.400 ;
        RECT 240.600 361.800 244.800 362.400 ;
        RECT 259.200 361.800 261.600 362.400 ;
        RECT 67.200 361.200 84.000 361.800 ;
        RECT 95.400 361.200 108.600 361.800 ;
        RECT 70.200 360.600 107.400 361.200 ;
        RECT 73.200 360.000 105.000 360.600 ;
        RECT 144.000 360.000 147.000 361.800 ;
        RECT 190.200 361.200 207.000 361.800 ;
        RECT 241.200 361.200 245.400 361.800 ;
        RECT 190.800 360.600 206.400 361.200 ;
        RECT 241.800 360.600 246.000 361.200 ;
        RECT 191.400 360.000 205.200 360.600 ;
        RECT 242.400 360.000 246.600 360.600 ;
        RECT 76.200 359.400 103.200 360.000 ;
        RECT 79.800 358.800 99.600 359.400 ;
        RECT 84.000 358.200 94.800 358.800 ;
        RECT 144.600 357.600 147.600 360.000 ;
        RECT 192.600 359.400 204.000 360.000 ;
        RECT 243.000 359.400 246.600 360.000 ;
        RECT 145.200 357.000 147.600 357.600 ;
        RECT 195.600 358.800 202.800 359.400 ;
        RECT 243.600 358.800 247.200 359.400 ;
        RECT 195.600 358.200 201.600 358.800 ;
        RECT 244.200 358.200 247.800 358.800 ;
        RECT 195.600 357.600 200.400 358.200 ;
        RECT 211.200 357.600 212.400 358.200 ;
        RECT 195.600 357.000 199.200 357.600 ;
        RECT 210.000 357.000 213.600 357.600 ;
        RECT 244.800 357.000 248.400 358.200 ;
        RECT 145.200 354.600 148.200 357.000 ;
        RECT 196.200 356.400 198.000 357.000 ;
        RECT 209.400 356.400 214.800 357.000 ;
        RECT 245.400 356.400 249.000 357.000 ;
        RECT 208.800 355.800 215.400 356.400 ;
        RECT 246.000 355.800 249.000 356.400 ;
        RECT 258.600 356.400 261.600 361.800 ;
        RECT 265.200 361.800 268.200 362.400 ;
        RECT 265.200 361.200 268.800 361.800 ;
        RECT 265.800 360.600 268.800 361.200 ;
        RECT 265.800 360.000 269.400 360.600 ;
        RECT 477.000 360.000 480.000 363.600 ;
        RECT 508.200 361.800 511.200 366.000 ;
        RECT 568.200 364.200 571.200 366.000 ;
        RECT 661.800 365.400 666.000 366.000 ;
        RECT 662.400 364.800 666.600 365.400 ;
        RECT 663.000 364.200 667.200 364.800 ;
        RECT 568.800 362.400 571.800 364.200 ;
        RECT 663.600 363.600 667.800 364.200 ;
        RECT 664.200 363.000 668.400 363.600 ;
        RECT 664.800 362.400 669.000 363.000 ;
        RECT 266.400 358.800 269.400 360.000 ;
        RECT 267.000 357.600 270.000 358.800 ;
        RECT 267.000 357.000 270.600 357.600 ;
        RECT 258.600 355.800 261.000 356.400 ;
        RECT 208.200 355.200 216.000 355.800 ;
        RECT 246.000 355.200 249.600 355.800 ;
        RECT 207.600 354.600 216.600 355.200 ;
        RECT 246.600 354.600 249.600 355.200 ;
        RECT 145.200 353.400 147.600 354.600 ;
        RECT 207.000 354.000 210.600 354.600 ;
        RECT 213.000 354.000 217.200 354.600 ;
        RECT 246.600 354.000 250.200 354.600 ;
        RECT 206.400 353.400 210.600 354.000 ;
        RECT 213.600 353.400 217.800 354.000 ;
        RECT 144.600 350.400 147.600 353.400 ;
        RECT 205.800 352.800 210.000 353.400 ;
        RECT 214.200 352.800 217.800 353.400 ;
        RECT 247.200 353.400 250.200 354.000 ;
        RECT 247.200 352.800 250.800 353.400 ;
        RECT 205.800 352.200 209.400 352.800 ;
        RECT 214.800 352.200 218.400 352.800 ;
        RECT 205.200 351.600 208.800 352.200 ;
        RECT 215.400 351.600 218.400 352.200 ;
        RECT 247.800 352.200 250.800 352.800 ;
        RECT 247.800 351.600 251.400 352.200 ;
        RECT 204.600 351.000 208.200 351.600 ;
        RECT 215.400 351.000 219.000 351.600 ;
        RECT 144.000 348.600 147.000 350.400 ;
        RECT 204.000 349.800 207.600 351.000 ;
        RECT 216.000 350.400 219.000 351.000 ;
        RECT 248.400 351.000 251.400 351.600 ;
        RECT 248.400 350.400 252.000 351.000 ;
        RECT 216.000 349.800 219.600 350.400 ;
        RECT 203.400 349.200 207.000 349.800 ;
        RECT 143.400 348.000 149.400 348.600 ;
        RECT 193.800 348.000 195.000 348.600 ;
        RECT 202.800 348.000 206.400 349.200 ;
        RECT 216.600 348.600 219.600 349.800 ;
        RECT 249.000 349.200 252.000 350.400 ;
        RECT 249.000 348.600 252.600 349.200 ;
        RECT 143.400 347.400 150.600 348.000 ;
        RECT 192.600 347.400 196.800 348.000 ;
        RECT 202.200 347.400 205.800 348.000 ;
        RECT 142.200 346.800 150.000 347.400 ;
        RECT 192.000 346.800 198.000 347.400 ;
        RECT 202.200 346.800 205.200 347.400 ;
        RECT 141.000 346.200 149.400 346.800 ;
        RECT 192.000 346.200 199.200 346.800 ;
        RECT 201.600 346.200 205.200 346.800 ;
        RECT 217.200 346.800 220.200 348.600 ;
        RECT 249.600 347.400 252.600 348.600 ;
        RECT 258.000 348.000 261.000 355.800 ;
        RECT 267.600 355.800 270.600 357.000 ;
        RECT 476.400 357.000 480.000 360.000 ;
        RECT 508.800 360.600 511.200 361.800 ;
        RECT 267.600 355.200 271.200 355.800 ;
        RECT 268.200 354.000 271.200 355.200 ;
        RECT 268.800 352.200 271.800 354.000 ;
        RECT 268.800 351.600 272.400 352.200 ;
        RECT 269.400 349.800 272.400 351.600 ;
        RECT 222.000 346.800 229.200 347.400 ;
        RECT 217.200 346.200 235.200 346.800 ;
        RECT 140.400 345.600 148.200 346.200 ;
        RECT 191.400 345.600 199.800 346.200 ;
        RECT 201.000 345.600 204.600 346.200 ;
        RECT 217.200 345.600 238.800 346.200 ;
        RECT 139.200 345.000 146.400 345.600 ;
        RECT 191.400 345.000 204.000 345.600 ;
        RECT 138.000 344.400 145.200 345.000 ;
        RECT 191.400 344.400 194.400 345.000 ;
        RECT 196.200 344.400 204.000 345.000 ;
        RECT 217.200 345.000 241.200 345.600 ;
        RECT 250.200 345.000 253.200 347.400 ;
        RECT 258.000 346.800 260.400 348.000 ;
        RECT 270.000 347.400 273.000 349.800 ;
        RECT 217.200 344.400 243.600 345.000 ;
        RECT 137.400 343.800 143.400 344.400 ;
        RECT 136.200 343.200 142.200 343.800 ;
        RECT 135.000 342.600 141.000 343.200 ;
        RECT 190.800 342.600 193.800 344.400 ;
        RECT 197.400 343.800 203.400 344.400 ;
        RECT 198.600 343.200 203.400 343.800 ;
        RECT 217.200 343.200 220.200 344.400 ;
        RECT 230.400 343.800 245.400 344.400 ;
        RECT 235.800 343.200 247.200 343.800 ;
        RECT 133.800 342.000 140.400 342.600 ;
        RECT 132.600 341.400 139.200 342.000 ;
        RECT 131.400 340.800 138.000 341.400 ;
        RECT 190.200 340.800 193.200 342.600 ;
        RECT 199.200 342.000 203.400 343.200 ;
        RECT 199.800 341.400 203.400 342.000 ;
        RECT 216.600 341.400 219.600 343.200 ;
        RECT 238.800 342.600 248.400 343.200 ;
        RECT 250.800 342.600 253.800 345.000 ;
        RECT 241.200 342.000 249.600 342.600 ;
        RECT 250.800 342.000 254.400 342.600 ;
        RECT 222.600 341.400 224.400 342.000 ;
        RECT 243.600 341.400 254.400 342.000 ;
        RECT 200.400 340.800 203.400 341.400 ;
        RECT 216.000 340.800 219.600 341.400 ;
        RECT 220.800 340.800 225.600 341.400 ;
        RECT 244.800 340.800 254.400 341.400 ;
        RECT 130.200 340.200 136.800 340.800 ;
        RECT 129.600 339.600 135.600 340.200 ;
        RECT 128.400 339.000 134.400 339.600 ;
        RECT 163.200 339.000 171.000 339.600 ;
        RECT 189.600 339.000 192.600 340.800 ;
        RECT 127.200 338.400 133.200 339.000 ;
        RECT 159.000 338.400 170.400 339.000 ;
        RECT 189.000 338.400 192.600 339.000 ;
        RECT 126.600 337.800 132.000 338.400 ;
        RECT 154.800 337.800 169.200 338.400 ;
        RECT 125.400 337.200 131.400 337.800 ;
        RECT 150.600 337.200 167.400 337.800 ;
        RECT 189.000 337.200 192.000 338.400 ;
        RECT 201.000 337.200 204.000 340.800 ;
        RECT 216.000 340.200 226.200 340.800 ;
        RECT 246.600 340.200 254.400 340.800 ;
        RECT 215.400 339.600 226.800 340.200 ;
        RECT 247.800 339.600 255.000 340.200 ;
        RECT 257.400 339.600 260.400 346.800 ;
        RECT 270.600 345.000 273.600 347.400 ;
        RECT 281.400 345.000 284.400 345.600 ;
        RECT 271.200 342.600 274.200 345.000 ;
        RECT 281.400 344.400 285.000 345.000 ;
        RECT 280.800 343.800 285.600 344.400 ;
        RECT 476.400 343.800 479.400 357.000 ;
        RECT 508.800 356.400 511.800 360.600 ;
        RECT 569.400 360.000 572.400 362.400 ;
        RECT 665.400 361.800 669.600 362.400 ;
        RECT 666.000 361.200 670.200 361.800 ;
        RECT 666.600 360.600 670.800 361.200 ;
        RECT 667.200 360.000 671.400 360.600 ;
        RECT 570.000 357.600 573.000 360.000 ;
        RECT 667.800 359.400 672.000 360.000 ;
        RECT 668.400 358.800 672.000 359.400 ;
        RECT 669.000 358.200 672.600 358.800 ;
        RECT 669.600 357.600 673.200 358.200 ;
        RECT 509.400 352.800 512.400 356.400 ;
        RECT 570.600 355.800 573.600 357.600 ;
        RECT 670.200 357.000 673.800 357.600 ;
        RECT 670.200 356.400 674.400 357.000 ;
        RECT 670.800 355.800 675.000 356.400 ;
        RECT 571.200 353.400 574.200 355.800 ;
        RECT 671.400 355.200 675.600 355.800 ;
        RECT 672.000 354.600 675.600 355.200 ;
        RECT 672.600 354.000 676.200 354.600 ;
        RECT 673.200 353.400 676.800 354.000 ;
        RECT 510.000 349.800 513.000 352.800 ;
        RECT 571.800 351.600 574.800 353.400 ;
        RECT 673.800 352.800 677.400 353.400 ;
        RECT 673.800 352.200 678.000 352.800 ;
        RECT 674.400 351.600 678.000 352.200 ;
        RECT 571.800 351.000 575.400 351.600 ;
        RECT 675.000 351.000 678.600 351.600 ;
        RECT 510.600 347.400 513.600 349.800 ;
        RECT 572.400 349.200 575.400 351.000 ;
        RECT 675.600 350.400 679.200 351.000 ;
        RECT 676.200 349.800 679.800 350.400 ;
        RECT 676.200 349.200 680.400 349.800 ;
        RECT 511.200 345.600 514.200 347.400 ;
        RECT 573.000 346.800 576.000 349.200 ;
        RECT 676.800 348.600 680.400 349.200 ;
        RECT 677.400 348.000 681.000 348.600 ;
        RECT 678.000 347.400 681.600 348.000 ;
        RECT 678.000 346.800 682.200 347.400 ;
        RECT 511.800 344.400 514.800 345.600 ;
        RECT 573.600 345.000 576.600 346.800 ;
        RECT 678.600 346.200 682.200 346.800 ;
        RECT 679.200 345.600 682.800 346.200 ;
        RECT 573.600 344.400 577.200 345.000 ;
        RECT 679.800 344.400 683.400 345.600 ;
        RECT 280.200 342.600 286.200 343.800 ;
        RECT 477.000 343.200 479.400 343.800 ;
        RECT 512.400 343.800 514.800 344.400 ;
        RECT 271.800 339.600 274.800 342.600 ;
        RECT 279.600 342.000 286.800 342.600 ;
        RECT 279.600 341.400 282.600 342.000 ;
        RECT 279.000 340.800 282.600 341.400 ;
        RECT 283.800 341.400 286.800 342.000 ;
        RECT 283.800 340.800 287.400 341.400 ;
        RECT 279.000 340.200 282.000 340.800 ;
        RECT 278.400 339.600 282.000 340.200 ;
        RECT 284.400 339.600 287.400 340.800 ;
        RECT 214.800 339.000 226.800 339.600 ;
        RECT 249.600 339.000 255.000 339.600 ;
        RECT 256.800 339.000 260.400 339.600 ;
        RECT 214.800 338.400 222.600 339.000 ;
        RECT 213.600 337.800 220.800 338.400 ;
        RECT 213.000 337.200 219.600 337.800 ;
        RECT 124.800 336.600 130.200 337.200 ;
        RECT 148.200 336.600 165.000 337.200 ;
        RECT 189.000 336.600 191.400 337.200 ;
        RECT 201.000 336.600 203.400 337.200 ;
        RECT 212.400 336.600 218.400 337.200 ;
        RECT 123.600 336.000 129.000 336.600 ;
        RECT 146.400 336.000 162.000 336.600 ;
        RECT 189.600 336.000 190.800 336.600 ;
        RECT 212.400 336.000 217.200 336.600 ;
        RECT 223.800 336.000 226.800 339.000 ;
        RECT 250.200 338.400 259.800 339.000 ;
        RECT 251.400 337.800 259.800 338.400 ;
        RECT 252.600 337.200 259.800 337.800 ;
        RECT 272.400 337.200 275.400 339.600 ;
        RECT 278.400 339.000 281.400 339.600 ;
        RECT 277.800 338.400 281.400 339.000 ;
        RECT 277.800 337.200 280.800 338.400 ;
        RECT 285.000 337.800 288.000 339.600 ;
        RECT 477.000 339.000 480.000 343.200 ;
        RECT 512.400 342.600 515.400 343.800 ;
        RECT 574.200 342.600 577.200 344.400 ;
        RECT 680.400 343.800 684.000 344.400 ;
        RECT 680.400 343.200 684.600 343.800 ;
        RECT 681.000 342.600 684.600 343.200 ;
        RECT 513.000 342.000 515.400 342.600 ;
        RECT 513.000 340.800 516.000 342.000 ;
        RECT 574.800 340.800 577.800 342.600 ;
        RECT 681.600 342.000 685.200 342.600 ;
        RECT 681.600 341.400 685.800 342.000 ;
        RECT 682.200 340.800 685.800 341.400 ;
        RECT 513.600 339.000 516.600 340.800 ;
        RECT 574.800 340.200 578.400 340.800 ;
        RECT 477.600 338.400 480.000 339.000 ;
        RECT 253.200 336.600 259.800 337.200 ;
        RECT 254.400 336.000 259.800 336.600 ;
        RECT 123.000 335.400 128.400 336.000 ;
        RECT 147.000 335.400 158.400 336.000 ;
        RECT 212.400 335.400 216.000 336.000 ;
        RECT 223.200 335.400 226.800 336.000 ;
        RECT 255.000 335.400 259.800 336.000 ;
        RECT 273.000 336.000 276.000 337.200 ;
        RECT 277.200 336.600 280.800 337.200 ;
        RECT 277.200 336.000 280.200 336.600 ;
        RECT 273.000 335.400 280.200 336.000 ;
        RECT 285.600 336.000 288.600 337.800 ;
        RECT 285.600 335.400 289.200 336.000 ;
        RECT 477.600 335.400 480.600 338.400 ;
        RECT 514.200 337.200 517.200 339.000 ;
        RECT 575.400 338.400 578.400 340.200 ;
        RECT 682.800 339.600 686.400 340.800 ;
        RECT 683.400 339.000 687.000 339.600 ;
        RECT 514.800 336.000 517.800 337.200 ;
        RECT 576.000 336.600 579.000 338.400 ;
        RECT 684.000 337.800 687.600 339.000 ;
        RECT 684.600 336.600 688.200 337.800 ;
        RECT 514.800 335.400 518.400 336.000 ;
        RECT 122.400 334.800 127.200 335.400 ;
        RECT 223.200 334.800 226.200 335.400 ;
        RECT 256.200 334.800 260.400 335.400 ;
        RECT 121.800 334.200 126.600 334.800 ;
        RECT 222.600 334.200 226.200 334.800 ;
        RECT 256.800 334.200 261.000 334.800 ;
        RECT 273.000 334.200 279.600 335.400 ;
        RECT 120.600 333.600 125.400 334.200 ;
        RECT 222.000 333.600 225.600 334.200 ;
        RECT 257.400 333.600 261.600 334.200 ;
        RECT 120.000 333.000 124.800 333.600 ;
        RECT 220.800 333.000 225.600 333.600 ;
        RECT 258.000 333.000 262.200 333.600 ;
        RECT 119.400 332.400 124.200 333.000 ;
        RECT 219.000 332.400 225.600 333.000 ;
        RECT 259.200 332.400 262.800 333.000 ;
        RECT 273.600 332.400 279.000 334.200 ;
        RECT 286.200 333.000 289.200 335.400 ;
        RECT 118.800 331.800 123.000 332.400 ;
        RECT 193.800 331.800 208.800 332.400 ;
        RECT 218.400 331.800 227.400 332.400 ;
        RECT 259.800 331.800 263.400 332.400 ;
        RECT 273.600 331.800 278.400 332.400 ;
        RECT 118.200 331.200 122.400 331.800 ;
        RECT 189.600 331.200 212.400 331.800 ;
        RECT 218.400 331.200 228.600 331.800 ;
        RECT 260.400 331.200 264.000 331.800 ;
        RECT 117.600 330.600 121.800 331.200 ;
        RECT 186.600 330.600 214.800 331.200 ;
        RECT 218.400 330.600 229.800 331.200 ;
        RECT 261.000 330.600 264.600 331.200 ;
        RECT 274.200 330.600 278.400 331.800 ;
        RECT 286.800 330.600 289.800 333.000 ;
        RECT 478.200 332.400 481.200 335.400 ;
        RECT 515.400 334.200 518.400 335.400 ;
        RECT 576.600 334.800 579.600 336.600 ;
        RECT 685.200 336.000 688.800 336.600 ;
        RECT 685.800 335.400 688.800 336.000 ;
        RECT 685.800 334.800 689.400 335.400 ;
        RECT 576.600 334.200 580.200 334.800 ;
        RECT 516.000 333.000 519.000 334.200 ;
        RECT 577.200 333.000 580.200 334.200 ;
        RECT 686.400 334.200 689.400 334.800 ;
        RECT 686.400 333.600 690.000 334.200 ;
        RECT 687.000 333.000 690.000 333.600 ;
        RECT 516.000 332.400 519.600 333.000 ;
        RECT 577.200 332.400 580.800 333.000 ;
        RECT 687.000 332.400 690.600 333.000 ;
        RECT 478.200 331.800 481.800 332.400 ;
        RECT 117.000 330.000 121.200 330.600 ;
        RECT 184.200 330.000 216.600 330.600 ;
        RECT 218.400 330.000 230.400 330.600 ;
        RECT 261.000 330.000 265.200 330.600 ;
        RECT 116.400 329.400 120.600 330.000 ;
        RECT 181.800 329.400 199.800 330.000 ;
        RECT 202.800 329.400 220.200 330.000 ;
        RECT 225.600 329.400 231.000 330.000 ;
        RECT 261.600 329.400 265.800 330.000 ;
        RECT 115.800 328.800 120.000 329.400 ;
        RECT 180.000 328.800 193.200 329.400 ;
        RECT 208.800 328.800 220.200 329.400 ;
        RECT 226.800 328.800 231.600 329.400 ;
        RECT 262.200 328.800 265.800 329.400 ;
        RECT 274.200 328.800 277.800 330.600 ;
        RECT 287.400 330.000 289.800 330.600 ;
        RECT 478.800 330.000 481.800 331.800 ;
        RECT 516.600 331.200 519.600 332.400 ;
        RECT 577.800 331.200 580.800 332.400 ;
        RECT 687.600 331.800 691.200 332.400 ;
        RECT 688.200 331.200 691.200 331.800 ;
        RECT 517.200 330.000 520.200 331.200 ;
        RECT 577.800 330.600 581.400 331.200 ;
        RECT 115.800 328.200 119.400 328.800 ;
        RECT 178.200 328.200 189.600 328.800 ;
        RECT 212.400 328.200 221.400 328.800 ;
        RECT 115.200 327.600 118.800 328.200 ;
        RECT 177.600 327.600 186.600 328.200 ;
        RECT 214.200 327.600 223.200 328.200 ;
        RECT 114.600 327.000 118.200 327.600 ;
        RECT 177.000 327.000 183.600 327.600 ;
        RECT 216.600 327.000 224.400 327.600 ;
        RECT 228.000 327.000 231.600 328.800 ;
        RECT 262.800 328.200 266.400 328.800 ;
        RECT 263.400 327.600 267.000 328.200 ;
        RECT 114.000 326.400 117.600 327.000 ;
        RECT 178.200 326.400 180.600 327.000 ;
        RECT 218.400 326.400 225.600 327.000 ;
        RECT 226.800 326.400 231.600 327.000 ;
        RECT 264.000 326.400 267.600 327.600 ;
        RECT 274.200 327.000 277.200 328.800 ;
        RECT 273.600 326.400 277.200 327.000 ;
        RECT 287.400 326.400 290.400 330.000 ;
        RECT 478.800 329.400 482.400 330.000 ;
        RECT 517.200 329.400 520.800 330.000 ;
        RECT 479.400 327.600 482.400 329.400 ;
        RECT 517.800 328.800 520.800 329.400 ;
        RECT 578.400 329.400 581.400 330.600 ;
        RECT 688.200 330.000 691.800 331.200 ;
        RECT 675.000 329.400 687.000 330.000 ;
        RECT 688.200 329.400 692.400 330.000 ;
        RECT 578.400 328.800 582.000 329.400 ;
        RECT 670.800 328.800 692.400 329.400 ;
        RECT 517.800 328.200 521.400 328.800 ;
        RECT 518.400 327.600 521.400 328.200 ;
        RECT 579.000 327.600 582.000 328.800 ;
        RECT 669.600 328.200 692.400 328.800 ;
        RECT 669.000 327.600 693.000 328.200 ;
        RECT 479.400 327.000 483.000 327.600 ;
        RECT 518.400 327.000 522.000 327.600 ;
        RECT 579.000 327.000 582.600 327.600 ;
        RECT 113.400 325.800 117.600 326.400 ;
        RECT 219.600 325.800 231.000 326.400 ;
        RECT 264.600 325.800 268.200 326.400 ;
        RECT 113.400 325.200 117.000 325.800 ;
        RECT 221.400 325.200 230.400 325.800 ;
        RECT 265.200 325.200 268.200 325.800 ;
        RECT 112.800 324.600 116.400 325.200 ;
        RECT 222.600 324.600 229.800 325.200 ;
        RECT 265.200 324.600 268.800 325.200 ;
        RECT 273.600 324.600 276.600 326.400 ;
        RECT 112.200 323.400 115.800 324.600 ;
        RECT 223.800 324.000 229.800 324.600 ;
        RECT 265.800 324.000 269.400 324.600 ;
        RECT 225.000 323.400 229.800 324.000 ;
        RECT 266.400 323.400 269.400 324.000 ;
        RECT 111.600 322.800 115.200 323.400 ;
        RECT 225.600 322.800 230.400 323.400 ;
        RECT 266.400 322.800 270.000 323.400 ;
        RECT 111.600 322.200 114.600 322.800 ;
        RECT 226.800 322.200 231.600 322.800 ;
        RECT 267.000 322.200 270.000 322.800 ;
        RECT 273.000 322.200 276.000 324.600 ;
        RECT 111.000 321.600 114.600 322.200 ;
        RECT 227.400 321.600 232.200 322.200 ;
        RECT 267.000 321.600 270.600 322.200 ;
        RECT 111.000 321.000 114.000 321.600 ;
        RECT 228.000 321.000 232.800 321.600 ;
        RECT 267.600 321.000 270.600 321.600 ;
        RECT 110.400 319.800 113.400 321.000 ;
        RECT 153.600 320.400 156.600 321.000 ;
        RECT 229.200 320.400 233.400 321.000 ;
        RECT 267.600 320.400 271.200 321.000 ;
        RECT 152.400 319.800 159.000 320.400 ;
        RECT 229.800 319.800 234.000 320.400 ;
        RECT 109.800 318.600 112.800 319.800 ;
        RECT 151.800 319.200 161.400 319.800 ;
        RECT 230.400 319.200 234.600 319.800 ;
        RECT 268.200 319.200 271.200 320.400 ;
        RECT 272.400 319.200 275.400 322.200 ;
        RECT 288.000 321.600 291.000 326.400 ;
        RECT 303.600 325.800 306.000 326.400 ;
        RECT 302.400 325.200 307.200 325.800 ;
        RECT 480.000 325.200 483.000 327.000 ;
        RECT 519.000 325.800 522.000 327.000 ;
        RECT 579.600 325.800 582.600 327.000 ;
        RECT 668.400 327.000 693.000 327.600 ;
        RECT 668.400 325.800 678.600 327.000 ;
        RECT 684.000 326.400 693.000 327.000 ;
        RECT 687.000 325.800 693.000 326.400 ;
        RECT 301.800 324.600 307.800 325.200 ;
        RECT 480.000 324.600 483.600 325.200 ;
        RECT 301.200 323.400 308.400 324.600 ;
        RECT 480.600 323.400 483.600 324.600 ;
        RECT 519.600 324.600 522.600 325.800 ;
        RECT 579.600 325.200 583.200 325.800 ;
        RECT 669.600 325.200 681.000 325.800 ;
        RECT 688.800 325.200 693.000 325.800 ;
        RECT 519.600 324.000 523.200 324.600 ;
        RECT 580.200 324.000 583.200 325.200 ;
        RECT 671.400 324.600 682.800 325.200 ;
        RECT 690.600 324.600 692.400 325.200 ;
        RECT 673.800 324.000 684.600 324.600 ;
        RECT 520.200 323.400 523.200 324.000 ;
        RECT 300.600 322.800 304.200 323.400 ;
        RECT 305.400 322.800 309.000 323.400 ;
        RECT 300.000 322.200 303.600 322.800 ;
        RECT 306.000 322.200 309.600 322.800 ;
        RECT 480.600 322.200 484.200 323.400 ;
        RECT 520.200 322.800 523.800 323.400 ;
        RECT 154.800 318.600 162.600 319.200 ;
        RECT 231.000 318.600 235.200 319.200 ;
        RECT 109.200 318.000 112.800 318.600 ;
        RECT 156.600 318.000 164.400 318.600 ;
        RECT 231.600 318.000 235.200 318.600 ;
        RECT 268.800 318.600 275.400 319.200 ;
        RECT 109.200 316.800 112.200 318.000 ;
        RECT 158.400 317.400 166.200 318.000 ;
        RECT 232.200 317.400 235.800 318.000 ;
        RECT 268.800 317.400 274.800 318.600 ;
        RECT 160.200 316.800 167.400 317.400 ;
        RECT 232.800 316.800 236.400 317.400 ;
        RECT 108.600 315.000 111.600 316.800 ;
        RECT 161.400 316.200 168.600 316.800 ;
        RECT 163.200 315.600 170.400 316.200 ;
        RECT 233.400 315.600 237.000 316.800 ;
        RECT 269.400 315.600 274.800 317.400 ;
        RECT 164.400 315.000 171.600 315.600 ;
        RECT 234.000 315.000 237.600 315.600 ;
        RECT 108.600 313.800 111.000 315.000 ;
        RECT 165.600 314.400 172.800 315.000 ;
        RECT 234.600 314.400 237.600 315.000 ;
        RECT 270.000 314.400 274.200 315.600 ;
        RECT 288.600 315.000 291.600 321.600 ;
        RECT 299.400 321.000 303.000 322.200 ;
        RECT 306.600 321.000 309.600 322.200 ;
        RECT 481.200 321.600 484.200 322.200 ;
        RECT 520.800 322.200 523.800 322.800 ;
        RECT 580.800 322.800 583.800 324.000 ;
        RECT 676.200 323.400 685.800 324.000 ;
        RECT 678.600 322.800 687.000 323.400 ;
        RECT 580.800 322.200 584.400 322.800 ;
        RECT 681.000 322.200 688.200 322.800 ;
        RECT 520.800 321.600 524.400 322.200 ;
        RECT 298.800 320.400 302.400 321.000 ;
        RECT 306.600 320.400 310.200 321.000 ;
        RECT 481.200 320.400 484.800 321.600 ;
        RECT 521.400 321.000 524.400 321.600 ;
        RECT 581.400 321.600 584.400 322.200 ;
        RECT 682.800 321.600 688.800 322.200 ;
        RECT 521.400 320.400 525.000 321.000 ;
        RECT 581.400 320.400 585.000 321.600 ;
        RECT 684.000 321.000 690.000 321.600 ;
        RECT 685.200 320.400 690.600 321.000 ;
        RECT 298.800 319.800 301.800 320.400 ;
        RECT 298.200 319.200 301.800 319.800 ;
        RECT 307.200 319.200 310.200 320.400 ;
        RECT 481.800 319.200 484.800 320.400 ;
        RECT 522.000 319.800 525.000 320.400 ;
        RECT 582.000 319.800 585.000 320.400 ;
        RECT 686.400 319.800 691.200 320.400 ;
        RECT 522.000 319.200 525.600 319.800 ;
        RECT 582.000 319.200 585.600 319.800 ;
        RECT 687.600 319.200 691.800 319.800 ;
        RECT 297.600 318.000 301.200 319.200 ;
        RECT 297.000 317.400 300.600 318.000 ;
        RECT 297.000 316.800 300.000 317.400 ;
        RECT 307.800 316.800 310.800 319.200 ;
        RECT 481.800 318.600 485.400 319.200 ;
        RECT 522.600 318.600 525.600 319.200 ;
        RECT 582.600 318.600 585.600 319.200 ;
        RECT 688.200 318.600 691.800 319.200 ;
        RECT 482.400 317.400 485.400 318.600 ;
        RECT 523.200 318.000 526.200 318.600 ;
        RECT 523.200 317.400 526.800 318.000 ;
        RECT 582.600 317.400 586.200 318.600 ;
        RECT 622.200 317.400 623.400 318.000 ;
        RECT 688.800 317.400 691.800 318.600 ;
        RECT 482.400 316.800 486.000 317.400 ;
        RECT 296.400 316.200 300.000 316.800 ;
        RECT 296.400 315.600 299.400 316.200 ;
        RECT 166.800 313.800 174.000 314.400 ;
        RECT 234.600 313.800 238.200 314.400 ;
        RECT 270.000 313.800 273.600 314.400 ;
        RECT 108.000 312.000 111.000 313.800 ;
        RECT 168.600 313.200 175.200 313.800 ;
        RECT 235.200 313.200 238.200 313.800 ;
        RECT 169.800 312.600 176.400 313.200 ;
        RECT 171.000 312.000 177.600 312.600 ;
        RECT 235.800 312.000 238.800 313.200 ;
        RECT 108.600 310.800 111.000 312.000 ;
        RECT 172.200 311.400 178.800 312.000 ;
        RECT 235.800 311.400 239.400 312.000 ;
        RECT 173.400 310.800 180.000 311.400 ;
        RECT 236.400 310.800 239.400 311.400 ;
        RECT 108.600 307.200 111.600 310.800 ;
        RECT 174.600 310.200 181.200 310.800 ;
        RECT 236.400 310.200 240.000 310.800 ;
        RECT 270.600 310.200 273.600 313.800 ;
        RECT 175.800 309.600 182.400 310.200 ;
        RECT 177.000 309.000 183.600 309.600 ;
        RECT 237.000 309.000 240.000 310.200 ;
        RECT 271.200 309.600 273.600 310.200 ;
        RECT 289.200 313.800 291.600 315.000 ;
        RECT 295.800 315.000 299.400 315.600 ;
        RECT 295.800 314.400 298.800 315.000 ;
        RECT 295.200 313.800 298.800 314.400 ;
        RECT 308.400 313.800 311.400 316.800 ;
        RECT 483.000 315.000 486.000 316.800 ;
        RECT 523.800 316.800 526.800 317.400 ;
        RECT 583.200 316.800 586.200 317.400 ;
        RECT 613.800 316.800 624.600 317.400 ;
        RECT 523.800 316.200 527.400 316.800 ;
        RECT 583.200 316.200 586.800 316.800 ;
        RECT 610.200 316.200 624.600 316.800 ;
        RECT 524.400 315.600 527.400 316.200 ;
        RECT 524.400 315.000 528.000 315.600 ;
        RECT 583.800 315.000 586.800 316.200 ;
        RECT 606.600 315.600 624.600 316.200 ;
        RECT 603.600 315.000 624.600 315.600 ;
        RECT 289.200 309.600 292.200 313.800 ;
        RECT 295.200 313.200 298.200 313.800 ;
        RECT 294.600 312.600 298.200 313.200 ;
        RECT 309.000 313.200 311.400 313.800 ;
        RECT 483.600 313.200 486.600 315.000 ;
        RECT 525.000 313.800 528.600 315.000 ;
        RECT 584.400 313.800 587.400 315.000 ;
        RECT 601.200 314.400 623.400 315.000 ;
        RECT 689.400 314.400 692.400 317.400 ;
        RECT 598.800 313.800 621.600 314.400 ;
        RECT 525.600 313.200 529.200 313.800 ;
        RECT 584.400 313.200 588.000 313.800 ;
        RECT 597.000 313.200 609.600 313.800 ;
        RECT 613.200 313.200 620.400 313.800 ;
        RECT 294.600 312.000 297.600 312.600 ;
        RECT 294.000 311.400 297.600 312.000 ;
        RECT 294.000 310.800 297.000 311.400 ;
        RECT 293.400 310.200 297.000 310.800 ;
        RECT 293.400 309.600 296.400 310.200 ;
        RECT 178.200 308.400 184.800 309.000 ;
        RECT 237.000 308.400 240.600 309.000 ;
        RECT 179.400 307.800 185.400 308.400 ;
        RECT 180.600 307.200 186.600 307.800 ;
        RECT 109.200 304.800 112.200 307.200 ;
        RECT 181.800 306.600 187.800 307.200 ;
        RECT 237.600 306.600 240.600 308.400 ;
        RECT 183.000 306.000 189.000 306.600 ;
        RECT 184.200 305.400 189.600 306.000 ;
        RECT 184.800 304.800 190.800 305.400 ;
        RECT 109.800 303.000 112.800 304.800 ;
        RECT 186.000 304.200 191.400 304.800 ;
        RECT 238.200 304.200 241.200 306.600 ;
        RECT 271.200 304.800 274.200 309.600 ;
        RECT 289.200 309.000 296.400 309.600 ;
        RECT 289.200 307.800 295.800 309.000 ;
        RECT 289.200 306.600 295.200 307.800 ;
        RECT 289.200 305.400 294.600 306.600 ;
        RECT 271.200 304.200 273.600 304.800 ;
        RECT 187.200 303.600 192.600 304.200 ;
        RECT 187.800 303.000 193.800 303.600 ;
        RECT 110.400 301.800 113.400 303.000 ;
        RECT 189.000 302.400 194.400 303.000 ;
        RECT 190.200 301.800 195.600 302.400 ;
        RECT 110.400 301.200 114.000 301.800 ;
        RECT 190.800 301.200 196.200 301.800 ;
        RECT 111.000 300.600 114.000 301.200 ;
        RECT 192.000 300.600 196.800 301.200 ;
        RECT 238.800 300.600 241.800 304.200 ;
        RECT 270.600 301.200 273.600 304.200 ;
        RECT 289.200 304.200 294.000 305.400 ;
        RECT 289.200 303.000 293.400 304.200 ;
        RECT 289.200 301.800 292.800 303.000 ;
        RECT 111.000 299.400 114.600 300.600 ;
        RECT 192.600 300.000 198.000 300.600 ;
        RECT 239.400 300.000 241.800 300.600 ;
        RECT 193.800 299.400 198.600 300.000 ;
        RECT 111.600 298.200 115.200 299.400 ;
        RECT 194.400 298.800 199.200 299.400 ;
        RECT 195.600 298.200 200.400 298.800 ;
        RECT 112.200 297.600 115.800 298.200 ;
        RECT 196.200 297.600 201.000 298.200 ;
        RECT 112.800 297.000 116.400 297.600 ;
        RECT 196.800 297.000 201.600 297.600 ;
        RECT 112.800 296.400 117.000 297.000 ;
        RECT 198.000 296.400 202.800 297.000 ;
        RECT 113.400 295.200 117.600 296.400 ;
        RECT 198.600 295.800 203.400 296.400 ;
        RECT 199.200 295.200 205.200 295.800 ;
        RECT 105.000 294.600 118.800 295.200 ;
        RECT 200.400 294.600 206.400 295.200 ;
        RECT 100.800 294.000 123.000 294.600 ;
        RECT 201.000 294.000 207.600 294.600 ;
        RECT 99.000 293.400 126.000 294.000 ;
        RECT 201.600 293.400 208.800 294.000 ;
        RECT 97.200 292.800 129.000 293.400 ;
        RECT 202.200 292.800 210.000 293.400 ;
        RECT 96.600 292.200 131.400 292.800 ;
        RECT 202.800 292.200 210.600 292.800 ;
        RECT 96.000 291.600 104.400 292.200 ;
        RECT 119.400 291.600 133.200 292.200 ;
        RECT 203.400 291.600 211.800 292.200 ;
        RECT 95.400 291.000 100.800 291.600 ;
        RECT 123.600 291.000 134.400 291.600 ;
        RECT 204.000 291.000 213.000 291.600 ;
        RECT 95.400 290.400 99.000 291.000 ;
        RECT 126.600 290.400 135.600 291.000 ;
        RECT 204.600 290.400 214.200 291.000 ;
        RECT 95.400 289.200 98.400 290.400 ;
        RECT 129.000 289.800 136.200 290.400 ;
        RECT 205.200 289.800 214.800 290.400 ;
        RECT 239.400 289.800 242.400 300.000 ;
        RECT 270.000 299.400 273.000 301.200 ;
        RECT 289.200 300.600 292.200 301.800 ;
        RECT 288.600 299.400 291.600 300.600 ;
        RECT 269.400 298.200 272.400 299.400 ;
        RECT 288.000 298.200 291.000 299.400 ;
        RECT 268.800 297.600 272.400 298.200 ;
        RECT 287.400 297.600 291.000 298.200 ;
        RECT 268.800 297.000 273.000 297.600 ;
        RECT 287.400 297.000 290.400 297.600 ;
        RECT 309.000 297.000 312.000 313.200 ;
        RECT 484.200 312.000 487.200 313.200 ;
        RECT 526.200 312.600 529.200 313.200 ;
        RECT 526.200 312.000 529.800 312.600 ;
        RECT 484.200 311.400 487.800 312.000 ;
        RECT 484.800 310.200 487.800 311.400 ;
        RECT 526.800 311.400 529.800 312.000 ;
        RECT 585.000 312.000 588.000 313.200 ;
        RECT 595.200 312.600 606.600 313.200 ;
        RECT 613.200 312.600 619.200 313.200 ;
        RECT 593.400 312.000 603.600 312.600 ;
        RECT 612.000 312.000 618.000 312.600 ;
        RECT 585.000 311.400 588.600 312.000 ;
        RECT 591.600 311.400 601.200 312.000 ;
        RECT 611.400 311.400 616.800 312.000 ;
        RECT 690.000 311.400 693.000 314.400 ;
        RECT 526.800 310.800 530.400 311.400 ;
        RECT 527.400 310.200 530.400 310.800 ;
        RECT 585.600 310.800 588.600 311.400 ;
        RECT 590.400 310.800 598.800 311.400 ;
        RECT 610.200 310.800 616.200 311.400 ;
        RECT 585.600 310.200 597.000 310.800 ;
        RECT 609.000 310.200 615.000 310.800 ;
        RECT 484.800 309.600 488.400 310.200 ;
        RECT 527.400 309.600 531.000 310.200 ;
        RECT 586.200 309.600 595.200 310.200 ;
        RECT 608.400 309.600 613.800 310.200 ;
        RECT 485.400 309.000 488.400 309.600 ;
        RECT 528.000 309.000 531.600 309.600 ;
        RECT 586.200 309.000 593.400 309.600 ;
        RECT 607.200 309.000 612.600 309.600 ;
        RECT 485.400 308.400 489.000 309.000 ;
        RECT 486.000 307.200 489.000 308.400 ;
        RECT 528.600 308.400 531.600 309.000 ;
        RECT 586.800 308.400 592.200 309.000 ;
        RECT 606.600 308.400 612.000 309.000 ;
        RECT 690.600 308.400 693.600 311.400 ;
        RECT 528.600 307.800 532.200 308.400 ;
        RECT 587.400 307.800 590.400 308.400 ;
        RECT 605.400 307.800 610.800 308.400 ;
        RECT 691.200 307.800 693.600 308.400 ;
        RECT 486.600 306.000 489.600 307.200 ;
        RECT 529.200 306.600 532.800 307.800 ;
        RECT 604.200 307.200 610.200 307.800 ;
        RECT 603.600 306.600 609.000 307.200 ;
        RECT 529.800 306.000 533.400 306.600 ;
        RECT 602.400 306.000 607.800 306.600 ;
        RECT 486.600 305.400 490.200 306.000 ;
        RECT 487.200 304.800 490.200 305.400 ;
        RECT 530.400 305.400 533.400 306.000 ;
        RECT 601.800 305.400 607.200 306.000 ;
        RECT 530.400 304.800 534.000 305.400 ;
        RECT 600.600 304.800 606.000 305.400 ;
        RECT 487.200 304.200 490.800 304.800 ;
        RECT 487.800 303.600 490.800 304.200 ;
        RECT 531.000 303.600 534.600 304.800 ;
        RECT 600.000 304.200 605.400 304.800 ;
        RECT 691.200 304.200 694.200 307.800 ;
        RECT 598.800 303.600 604.200 304.200 ;
        RECT 691.800 303.600 694.200 304.200 ;
        RECT 487.800 303.000 491.400 303.600 ;
        RECT 531.600 303.000 535.200 303.600 ;
        RECT 597.600 303.000 603.000 303.600 ;
        RECT 488.400 301.800 491.400 303.000 ;
        RECT 532.200 301.800 535.800 303.000 ;
        RECT 597.000 302.400 602.400 303.000 ;
        RECT 595.800 301.800 601.200 302.400 ;
        RECT 489.000 300.600 492.000 301.800 ;
        RECT 532.800 301.200 536.400 301.800 ;
        RECT 595.200 301.200 600.600 301.800 ;
        RECT 533.400 300.600 536.400 301.200 ;
        RECT 594.000 300.600 599.400 301.200 ;
        RECT 489.000 300.000 492.600 300.600 ;
        RECT 533.400 300.000 537.000 300.600 ;
        RECT 592.800 300.000 598.800 300.600 ;
        RECT 489.600 299.400 492.600 300.000 ;
        RECT 534.000 299.400 537.600 300.000 ;
        RECT 592.200 299.400 597.600 300.000 ;
        RECT 489.600 298.800 493.200 299.400 ;
        RECT 490.200 298.200 493.200 298.800 ;
        RECT 534.600 298.800 537.600 299.400 ;
        RECT 591.000 298.800 596.400 299.400 ;
        RECT 534.600 298.200 538.200 298.800 ;
        RECT 590.400 298.200 595.800 298.800 ;
        RECT 691.800 298.200 694.800 303.600 ;
        RECT 490.200 297.600 493.800 298.200 ;
        RECT 490.800 297.000 493.800 297.600 ;
        RECT 535.200 297.000 538.800 298.200 ;
        RECT 589.200 297.600 594.600 298.200 ;
        RECT 692.400 297.600 694.800 298.200 ;
        RECT 588.600 297.000 594.000 297.600 ;
        RECT 268.200 296.400 273.000 297.000 ;
        RECT 286.800 296.400 290.400 297.000 ;
        RECT 268.200 295.800 273.600 296.400 ;
        RECT 267.600 294.600 274.200 295.800 ;
        RECT 286.800 295.200 289.800 296.400 ;
        RECT 267.000 294.000 274.800 294.600 ;
        RECT 286.200 294.000 289.200 295.200 ;
        RECT 266.400 293.400 270.000 294.000 ;
        RECT 265.800 292.800 270.000 293.400 ;
        RECT 271.800 292.800 274.800 294.000 ;
        RECT 285.600 293.400 289.200 294.000 ;
        RECT 265.200 292.200 269.400 292.800 ;
        RECT 264.600 291.600 268.800 292.200 ;
        RECT 272.400 291.600 275.400 292.800 ;
        RECT 285.600 292.200 288.600 293.400 ;
        RECT 308.400 292.200 311.400 297.000 ;
        RECT 490.800 296.400 494.400 297.000 ;
        RECT 535.800 296.400 539.400 297.000 ;
        RECT 587.400 296.400 592.800 297.000 ;
        RECT 491.400 295.800 494.400 296.400 ;
        RECT 491.400 295.200 495.000 295.800 ;
        RECT 536.400 295.200 540.000 296.400 ;
        RECT 586.800 295.800 591.600 296.400 ;
        RECT 585.600 295.200 591.000 295.800 ;
        RECT 492.000 294.600 495.000 295.200 ;
        RECT 537.000 294.600 540.600 295.200 ;
        RECT 585.000 294.600 589.800 295.200 ;
        RECT 492.000 294.000 495.600 294.600 ;
        RECT 492.600 293.400 496.200 294.000 ;
        RECT 537.600 293.400 541.200 294.600 ;
        RECT 585.000 293.400 589.200 294.600 ;
        RECT 493.200 292.800 496.200 293.400 ;
        RECT 538.200 292.800 541.800 293.400 ;
        RECT 585.000 292.800 589.800 293.400 ;
        RECT 493.200 292.200 496.800 292.800 ;
        RECT 264.000 291.000 268.200 291.600 ;
        RECT 272.400 291.000 276.000 291.600 ;
        RECT 285.000 291.000 288.000 292.200 ;
        RECT 263.400 290.400 267.600 291.000 ;
        RECT 262.800 289.800 267.600 290.400 ;
        RECT 273.000 289.800 276.000 291.000 ;
        RECT 284.400 290.400 288.000 291.000 ;
        RECT 130.800 289.200 136.800 289.800 ;
        RECT 205.800 289.200 216.000 289.800 ;
        RECT 239.400 289.200 241.800 289.800 ;
        RECT 261.600 289.200 267.000 289.800 ;
        RECT 95.400 288.600 99.000 289.200 ;
        RECT 133.200 288.600 136.800 289.200 ;
        RECT 206.400 288.600 217.200 289.200 ;
        RECT 96.000 287.400 99.600 288.600 ;
        RECT 135.000 288.000 136.200 288.600 ;
        RECT 207.000 288.000 211.200 288.600 ;
        RECT 212.400 288.000 218.400 288.600 ;
        RECT 207.600 287.400 211.200 288.000 ;
        RECT 213.600 287.400 219.000 288.000 ;
        RECT 96.600 286.800 100.800 287.400 ;
        RECT 208.200 286.800 211.800 287.400 ;
        RECT 214.200 286.800 220.200 287.400 ;
        RECT 97.200 286.200 101.400 286.800 ;
        RECT 208.800 286.200 212.400 286.800 ;
        RECT 215.400 286.200 221.400 286.800 ;
        RECT 238.800 286.200 241.800 289.200 ;
        RECT 261.000 288.600 266.400 289.200 ;
        RECT 273.600 288.600 276.600 289.800 ;
        RECT 284.400 289.200 287.400 290.400 ;
        RECT 260.400 288.000 265.800 288.600 ;
        RECT 273.600 288.000 277.200 288.600 ;
        RECT 283.800 288.000 286.800 289.200 ;
        RECT 307.800 288.600 310.800 292.200 ;
        RECT 493.800 291.600 496.800 292.200 ;
        RECT 538.800 291.600 542.400 292.800 ;
        RECT 585.600 292.200 590.400 292.800 ;
        RECT 586.200 291.600 591.000 292.200 ;
        RECT 493.800 291.000 497.400 291.600 ;
        RECT 539.400 291.000 543.000 291.600 ;
        RECT 587.400 291.000 591.600 291.600 ;
        RECT 494.400 290.400 497.400 291.000 ;
        RECT 494.400 289.800 498.000 290.400 ;
        RECT 540.000 289.800 543.600 291.000 ;
        RECT 588.000 290.400 592.200 291.000 ;
        RECT 588.600 289.800 592.800 290.400 ;
        RECT 495.000 289.200 498.000 289.800 ;
        RECT 540.600 289.200 544.200 289.800 ;
        RECT 589.200 289.200 593.400 289.800 ;
        RECT 495.000 288.600 498.600 289.200 ;
        RECT 259.800 287.400 265.200 288.000 ;
        RECT 259.200 286.800 264.000 287.400 ;
        RECT 274.200 286.800 277.200 288.000 ;
        RECT 283.200 287.400 286.800 288.000 ;
        RECT 258.000 286.200 263.400 286.800 ;
        RECT 274.200 286.200 277.800 286.800 ;
        RECT 283.200 286.200 286.200 287.400 ;
        RECT 97.800 285.600 102.000 286.200 ;
        RECT 209.400 285.600 212.400 286.200 ;
        RECT 216.600 285.600 222.600 286.200 ;
        RECT 98.400 285.000 102.600 285.600 ;
        RECT 99.000 284.400 103.800 285.000 ;
        RECT 210.000 284.400 213.000 285.600 ;
        RECT 217.800 285.000 223.200 285.600 ;
        RECT 238.200 285.000 241.200 286.200 ;
        RECT 257.400 285.600 262.800 286.200 ;
        RECT 256.200 285.000 262.200 285.600 ;
        RECT 274.800 285.000 277.800 286.200 ;
        RECT 218.400 284.400 224.400 285.000 ;
        RECT 99.600 283.800 104.400 284.400 ;
        RECT 210.600 283.800 213.600 284.400 ;
        RECT 219.600 283.800 225.600 284.400 ;
        RECT 237.600 283.800 241.200 285.000 ;
        RECT 255.000 284.400 261.000 285.000 ;
        RECT 274.800 284.400 278.400 285.000 ;
        RECT 282.600 284.400 285.600 286.200 ;
        RECT 307.200 285.600 310.200 288.600 ;
        RECT 495.600 288.000 499.200 288.600 ;
        RECT 541.200 288.000 544.800 289.200 ;
        RECT 589.800 288.600 594.000 289.200 ;
        RECT 590.400 288.000 594.600 288.600 ;
        RECT 496.200 287.400 499.200 288.000 ;
        RECT 541.800 287.400 545.400 288.000 ;
        RECT 591.000 287.400 595.200 288.000 ;
        RECT 496.200 286.800 499.800 287.400 ;
        RECT 496.800 286.200 499.800 286.800 ;
        RECT 542.400 286.200 546.000 287.400 ;
        RECT 591.600 286.800 595.800 287.400 ;
        RECT 592.200 286.200 596.400 286.800 ;
        RECT 496.800 285.600 500.400 286.200 ;
        RECT 543.000 285.600 546.600 286.200 ;
        RECT 592.800 285.600 597.600 286.200 ;
        RECT 253.800 283.800 260.400 284.400 ;
        RECT 100.200 283.200 105.600 283.800 ;
        RECT 211.200 283.200 213.600 283.800 ;
        RECT 220.800 283.200 226.200 283.800 ;
        RECT 237.600 283.200 240.600 283.800 ;
        RECT 252.600 283.200 259.200 283.800 ;
        RECT 100.800 282.600 106.200 283.200 ;
        RECT 211.800 282.600 214.200 283.200 ;
        RECT 221.400 282.600 227.400 283.200 ;
        RECT 237.000 282.600 240.600 283.200 ;
        RECT 251.400 282.600 258.000 283.200 ;
        RECT 275.400 282.600 278.400 284.400 ;
        RECT 282.000 283.200 285.000 284.400 ;
        RECT 306.600 283.200 309.600 285.600 ;
        RECT 497.400 285.000 501.000 285.600 ;
        RECT 543.600 285.000 547.200 285.600 ;
        RECT 593.400 285.000 598.200 285.600 ;
        RECT 498.000 284.400 501.000 285.000 ;
        RECT 544.200 284.400 547.200 285.000 ;
        RECT 594.600 284.400 598.800 285.000 ;
        RECT 498.000 283.800 501.600 284.400 ;
        RECT 544.200 283.800 547.800 284.400 ;
        RECT 595.200 283.800 599.400 284.400 ;
        RECT 498.600 283.200 501.600 283.800 ;
        RECT 544.800 283.200 548.400 283.800 ;
        RECT 595.800 283.200 600.000 283.800 ;
        RECT 281.400 282.600 285.000 283.200 ;
        RECT 102.000 282.000 107.400 282.600 ;
        RECT 212.400 282.000 214.200 282.600 ;
        RECT 222.600 282.000 228.000 282.600 ;
        RECT 237.000 282.000 240.000 282.600 ;
        RECT 250.200 282.000 256.800 282.600 ;
        RECT 102.600 281.400 108.600 282.000 ;
        RECT 103.800 280.800 109.200 281.400 ;
        RECT 213.000 280.800 214.800 282.000 ;
        RECT 223.800 281.400 229.200 282.000 ;
        RECT 224.400 280.800 230.400 281.400 ;
        RECT 236.400 280.800 240.000 282.000 ;
        RECT 248.400 281.400 255.600 282.000 ;
        RECT 247.200 280.800 255.000 281.400 ;
        RECT 104.400 280.200 110.400 280.800 ;
        RECT 213.600 280.200 214.800 280.800 ;
        RECT 225.600 280.200 231.000 280.800 ;
        RECT 236.400 280.200 239.400 280.800 ;
        RECT 105.600 279.600 112.200 280.200 ;
        RECT 214.200 279.600 215.400 280.200 ;
        RECT 226.800 279.600 232.200 280.200 ;
        RECT 235.800 279.600 239.400 280.200 ;
        RECT 246.000 280.200 253.800 280.800 ;
        RECT 276.000 280.200 279.000 282.600 ;
        RECT 281.400 281.400 284.400 282.600 ;
        RECT 246.000 279.600 252.600 280.200 ;
        RECT 276.600 279.600 279.600 280.200 ;
        RECT 280.800 279.600 283.800 281.400 ;
        RECT 306.000 280.800 309.000 283.200 ;
        RECT 498.600 282.600 502.200 283.200 ;
        RECT 499.200 282.000 502.800 282.600 ;
        RECT 545.400 282.000 549.000 283.200 ;
        RECT 596.400 282.600 600.600 283.200 ;
        RECT 597.000 282.000 601.200 282.600 ;
        RECT 692.400 282.000 695.400 297.600 ;
        RECT 499.800 281.400 502.800 282.000 ;
        RECT 546.000 281.400 549.600 282.000 ;
        RECT 597.600 281.400 601.800 282.000 ;
        RECT 499.800 280.800 503.400 281.400 ;
        RECT 106.800 279.000 113.400 279.600 ;
        RECT 214.800 279.000 215.400 279.600 ;
        RECT 227.400 279.000 232.800 279.600 ;
        RECT 235.800 279.000 238.800 279.600 ;
        RECT 246.000 279.000 250.800 279.600 ;
        RECT 108.000 278.400 114.600 279.000 ;
        RECT 228.600 278.400 234.000 279.000 ;
        RECT 235.200 278.400 238.800 279.000 ;
        RECT 246.600 278.400 249.600 279.000 ;
        RECT 109.200 277.800 116.400 278.400 ;
        RECT 229.200 277.800 238.200 278.400 ;
        RECT 110.400 277.200 118.200 277.800 ;
        RECT 230.400 277.200 238.200 277.800 ;
        RECT 247.200 277.800 249.600 278.400 ;
        RECT 276.600 277.800 283.200 279.600 ;
        RECT 305.400 278.400 308.400 280.800 ;
        RECT 500.400 280.200 503.400 280.800 ;
        RECT 546.600 280.200 550.200 281.400 ;
        RECT 598.200 280.800 602.400 281.400 ;
        RECT 692.400 280.800 694.800 282.000 ;
        RECT 598.800 280.200 603.000 280.800 ;
        RECT 500.400 279.600 504.000 280.200 ;
        RECT 547.200 279.600 550.800 280.200 ;
        RECT 599.400 279.600 603.600 280.200 ;
        RECT 501.000 279.000 504.600 279.600 ;
        RECT 547.800 279.000 551.400 279.600 ;
        RECT 600.000 279.000 604.200 279.600 ;
        RECT 501.600 278.400 504.600 279.000 ;
        RECT 247.200 277.200 250.200 277.800 ;
        RECT 111.600 276.600 119.400 277.200 ;
        RECT 231.000 276.600 238.200 277.200 ;
        RECT 112.800 276.000 121.800 276.600 ;
        RECT 232.200 276.000 238.200 276.600 ;
        RECT 114.600 275.400 123.600 276.000 ;
        RECT 232.800 275.400 238.200 276.000 ;
        RECT 247.800 276.600 250.200 277.200 ;
        RECT 247.800 275.400 250.800 276.600 ;
        RECT 277.200 276.000 282.600 277.800 ;
        RECT 304.800 276.000 307.800 278.400 ;
        RECT 501.600 277.800 505.200 278.400 ;
        RECT 548.400 277.800 552.000 279.000 ;
        RECT 600.600 278.400 605.400 279.000 ;
        RECT 601.200 277.800 606.000 278.400 ;
        RECT 502.200 277.200 505.800 277.800 ;
        RECT 549.000 277.200 552.600 277.800 ;
        RECT 601.800 277.200 606.600 277.800 ;
        RECT 502.200 276.600 506.400 277.200 ;
        RECT 502.800 276.000 506.400 276.600 ;
        RECT 549.600 276.000 553.200 277.200 ;
        RECT 603.000 276.600 607.200 277.200 ;
        RECT 603.600 276.000 607.800 276.600 ;
        RECT 277.200 275.400 282.000 276.000 ;
        RECT 115.800 274.800 126.000 275.400 ;
        RECT 234.000 274.800 239.400 275.400 ;
        RECT 117.600 274.200 128.400 274.800 ;
        RECT 234.600 274.200 240.000 274.800 ;
        RECT 248.400 274.200 251.400 275.400 ;
        RECT 277.800 274.800 282.000 275.400 ;
        RECT 119.400 273.600 130.800 274.200 ;
        RECT 235.800 273.600 240.600 274.200 ;
        RECT 248.400 273.600 252.000 274.200 ;
        RECT 121.200 273.000 133.200 273.600 ;
        RECT 236.400 273.000 241.800 273.600 ;
        RECT 122.400 272.400 135.600 273.000 ;
        RECT 237.600 272.400 242.400 273.000 ;
        RECT 249.000 272.400 252.000 273.600 ;
        RECT 277.800 273.000 281.400 274.800 ;
        RECT 304.200 274.200 307.200 276.000 ;
        RECT 503.400 274.800 507.000 276.000 ;
        RECT 550.200 275.400 553.800 276.000 ;
        RECT 604.200 275.400 608.400 276.000 ;
        RECT 550.800 274.800 554.400 275.400 ;
        RECT 604.800 274.800 609.000 275.400 ;
        RECT 691.800 274.800 694.800 280.800 ;
        RECT 504.000 274.200 507.600 274.800 ;
        RECT 124.800 271.800 138.600 272.400 ;
        RECT 238.200 271.800 243.000 272.400 ;
        RECT 126.600 271.200 141.000 271.800 ;
        RECT 239.400 271.200 244.200 271.800 ;
        RECT 249.600 271.200 252.600 272.400 ;
        RECT 126.600 270.600 154.200 271.200 ;
        RECT 240.000 270.600 244.800 271.200 ;
        RECT 114.000 270.000 159.600 270.600 ;
        RECT 240.600 270.000 246.000 270.600 ;
        RECT 250.200 270.000 253.200 271.200 ;
        RECT 278.400 270.000 281.400 273.000 ;
        RECT 303.600 273.600 307.200 274.200 ;
        RECT 303.600 271.800 306.600 273.600 ;
        RECT 504.600 273.000 508.200 274.200 ;
        RECT 551.400 273.600 555.000 274.800 ;
        RECT 605.400 274.200 609.600 274.800 ;
        RECT 606.000 273.600 610.200 274.200 ;
        RECT 552.000 273.000 555.600 273.600 ;
        RECT 606.600 273.000 610.800 273.600 ;
        RECT 505.200 272.400 508.800 273.000 ;
        RECT 303.000 270.000 306.000 271.800 ;
        RECT 505.800 271.200 509.400 272.400 ;
        RECT 552.600 271.800 556.200 273.000 ;
        RECT 607.200 272.400 611.400 273.000 ;
        RECT 607.800 271.800 612.600 272.400 ;
        RECT 553.200 271.200 556.800 271.800 ;
        RECT 608.400 271.200 613.200 271.800 ;
        RECT 506.400 270.600 510.000 271.200 ;
        RECT 553.800 270.600 557.400 271.200 ;
        RECT 609.600 270.600 613.800 271.200 ;
        RECT 691.200 270.600 694.200 274.800 ;
        RECT 507.000 270.000 510.000 270.600 ;
        RECT 106.200 269.400 160.200 270.000 ;
        RECT 241.800 269.400 246.600 270.000 ;
        RECT 250.800 269.400 253.800 270.000 ;
        RECT 100.200 268.800 160.800 269.400 ;
        RECT 242.400 268.800 247.200 269.400 ;
        RECT 250.800 268.800 254.400 269.400 ;
        RECT 95.400 268.200 160.800 268.800 ;
        RECT 243.000 268.200 247.800 268.800 ;
        RECT 251.400 268.200 254.400 268.800 ;
        RECT 91.200 267.600 126.000 268.200 ;
        RECT 156.000 267.600 160.200 268.200 ;
        RECT 244.200 267.600 249.000 268.200 ;
        RECT 251.400 267.600 255.000 268.200 ;
        RECT 87.600 267.000 112.800 267.600 ;
        RECT 244.800 267.000 249.600 267.600 ;
        RECT 252.000 267.000 255.000 267.600 ;
        RECT 84.000 266.400 105.600 267.000 ;
        RECT 245.400 266.400 250.200 267.000 ;
        RECT 81.000 265.800 99.600 266.400 ;
        RECT 246.600 265.800 250.800 266.400 ;
        RECT 252.000 265.800 255.600 267.000 ;
        RECT 279.000 266.400 282.000 270.000 ;
        RECT 302.400 268.200 305.400 270.000 ;
        RECT 507.000 269.400 510.600 270.000 ;
        RECT 554.400 269.400 558.000 270.600 ;
        RECT 610.200 270.000 614.400 270.600 ;
        RECT 691.200 270.000 693.600 270.600 ;
        RECT 610.800 269.400 615.000 270.000 ;
        RECT 507.600 268.800 511.200 269.400 ;
        RECT 555.000 268.800 558.600 269.400 ;
        RECT 611.400 268.800 615.600 269.400 ;
        RECT 301.800 267.600 305.400 268.200 ;
        RECT 508.200 268.200 511.200 268.800 ;
        RECT 555.600 268.200 559.200 268.800 ;
        RECT 612.000 268.200 616.200 268.800 ;
        RECT 508.200 267.600 511.800 268.200 ;
        RECT 301.800 266.400 304.800 267.600 ;
        RECT 508.800 267.000 511.800 267.600 ;
        RECT 556.200 267.000 559.800 268.200 ;
        RECT 612.600 267.600 616.800 268.200 ;
        RECT 613.200 267.000 617.400 267.600 ;
        RECT 314.400 266.400 327.000 267.000 ;
        RECT 508.800 266.400 512.400 267.000 ;
        RECT 556.800 266.400 560.400 267.000 ;
        RECT 613.800 266.400 618.000 267.000 ;
        RECT 690.600 266.400 693.600 270.000 ;
        RECT 279.600 265.800 282.000 266.400 ;
        RECT 301.200 265.800 304.800 266.400 ;
        RECT 309.000 265.800 331.800 266.400 ;
        RECT 509.400 265.800 513.000 266.400 ;
        RECT 78.600 265.200 94.800 265.800 ;
        RECT 247.200 265.200 256.200 265.800 ;
        RECT 76.200 264.600 91.200 265.200 ;
        RECT 247.800 264.600 256.800 265.200 ;
        RECT 74.400 264.000 87.000 264.600 ;
        RECT 248.400 264.000 256.800 264.600 ;
        RECT 72.600 263.400 84.000 264.000 ;
        RECT 249.600 263.400 257.400 264.000 ;
        RECT 70.800 262.800 81.000 263.400 ;
        RECT 250.200 262.800 258.000 263.400 ;
        RECT 69.600 262.200 78.600 262.800 ;
        RECT 250.800 262.200 258.000 262.800 ;
        RECT 68.400 261.600 76.200 262.200 ;
        RECT 251.400 261.600 258.600 262.200 ;
        RECT 67.800 261.000 74.400 261.600 ;
        RECT 252.600 261.000 259.200 261.600 ;
        RECT 67.200 260.400 72.600 261.000 ;
        RECT 253.200 260.400 259.800 261.000 ;
        RECT 66.600 259.800 71.400 260.400 ;
        RECT 253.800 259.800 259.800 260.400 ;
        RECT 279.600 259.800 282.600 265.800 ;
        RECT 301.200 265.200 334.200 265.800 ;
        RECT 510.000 265.200 513.000 265.800 ;
        RECT 557.400 265.800 561.000 266.400 ;
        RECT 614.400 265.800 618.600 266.400 ;
        RECT 557.400 265.200 561.600 265.800 ;
        RECT 615.000 265.200 619.200 265.800 ;
        RECT 301.200 264.600 336.600 265.200 ;
        RECT 510.000 264.600 513.600 265.200 ;
        RECT 558.000 264.600 561.600 265.200 ;
        RECT 615.600 264.600 619.800 265.200 ;
        RECT 300.000 264.000 339.000 264.600 ;
        RECT 510.600 264.000 513.600 264.600 ;
        RECT 558.600 264.000 562.200 264.600 ;
        RECT 616.200 264.000 620.400 264.600 ;
        RECT 297.600 263.400 313.800 264.000 ;
        RECT 327.600 263.400 340.800 264.000 ;
        RECT 510.600 263.400 514.200 264.000 ;
        RECT 559.200 263.400 562.800 264.000 ;
        RECT 616.800 263.400 621.000 264.000 ;
        RECT 690.000 263.400 693.000 266.400 ;
        RECT 295.200 262.800 308.400 263.400 ;
        RECT 331.800 262.800 342.600 263.400 ;
        RECT 511.200 262.800 514.800 263.400 ;
        RECT 559.200 262.800 563.400 263.400 ;
        RECT 617.400 262.800 621.600 263.400 ;
        RECT 690.000 262.800 692.400 263.400 ;
        RECT 292.800 262.200 305.400 262.800 ;
        RECT 334.800 262.200 344.400 262.800 ;
        RECT 511.800 262.200 514.800 262.800 ;
        RECT 559.800 262.200 563.400 262.800 ;
        RECT 618.000 262.200 622.200 262.800 ;
        RECT 291.000 261.600 301.800 262.200 ;
        RECT 336.600 261.600 346.200 262.200 ;
        RECT 511.800 261.600 515.400 262.200 ;
        RECT 288.600 261.000 299.400 261.600 ;
        RECT 339.000 261.000 347.400 261.600 ;
        RECT 512.400 261.000 515.400 261.600 ;
        RECT 560.400 261.600 564.000 262.200 ;
        RECT 618.600 261.600 622.800 262.200 ;
        RECT 560.400 261.000 564.600 261.600 ;
        RECT 619.200 261.000 623.400 261.600 ;
        RECT 286.800 260.400 297.600 261.000 ;
        RECT 340.800 260.400 348.600 261.000 ;
        RECT 512.400 260.400 516.000 261.000 ;
        RECT 561.000 260.400 564.600 261.000 ;
        RECT 619.800 260.400 624.000 261.000 ;
        RECT 285.000 259.800 295.200 260.400 ;
        RECT 342.600 259.800 349.800 260.400 ;
        RECT 513.000 259.800 516.000 260.400 ;
        RECT 561.600 259.800 565.200 260.400 ;
        RECT 620.400 259.800 624.600 260.400 ;
        RECT 689.400 259.800 692.400 262.800 ;
        RECT 66.600 259.200 70.200 259.800 ;
        RECT 254.400 259.200 260.400 259.800 ;
        RECT 280.200 259.200 292.800 259.800 ;
        RECT 343.800 259.200 351.000 259.800 ;
        RECT 513.000 259.200 516.600 259.800 ;
        RECT 562.200 259.200 565.800 259.800 ;
        RECT 621.000 259.200 625.200 259.800 ;
        RECT 66.000 258.600 70.200 259.200 ;
        RECT 255.000 258.600 261.000 259.200 ;
        RECT 280.200 258.600 291.000 259.200 ;
        RECT 345.600 258.600 352.200 259.200 ;
        RECT 513.600 258.600 517.200 259.200 ;
        RECT 66.600 258.000 70.200 258.600 ;
        RECT 255.600 258.000 261.000 258.600 ;
        RECT 279.600 258.000 289.200 258.600 ;
        RECT 346.800 258.000 353.400 258.600 ;
        RECT 514.200 258.000 517.200 258.600 ;
        RECT 562.800 258.600 565.800 259.200 ;
        RECT 621.600 258.600 625.800 259.200 ;
        RECT 562.800 258.000 566.400 258.600 ;
        RECT 622.200 258.000 626.400 258.600 ;
        RECT 66.600 257.400 71.400 258.000 ;
        RECT 256.800 257.400 261.600 258.000 ;
        RECT 278.400 257.400 287.400 258.000 ;
        RECT 348.000 257.400 354.600 258.000 ;
        RECT 514.200 257.400 517.800 258.000 ;
        RECT 563.400 257.400 567.000 258.000 ;
        RECT 622.800 257.400 627.000 258.000 ;
        RECT 688.800 257.400 691.800 259.800 ;
        RECT 67.200 256.800 72.600 257.400 ;
        RECT 257.400 256.800 261.600 257.400 ;
        RECT 276.600 256.800 285.600 257.400 ;
        RECT 349.200 256.800 355.200 257.400 ;
        RECT 514.800 256.800 517.800 257.400 ;
        RECT 564.000 256.800 567.000 257.400 ;
        RECT 623.400 256.800 627.600 257.400 ;
        RECT 688.800 256.800 691.200 257.400 ;
        RECT 67.200 256.200 74.400 256.800 ;
        RECT 183.600 256.200 194.400 256.800 ;
        RECT 258.000 256.200 262.200 256.800 ;
        RECT 275.400 256.200 283.800 256.800 ;
        RECT 350.400 256.200 356.400 256.800 ;
        RECT 514.800 256.200 518.400 256.800 ;
        RECT 564.000 256.200 567.600 256.800 ;
        RECT 624.000 256.200 628.200 256.800 ;
        RECT 68.400 255.600 76.800 256.200 ;
        RECT 177.600 255.600 195.600 256.200 ;
        RECT 258.600 255.600 262.800 256.200 ;
        RECT 274.200 255.600 282.000 256.200 ;
        RECT 351.600 255.600 357.000 256.200 ;
        RECT 515.400 255.600 518.400 256.200 ;
        RECT 564.600 255.600 568.200 256.200 ;
        RECT 624.600 255.600 628.800 256.200 ;
        RECT 69.600 255.000 78.600 255.600 ;
        RECT 172.800 255.000 195.600 255.600 ;
        RECT 259.200 255.000 263.400 255.600 ;
        RECT 272.400 255.000 280.200 255.600 ;
        RECT 352.800 255.000 358.200 255.600 ;
        RECT 515.400 255.000 519.000 255.600 ;
        RECT 70.800 254.400 81.600 255.000 ;
        RECT 168.000 254.400 195.600 255.000 ;
        RECT 259.800 254.400 264.000 255.000 ;
        RECT 271.800 254.400 278.400 255.000 ;
        RECT 353.400 254.400 358.800 255.000 ;
        RECT 516.000 254.400 519.000 255.000 ;
        RECT 565.200 255.000 568.200 255.600 ;
        RECT 625.200 255.000 629.400 255.600 ;
        RECT 565.200 254.400 568.800 255.000 ;
        RECT 625.800 254.400 630.000 255.000 ;
        RECT 688.200 254.400 691.200 256.800 ;
        RECT 72.600 253.800 84.000 254.400 ;
        RECT 163.800 253.800 190.800 254.400 ;
        RECT 260.400 253.800 264.600 254.400 ;
        RECT 270.600 253.800 277.200 254.400 ;
        RECT 354.600 253.800 359.400 254.400 ;
        RECT 516.000 253.800 519.600 254.400 ;
        RECT 74.400 253.200 87.000 253.800 ;
        RECT 160.200 253.200 183.000 253.800 ;
        RECT 261.000 253.200 265.200 253.800 ;
        RECT 269.400 253.200 276.000 253.800 ;
        RECT 355.200 253.200 360.000 253.800 ;
        RECT 516.600 253.200 519.600 253.800 ;
        RECT 565.800 253.800 569.400 254.400 ;
        RECT 626.400 253.800 630.600 254.400 ;
        RECT 565.800 253.200 570.000 253.800 ;
        RECT 627.000 253.200 631.200 253.800 ;
        RECT 76.800 252.600 90.000 253.200 ;
        RECT 156.000 252.600 177.000 253.200 ;
        RECT 261.600 252.600 265.800 253.200 ;
        RECT 268.200 252.600 274.800 253.200 ;
        RECT 356.400 252.600 360.600 253.200 ;
        RECT 516.600 252.600 520.200 253.200 ;
        RECT 566.400 252.600 570.000 253.200 ;
        RECT 627.600 252.600 631.800 253.200 ;
        RECT 78.600 252.000 93.000 252.600 ;
        RECT 152.400 252.000 172.200 252.600 ;
        RECT 262.800 252.000 265.800 252.600 ;
        RECT 267.000 252.000 273.600 252.600 ;
        RECT 357.000 252.000 361.200 252.600 ;
        RECT 517.200 252.000 520.200 252.600 ;
        RECT 81.000 251.400 96.600 252.000 ;
        RECT 148.800 251.400 168.000 252.000 ;
        RECT 263.400 251.400 272.400 252.000 ;
        RECT 357.600 251.400 361.200 252.000 ;
        RECT 517.800 251.400 520.800 252.000 ;
        RECT 567.000 251.400 570.600 252.600 ;
        RECT 628.200 252.000 632.400 252.600 ;
        RECT 687.600 252.000 690.600 254.400 ;
        RECT 628.800 251.400 633.000 252.000 ;
        RECT 84.000 250.800 100.800 251.400 ;
        RECT 145.200 250.800 163.800 251.400 ;
        RECT 264.000 250.800 271.200 251.400 ;
        RECT 358.200 250.800 361.800 251.400 ;
        RECT 517.800 250.800 521.400 251.400 ;
        RECT 567.600 250.800 571.200 251.400 ;
        RECT 629.400 250.800 633.600 251.400 ;
        RECT 87.000 250.200 105.600 250.800 ;
        RECT 141.600 250.200 159.600 250.800 ;
        RECT 264.000 250.200 270.000 250.800 ;
        RECT 358.200 250.200 362.400 250.800 ;
        RECT 90.000 249.600 112.800 250.200 ;
        RECT 137.400 249.600 156.000 250.200 ;
        RECT 218.400 249.600 225.000 250.200 ;
        RECT 263.400 249.600 268.800 250.200 ;
        RECT 358.800 249.600 362.400 250.200 ;
        RECT 518.400 250.200 521.400 250.800 ;
        RECT 568.200 250.200 571.200 250.800 ;
        RECT 630.000 250.200 634.200 250.800 ;
        RECT 518.400 249.600 522.000 250.200 ;
        RECT 568.200 249.600 571.800 250.200 ;
        RECT 630.600 249.600 634.800 250.200 ;
        RECT 687.000 249.600 690.000 252.000 ;
        RECT 93.000 249.000 152.400 249.600 ;
        RECT 215.400 249.000 225.000 249.600 ;
        RECT 262.200 249.000 267.600 249.600 ;
        RECT 96.600 248.400 148.800 249.000 ;
        RECT 213.000 248.400 225.000 249.000 ;
        RECT 261.600 248.400 267.000 249.000 ;
        RECT 359.400 248.400 363.000 249.600 ;
        RECT 519.000 249.000 522.000 249.600 ;
        RECT 568.800 249.000 571.800 249.600 ;
        RECT 631.200 249.000 635.400 249.600 ;
        RECT 519.000 248.400 522.600 249.000 ;
        RECT 568.800 248.400 572.400 249.000 ;
        RECT 631.800 248.400 636.000 249.000 ;
        RECT 100.800 247.800 145.200 248.400 ;
        RECT 210.600 247.800 223.800 248.400 ;
        RECT 260.400 247.800 265.800 248.400 ;
        RECT 360.000 247.800 363.000 248.400 ;
        RECT 106.200 247.200 141.600 247.800 ;
        RECT 208.800 247.200 221.400 247.800 ;
        RECT 259.800 247.200 264.600 247.800 ;
        RECT 360.000 247.200 363.600 247.800 ;
        RECT 519.600 247.200 522.600 248.400 ;
        RECT 569.400 247.800 573.000 248.400 ;
        RECT 632.400 247.800 636.000 248.400 ;
        RECT 570.000 247.200 573.000 247.800 ;
        RECT 633.000 247.200 636.600 247.800 ;
        RECT 686.400 247.200 689.400 249.600 ;
        RECT 114.000 246.600 138.000 247.200 ;
        RECT 206.400 246.600 218.400 247.200 ;
        RECT 258.600 246.600 264.000 247.200 ;
        RECT 360.600 246.600 363.600 247.200 ;
        RECT 114.000 246.000 134.400 246.600 ;
        RECT 204.600 246.000 215.400 246.600 ;
        RECT 258.000 246.000 262.800 246.600 ;
        RECT 360.600 246.000 364.200 246.600 ;
        RECT 114.000 245.400 130.800 246.000 ;
        RECT 202.200 245.400 213.000 246.000 ;
        RECT 257.400 245.400 262.200 246.000 ;
        RECT 361.200 245.400 364.200 246.000 ;
        RECT 520.200 246.000 523.200 247.200 ;
        RECT 570.000 246.600 573.600 247.200 ;
        RECT 633.600 246.600 637.200 247.200 ;
        RECT 570.600 246.000 573.600 246.600 ;
        RECT 634.200 246.000 637.800 246.600 ;
        RECT 520.200 245.400 523.800 246.000 ;
        RECT 570.600 245.400 574.200 246.000 ;
        RECT 111.000 244.800 127.800 245.400 ;
        RECT 200.400 244.800 210.600 245.400 ;
        RECT 256.200 244.800 261.000 245.400 ;
        RECT 361.200 244.800 364.800 245.400 ;
        RECT 108.000 244.200 124.200 244.800 ;
        RECT 198.600 244.200 208.800 244.800 ;
        RECT 255.600 244.200 260.400 244.800 ;
        RECT 361.800 244.200 364.800 244.800 ;
        RECT 520.800 244.800 523.800 245.400 ;
        RECT 571.200 244.800 574.200 245.400 ;
        RECT 634.800 245.400 638.400 246.000 ;
        RECT 634.800 244.800 639.000 245.400 ;
        RECT 685.800 244.800 688.800 247.200 ;
        RECT 520.800 244.200 524.400 244.800 ;
        RECT 571.200 244.200 574.800 244.800 ;
        RECT 635.400 244.200 639.600 244.800 ;
        RECT 104.400 243.600 120.600 244.200 ;
        RECT 196.800 243.600 206.400 244.200 ;
        RECT 255.000 243.600 259.800 244.200 ;
        RECT 361.800 243.600 365.400 244.200 ;
        RECT 101.400 243.000 117.600 243.600 ;
        RECT 195.000 243.000 204.600 243.600 ;
        RECT 254.400 243.000 258.600 243.600 ;
        RECT 98.400 242.400 114.000 243.000 ;
        RECT 193.200 242.400 202.800 243.000 ;
        RECT 253.200 242.400 258.000 243.000 ;
        RECT 362.400 242.400 365.400 243.600 ;
        RECT 521.400 243.600 524.400 244.200 ;
        RECT 571.800 243.600 574.800 244.200 ;
        RECT 636.000 243.600 640.200 244.200 ;
        RECT 521.400 243.000 525.000 243.600 ;
        RECT 571.800 243.000 575.400 243.600 ;
        RECT 636.600 243.000 640.800 243.600 ;
        RECT 685.200 243.000 688.200 244.800 ;
        RECT 522.000 242.400 525.000 243.000 ;
        RECT 572.400 242.400 575.400 243.000 ;
        RECT 637.200 242.400 640.800 243.000 ;
        RECT 684.600 242.400 688.200 243.000 ;
        RECT 95.400 241.800 111.000 242.400 ;
        RECT 191.400 241.800 200.400 242.400 ;
        RECT 252.600 241.800 257.400 242.400 ;
        RECT 93.000 241.200 107.400 241.800 ;
        RECT 189.600 241.200 198.600 241.800 ;
        RECT 252.000 241.200 256.800 241.800 ;
        RECT 363.000 241.200 366.000 242.400 ;
        RECT 522.000 241.800 525.600 242.400 ;
        RECT 572.400 241.800 576.000 242.400 ;
        RECT 637.800 241.800 641.400 242.400 ;
        RECT 90.000 240.600 104.400 241.200 ;
        RECT 187.800 240.600 196.800 241.200 ;
        RECT 251.400 240.600 255.600 241.200 ;
        RECT 363.000 240.600 366.600 241.200 ;
        RECT 522.600 240.600 525.600 241.800 ;
        RECT 573.000 241.200 576.000 241.800 ;
        RECT 638.400 241.200 642.000 241.800 ;
        RECT 573.000 240.600 576.600 241.200 ;
        RECT 87.000 240.000 101.400 240.600 ;
        RECT 186.000 240.000 195.000 240.600 ;
        RECT 250.800 240.000 255.000 240.600 ;
        RECT 84.600 239.400 98.400 240.000 ;
        RECT 184.800 239.400 193.200 240.000 ;
        RECT 250.200 239.400 254.400 240.000 ;
        RECT 363.600 239.400 366.600 240.600 ;
        RECT 523.200 239.400 526.200 240.600 ;
        RECT 573.600 240.000 576.600 240.600 ;
        RECT 639.000 240.600 642.600 241.200 ;
        RECT 684.600 240.600 687.600 242.400 ;
        RECT 639.000 240.000 643.200 240.600 ;
        RECT 573.600 239.400 577.200 240.000 ;
        RECT 639.600 239.400 643.800 240.000 ;
        RECT 82.200 238.800 95.400 239.400 ;
        RECT 183.000 238.800 191.400 239.400 ;
        RECT 249.600 238.800 253.800 239.400 ;
        RECT 363.600 238.800 367.200 239.400 ;
        RECT 523.200 238.800 526.800 239.400 ;
        RECT 79.800 238.200 93.000 238.800 ;
        RECT 181.200 238.200 190.200 238.800 ;
        RECT 249.000 238.200 253.200 238.800 ;
        RECT 77.400 237.600 90.000 238.200 ;
        RECT 180.000 237.600 188.400 238.200 ;
        RECT 248.400 237.600 252.600 238.200 ;
        RECT 75.000 237.000 87.600 237.600 ;
        RECT 178.200 237.000 186.600 237.600 ;
        RECT 247.800 237.000 252.000 237.600 ;
        RECT 364.200 237.000 367.200 238.800 ;
        RECT 523.800 238.200 526.800 238.800 ;
        RECT 574.200 238.800 577.200 239.400 ;
        RECT 640.200 238.800 644.400 239.400 ;
        RECT 684.000 238.800 687.000 240.600 ;
        RECT 574.200 238.200 577.800 238.800 ;
        RECT 640.800 238.200 644.400 238.800 ;
        RECT 683.400 238.200 687.000 238.800 ;
        RECT 523.800 237.600 527.400 238.200 ;
        RECT 73.200 236.400 84.600 237.000 ;
        RECT 176.400 236.400 184.800 237.000 ;
        RECT 247.200 236.400 251.400 237.000 ;
        RECT 70.800 235.800 82.200 236.400 ;
        RECT 175.200 235.800 183.600 236.400 ;
        RECT 246.600 235.800 250.800 236.400 ;
        RECT 69.000 235.200 79.800 235.800 ;
        RECT 173.400 235.200 181.800 235.800 ;
        RECT 246.000 235.200 250.200 235.800 ;
        RECT 364.800 235.200 367.800 237.000 ;
        RECT 524.400 236.400 527.400 237.600 ;
        RECT 574.800 237.600 577.800 238.200 ;
        RECT 641.400 237.600 645.000 238.200 ;
        RECT 574.800 237.000 578.400 237.600 ;
        RECT 642.000 237.000 645.600 237.600 ;
        RECT 683.400 237.000 686.400 238.200 ;
        RECT 575.400 236.400 578.400 237.000 ;
        RECT 642.600 236.400 646.200 237.000 ;
        RECT 682.800 236.400 686.400 237.000 ;
        RECT 525.000 235.200 528.000 236.400 ;
        RECT 575.400 235.800 579.000 236.400 ;
        RECT 642.600 235.800 646.800 236.400 ;
        RECT 66.600 234.600 77.400 235.200 ;
        RECT 172.200 234.600 180.000 235.200 ;
        RECT 245.400 234.600 249.600 235.200 ;
        RECT 64.800 234.000 75.000 234.600 ;
        RECT 170.400 234.000 178.800 234.600 ;
        RECT 244.800 234.000 249.000 234.600 ;
        RECT 63.000 233.400 73.200 234.000 ;
        RECT 169.200 233.400 177.000 234.000 ;
        RECT 244.200 233.400 248.400 234.000 ;
        RECT 61.200 232.800 70.800 233.400 ;
        RECT 167.400 232.800 175.800 233.400 ;
        RECT 243.600 232.800 247.800 233.400 ;
        RECT 365.400 232.800 368.400 235.200 ;
        RECT 525.000 234.600 528.600 235.200 ;
        RECT 576.000 234.600 579.000 235.800 ;
        RECT 643.200 235.200 647.400 235.800 ;
        RECT 643.800 234.600 647.400 235.200 ;
        RECT 682.800 234.600 685.800 236.400 ;
        RECT 525.600 233.400 528.600 234.600 ;
        RECT 576.600 233.400 579.600 234.600 ;
        RECT 644.400 234.000 648.000 234.600 ;
        RECT 645.000 233.400 648.600 234.000 ;
        RECT 525.600 232.800 529.200 233.400 ;
        RECT 576.600 232.800 580.200 233.400 ;
        RECT 645.000 232.800 649.200 233.400 ;
        RECT 682.200 232.800 685.200 234.600 ;
        RECT 59.400 232.200 69.000 232.800 ;
        RECT 166.200 232.200 174.000 232.800 ;
        RECT 243.600 232.200 247.200 232.800 ;
        RECT 58.200 231.600 67.200 232.200 ;
        RECT 165.000 231.600 172.800 232.200 ;
        RECT 243.000 231.600 246.600 232.200 ;
        RECT 57.000 231.000 65.400 231.600 ;
        RECT 163.200 231.000 171.000 231.600 ;
        RECT 242.400 231.000 246.000 231.600 ;
        RECT 55.800 230.400 63.600 231.000 ;
        RECT 162.000 230.400 169.800 231.000 ;
        RECT 241.800 230.400 245.400 231.000 ;
        RECT 366.000 230.400 369.000 232.800 ;
        RECT 526.200 231.600 529.200 232.800 ;
        RECT 577.200 232.200 580.200 232.800 ;
        RECT 645.600 232.200 649.800 232.800 ;
        RECT 577.200 231.600 580.800 232.200 ;
        RECT 646.200 231.600 649.800 232.200 ;
        RECT 54.600 229.800 61.800 230.400 ;
        RECT 160.200 229.800 168.000 230.400 ;
        RECT 241.200 229.800 245.400 230.400 ;
        RECT 54.000 229.200 60.000 229.800 ;
        RECT 159.000 229.200 166.800 229.800 ;
        RECT 240.600 229.200 244.800 229.800 ;
        RECT 53.400 228.600 58.800 229.200 ;
        RECT 157.800 228.600 165.000 229.200 ;
        RECT 240.600 228.600 244.200 229.200 ;
        RECT 52.800 228.000 57.600 228.600 ;
        RECT 156.000 228.000 163.800 228.600 ;
        RECT 240.000 228.000 243.600 228.600 ;
        RECT 366.600 228.000 369.600 230.400 ;
        RECT 526.800 229.800 529.800 231.600 ;
        RECT 577.800 230.400 580.800 231.600 ;
        RECT 646.800 231.000 650.400 231.600 ;
        RECT 681.600 231.000 684.600 232.800 ;
        RECT 647.400 230.400 651.000 231.000 ;
        RECT 527.400 228.000 530.400 229.800 ;
        RECT 578.400 229.200 581.400 230.400 ;
        RECT 648.000 229.800 651.600 230.400 ;
        RECT 681.000 229.800 684.000 231.000 ;
        RECT 648.000 229.200 652.200 229.800 ;
        RECT 578.400 228.600 582.000 229.200 ;
        RECT 648.600 228.600 652.200 229.200 ;
        RECT 680.400 229.200 684.000 229.800 ;
        RECT 52.200 227.400 56.400 228.000 ;
        RECT 154.800 227.400 162.000 228.000 ;
        RECT 239.400 227.400 243.000 228.000 ;
        RECT 51.600 226.800 55.800 227.400 ;
        RECT 153.600 226.800 160.800 227.400 ;
        RECT 51.600 225.600 55.200 226.800 ;
        RECT 151.800 226.200 159.600 226.800 ;
        RECT 238.800 226.200 242.400 227.400 ;
        RECT 150.600 225.600 157.800 226.200 ;
        RECT 238.200 225.600 241.800 226.200 ;
        RECT 51.600 225.000 55.800 225.600 ;
        RECT 149.400 225.000 156.600 225.600 ;
        RECT 237.600 225.000 241.200 225.600 ;
        RECT 367.200 225.000 370.200 228.000 ;
        RECT 528.000 226.200 531.000 228.000 ;
        RECT 579.000 227.400 582.000 228.600 ;
        RECT 649.200 228.000 652.800 228.600 ;
        RECT 680.400 228.000 683.400 229.200 ;
        RECT 649.800 227.400 653.400 228.000 ;
        RECT 679.800 227.400 683.400 228.000 ;
        RECT 579.000 226.800 582.600 227.400 ;
        RECT 52.200 224.400 57.600 225.000 ;
        RECT 148.200 224.400 154.800 225.000 ;
        RECT 52.200 223.800 59.400 224.400 ;
        RECT 146.400 223.800 153.000 224.400 ;
        RECT 237.000 223.800 240.600 225.000 ;
        RECT 53.400 223.200 61.200 223.800 ;
        RECT 145.200 223.200 151.800 223.800 ;
        RECT 236.400 223.200 240.000 223.800 ;
        RECT 54.000 222.600 63.600 223.200 ;
        RECT 144.000 222.600 150.600 223.200 ;
        RECT 55.200 222.000 66.600 222.600 ;
        RECT 142.800 222.000 149.400 222.600 ;
        RECT 235.800 222.000 239.400 223.200 ;
        RECT 57.000 221.400 70.200 222.000 ;
        RECT 141.600 221.400 148.200 222.000 ;
        RECT 234.600 221.400 238.800 222.000 ;
        RECT 58.800 220.800 73.800 221.400 ;
        RECT 139.800 220.800 147.600 221.400 ;
        RECT 233.400 220.800 238.200 221.400 ;
        RECT 61.200 220.200 78.600 220.800 ;
        RECT 135.600 220.200 146.400 220.800 ;
        RECT 231.600 220.200 238.200 220.800 ;
        RECT 334.200 220.200 334.800 222.000 ;
        RECT 367.800 221.400 370.800 225.000 ;
        RECT 528.600 223.800 531.600 226.200 ;
        RECT 579.600 225.600 582.600 226.800 ;
        RECT 650.400 226.800 654.000 227.400 ;
        RECT 650.400 226.200 654.600 226.800 ;
        RECT 679.800 226.200 682.800 227.400 ;
        RECT 651.000 225.600 654.600 226.200 ;
        RECT 679.200 225.600 682.800 226.200 ;
        RECT 580.200 223.800 583.200 225.600 ;
        RECT 651.600 225.000 655.200 225.600 ;
        RECT 652.200 224.400 655.800 225.000 ;
        RECT 679.200 224.400 682.200 225.600 ;
        RECT 652.800 223.800 656.400 224.400 ;
        RECT 529.200 222.000 532.200 223.800 ;
        RECT 580.800 222.000 583.800 223.800 ;
        RECT 652.800 223.200 657.000 223.800 ;
        RECT 678.600 223.200 681.600 224.400 ;
        RECT 653.400 222.600 657.000 223.200 ;
        RECT 678.000 222.600 681.600 223.200 ;
        RECT 654.000 222.000 657.600 222.600 ;
        RECT 529.200 221.400 532.800 222.000 ;
        RECT 63.600 219.600 84.000 220.200 ;
        RECT 128.400 219.600 144.600 220.200 ;
        RECT 230.400 219.600 237.600 220.200 ;
        RECT 334.200 219.600 335.400 220.200 ;
        RECT 66.600 219.000 91.200 219.600 ;
        RECT 120.000 219.000 143.400 219.600 ;
        RECT 228.600 219.000 237.000 219.600 ;
        RECT 70.200 218.400 141.600 219.000 ;
        RECT 227.400 218.400 237.000 219.000 ;
        RECT 74.400 217.800 140.400 218.400 ;
        RECT 225.600 217.800 236.400 218.400 ;
        RECT 78.600 217.200 129.600 217.800 ;
        RECT 130.800 217.200 139.200 217.800 ;
        RECT 224.400 217.200 235.800 217.800 ;
        RECT 84.600 216.600 124.800 217.200 ;
        RECT 130.800 216.600 138.000 217.200 ;
        RECT 222.600 216.600 229.800 217.200 ;
        RECT 232.200 216.600 235.800 217.200 ;
        RECT 333.600 216.600 335.400 219.600 ;
        RECT 368.400 217.800 371.400 221.400 ;
        RECT 529.800 219.000 532.800 221.400 ;
        RECT 581.400 220.200 584.400 222.000 ;
        RECT 654.600 221.400 658.200 222.000 ;
        RECT 678.000 221.400 681.000 222.600 ;
        RECT 655.200 220.800 658.800 221.400 ;
        RECT 677.400 220.800 681.000 221.400 ;
        RECT 655.200 220.200 659.400 220.800 ;
        RECT 581.400 219.600 585.000 220.200 ;
        RECT 655.800 219.600 659.400 220.200 ;
        RECT 677.400 219.600 680.400 220.800 ;
        RECT 91.800 216.000 118.200 216.600 ;
        RECT 129.600 216.000 136.800 216.600 ;
        RECT 220.800 216.000 228.600 216.600 ;
        RECT 232.200 216.000 235.200 216.600 ;
        RECT 128.400 215.400 135.600 216.000 ;
        RECT 219.600 215.400 226.800 216.000 ;
        RECT 231.600 215.400 235.200 216.000 ;
        RECT 127.200 214.800 134.400 215.400 ;
        RECT 217.800 214.800 225.600 215.400 ;
        RECT 231.600 214.800 234.600 215.400 ;
        RECT 126.000 214.200 132.600 214.800 ;
        RECT 216.000 214.200 223.800 214.800 ;
        RECT 231.000 214.200 234.600 214.800 ;
        RECT 124.800 213.600 131.400 214.200 ;
        RECT 214.800 213.600 222.600 214.200 ;
        RECT 231.000 213.600 234.000 214.200 ;
        RECT 123.600 213.000 130.200 213.600 ;
        RECT 213.000 213.000 220.800 213.600 ;
        RECT 230.400 213.000 234.000 213.600 ;
        RECT 333.000 213.000 335.400 216.600 ;
        RECT 369.000 214.200 372.000 217.800 ;
        RECT 530.400 216.600 533.400 219.000 ;
        RECT 582.000 217.800 585.000 219.600 ;
        RECT 656.400 219.000 660.000 219.600 ;
        RECT 657.000 218.400 660.600 219.000 ;
        RECT 676.800 218.400 679.800 219.600 ;
        RECT 657.600 217.800 661.200 218.400 ;
        RECT 676.200 217.800 679.800 218.400 ;
        RECT 122.400 212.400 129.000 213.000 ;
        RECT 211.200 212.400 219.600 213.000 ;
        RECT 230.400 212.400 233.400 213.000 ;
        RECT 121.200 211.800 127.800 212.400 ;
        RECT 209.400 211.800 217.800 212.400 ;
        RECT 229.800 211.800 233.400 212.400 ;
        RECT 332.400 212.400 335.400 213.000 ;
        RECT 369.600 213.600 372.000 214.200 ;
        RECT 120.000 211.200 126.600 211.800 ;
        RECT 207.600 211.200 216.600 211.800 ;
        RECT 229.800 211.200 232.800 211.800 ;
        RECT 118.800 210.600 125.400 211.200 ;
        RECT 205.800 210.600 214.800 211.200 ;
        RECT 229.200 210.600 232.800 211.200 ;
        RECT 117.600 210.000 124.200 210.600 ;
        RECT 204.600 210.000 213.000 210.600 ;
        RECT 229.200 210.000 232.200 210.600 ;
        RECT 116.400 209.400 123.000 210.000 ;
        RECT 202.800 209.400 211.200 210.000 ;
        RECT 228.600 209.400 232.200 210.000 ;
        RECT 332.400 209.400 334.800 212.400 ;
        RECT 369.600 209.400 372.600 213.600 ;
        RECT 531.000 213.000 534.000 216.600 ;
        RECT 582.600 215.400 585.600 217.800 ;
        RECT 657.600 217.200 661.800 217.800 ;
        RECT 676.200 217.200 679.200 217.800 ;
        RECT 658.200 216.600 661.800 217.200 ;
        RECT 675.600 216.600 679.200 217.200 ;
        RECT 658.800 216.000 662.400 216.600 ;
        RECT 659.400 215.400 663.000 216.000 ;
        RECT 675.600 215.400 678.600 216.600 ;
        RECT 583.200 213.000 586.200 215.400 ;
        RECT 660.000 214.800 663.600 215.400 ;
        RECT 675.000 214.800 678.600 215.400 ;
        RECT 660.000 214.200 664.200 214.800 ;
        RECT 675.000 214.200 678.000 214.800 ;
        RECT 660.600 213.600 664.200 214.200 ;
        RECT 674.400 213.600 678.000 214.200 ;
        RECT 661.200 213.000 664.800 213.600 ;
        RECT 674.400 213.000 677.400 213.600 ;
        RECT 115.200 208.800 121.800 209.400 ;
        RECT 200.400 208.800 210.000 209.400 ;
        RECT 228.600 208.800 231.600 209.400 ;
        RECT 114.000 208.200 120.600 208.800 ;
        RECT 198.600 208.200 208.200 208.800 ;
        RECT 228.000 208.200 231.600 208.800 ;
        RECT 113.400 207.600 119.400 208.200 ;
        RECT 196.800 207.600 206.400 208.200 ;
        RECT 228.000 207.600 231.000 208.200 ;
        RECT 112.200 207.000 118.200 207.600 ;
        RECT 195.000 207.000 204.600 207.600 ;
        RECT 227.400 207.000 231.000 207.600 ;
        RECT 111.000 206.400 117.000 207.000 ;
        RECT 193.200 206.400 202.800 207.000 ;
        RECT 109.800 205.800 115.800 206.400 ;
        RECT 190.800 205.800 201.000 206.400 ;
        RECT 227.400 205.800 230.400 207.000 ;
        RECT 331.800 206.400 334.800 209.400 ;
        RECT 370.200 208.800 372.600 209.400 ;
        RECT 531.600 208.800 534.600 213.000 ;
        RECT 583.800 210.000 586.800 213.000 ;
        RECT 661.800 212.400 665.400 213.000 ;
        RECT 673.800 212.400 677.400 213.000 ;
        RECT 662.400 211.800 666.000 212.400 ;
        RECT 662.400 211.200 666.600 211.800 ;
        RECT 673.800 211.200 676.800 212.400 ;
        RECT 663.000 210.600 666.600 211.200 ;
        RECT 663.600 210.000 667.200 210.600 ;
        RECT 673.200 210.000 676.200 211.200 ;
        RECT 331.800 205.800 334.200 206.400 ;
        RECT 108.600 205.200 114.600 205.800 ;
        RECT 189.000 205.200 199.200 205.800 ;
        RECT 107.400 204.600 114.000 205.200 ;
        RECT 186.600 204.600 196.800 205.200 ;
        RECT 226.800 204.600 229.800 205.800 ;
        RECT 106.800 204.000 112.800 204.600 ;
        RECT 184.800 204.000 195.000 204.600 ;
        RECT 226.200 204.000 229.800 204.600 ;
        RECT 105.600 203.400 111.600 204.000 ;
        RECT 182.400 203.400 193.200 204.000 ;
        RECT 104.400 202.800 110.400 203.400 ;
        RECT 180.000 202.800 191.400 203.400 ;
        RECT 226.200 202.800 229.200 204.000 ;
        RECT 331.200 202.800 334.200 205.800 ;
        RECT 370.200 203.400 373.200 208.800 ;
        RECT 531.600 208.200 535.200 208.800 ;
        RECT 532.200 205.800 535.200 208.200 ;
        RECT 584.400 207.000 587.400 210.000 ;
        RECT 664.200 209.400 667.800 210.000 ;
        RECT 672.600 209.400 676.200 210.000 ;
        RECT 664.200 208.800 668.400 209.400 ;
        RECT 672.600 208.800 675.600 209.400 ;
        RECT 664.800 208.200 668.400 208.800 ;
        RECT 672.000 208.200 675.600 208.800 ;
        RECT 665.400 207.600 669.000 208.200 ;
        RECT 672.000 207.600 675.000 208.200 ;
        RECT 666.000 207.000 669.600 207.600 ;
        RECT 671.400 207.000 675.000 207.600 ;
        RECT 532.200 204.000 534.600 205.800 ;
        RECT 103.200 202.200 109.200 202.800 ;
        RECT 177.600 202.200 189.000 202.800 ;
        RECT 225.600 202.200 229.200 202.800 ;
        RECT 102.600 201.600 108.000 202.200 ;
        RECT 175.800 201.600 187.200 202.200 ;
        RECT 101.400 201.000 107.400 201.600 ;
        RECT 172.800 201.000 184.800 201.600 ;
        RECT 225.600 201.000 228.600 202.200 ;
        RECT 100.200 200.400 106.200 201.000 ;
        RECT 170.400 200.400 184.800 201.000 ;
        RECT 99.600 199.800 105.000 200.400 ;
        RECT 168.000 199.800 180.000 200.400 ;
        RECT 98.400 199.200 103.800 199.800 ;
        RECT 165.000 199.200 178.200 199.800 ;
        RECT 97.800 198.600 103.200 199.200 ;
        RECT 162.600 198.600 175.800 199.200 ;
        RECT 96.600 198.000 102.000 198.600 ;
        RECT 159.600 198.000 173.400 198.600 ;
        RECT 96.000 197.400 100.800 198.000 ;
        RECT 156.600 197.400 170.400 198.000 ;
        RECT 94.800 196.800 100.200 197.400 ;
        RECT 153.600 196.800 168.000 197.400 ;
        RECT 94.200 196.200 99.000 196.800 ;
        RECT 150.000 196.200 165.000 196.800 ;
        RECT 93.600 195.600 98.400 196.200 ;
        RECT 147.000 195.600 162.600 196.200 ;
        RECT 93.000 195.000 97.200 195.600 ;
        RECT 142.800 195.000 159.600 195.600 ;
        RECT 92.400 194.400 96.600 195.000 ;
        RECT 139.200 194.400 156.600 195.000 ;
        RECT 92.400 193.800 96.000 194.400 ;
        RECT 135.000 193.800 153.600 194.400 ;
        RECT 91.800 192.600 95.400 193.800 ;
        RECT 129.600 193.200 150.000 193.800 ;
        RECT 124.200 192.600 146.400 193.200 ;
        RECT 91.800 192.000 97.200 192.600 ;
        RECT 117.600 192.000 142.800 192.600 ;
        RECT 92.400 191.400 138.600 192.000 ;
        RECT 92.400 190.800 134.400 191.400 ;
        RECT 93.600 190.200 129.600 190.800 ;
        RECT 94.800 189.600 123.600 190.200 ;
        RECT 97.800 189.000 116.400 189.600 ;
        RECT 181.800 180.600 184.800 200.400 ;
        RECT 225.000 199.200 228.000 201.000 ;
        RECT 330.600 199.800 333.600 202.800 ;
        RECT 370.200 201.000 373.800 203.400 ;
        RECT 224.400 196.800 227.400 199.200 ;
        RECT 330.000 197.400 333.000 199.800 ;
        RECT 370.800 199.200 373.800 201.000 ;
        RECT 401.400 199.800 415.200 200.400 ;
        RECT 392.400 199.200 416.400 199.800 ;
        RECT 370.800 198.600 378.600 199.200 ;
        RECT 385.200 198.600 417.000 199.200 ;
        RECT 370.800 198.000 417.600 198.600 ;
        RECT 370.800 197.400 418.200 198.000 ;
        RECT 329.400 196.800 333.000 197.400 ;
        RECT 371.400 196.800 400.200 197.400 ;
        RECT 414.600 196.800 419.400 197.400 ;
        RECT 531.600 196.800 534.600 204.000 ;
        RECT 585.000 202.800 588.000 207.000 ;
        RECT 666.600 206.400 670.200 207.000 ;
        RECT 671.400 206.400 674.400 207.000 ;
        RECT 667.200 205.800 674.400 206.400 ;
        RECT 667.200 205.200 673.800 205.800 ;
        RECT 667.800 204.600 673.800 205.200 ;
        RECT 668.400 204.000 673.200 204.600 ;
        RECT 669.600 203.400 673.200 204.000 ;
        RECT 670.200 202.800 672.600 203.400 ;
        RECT 585.600 196.800 588.600 202.800 ;
        RECT 670.800 202.200 672.000 202.800 ;
        RECT 223.800 194.400 226.800 196.800 ;
        RECT 329.400 195.600 333.600 196.800 ;
        RECT 371.400 196.200 373.800 196.800 ;
        RECT 375.000 196.200 391.800 196.800 ;
        RECT 415.200 196.200 421.200 196.800 ;
        RECT 531.600 196.200 534.000 196.800 ;
        RECT 372.000 195.600 373.200 196.200 ;
        RECT 378.600 195.600 384.000 196.200 ;
        RECT 415.800 195.600 421.800 196.200 ;
        RECT 329.400 195.000 334.200 195.600 ;
        RECT 416.400 195.000 423.000 195.600 ;
        RECT 328.800 194.400 334.800 195.000 ;
        RECT 416.400 194.400 423.600 195.000 ;
        RECT 223.800 193.800 226.200 194.400 ;
        RECT 223.200 192.000 226.200 193.800 ;
        RECT 328.800 193.800 335.400 194.400 ;
        RECT 405.000 193.800 411.600 194.400 ;
        RECT 415.800 193.800 424.800 194.400 ;
        RECT 328.800 193.200 336.000 193.800 ;
        RECT 328.800 192.600 336.600 193.200 ;
        RECT 403.800 192.600 418.800 193.800 ;
        RECT 420.600 193.200 425.400 193.800 ;
        RECT 420.600 192.600 426.000 193.200 ;
        RECT 223.800 190.800 225.600 192.000 ;
        RECT 328.200 190.800 331.200 192.600 ;
        RECT 333.000 192.000 337.200 192.600 ;
        RECT 404.400 192.000 426.600 192.600 ;
        RECT 531.000 192.000 534.000 196.200 ;
        RECT 586.200 195.600 588.600 196.800 ;
        RECT 333.600 191.400 337.800 192.000 ;
        RECT 405.600 191.400 426.600 192.000 ;
        RECT 334.200 190.800 338.400 191.400 ;
        RECT 411.000 190.800 427.200 191.400 ;
        RECT 327.600 190.200 331.200 190.800 ;
        RECT 334.800 190.200 339.600 190.800 ;
        RECT 414.000 190.200 430.200 190.800 ;
        RECT 327.600 189.000 330.600 190.200 ;
        RECT 335.400 189.600 340.200 190.200 ;
        RECT 418.200 189.600 432.600 190.200 ;
        RECT 336.000 189.000 340.800 189.600 ;
        RECT 421.200 189.000 435.000 189.600 ;
        RECT 530.400 189.000 533.400 192.000 ;
        RECT 327.000 188.400 330.600 189.000 ;
        RECT 337.200 188.400 342.000 189.000 ;
        RECT 423.600 188.400 437.400 189.000 ;
        RECT 327.000 186.600 330.000 188.400 ;
        RECT 337.800 187.800 342.600 188.400 ;
        RECT 426.600 187.800 439.800 188.400 ;
        RECT 338.400 187.200 343.800 187.800 ;
        RECT 429.000 187.200 442.200 187.800 ;
        RECT 339.000 186.600 344.400 187.200 ;
        RECT 432.000 186.600 444.000 187.200 ;
        RECT 326.400 185.400 329.400 186.600 ;
        RECT 340.200 186.000 345.600 186.600 ;
        RECT 434.400 186.000 445.800 186.600 ;
        RECT 529.800 186.000 532.800 189.000 ;
        RECT 586.200 187.200 589.200 195.600 ;
        RECT 340.800 185.400 346.800 186.000 ;
        RECT 437.400 185.400 448.200 186.000 ;
        RECT 325.800 184.800 329.400 185.400 ;
        RECT 342.000 184.800 347.400 185.400 ;
        RECT 439.800 184.800 449.400 185.400 ;
        RECT 325.800 183.600 328.800 184.800 ;
        RECT 342.600 184.200 348.600 184.800 ;
        RECT 442.200 184.200 451.200 184.800 ;
        RECT 343.800 183.600 349.800 184.200 ;
        RECT 444.000 183.600 453.000 184.200 ;
        RECT 529.200 183.600 532.200 186.000 ;
        RECT 586.200 185.400 588.600 187.200 ;
        RECT 325.200 183.000 328.800 183.600 ;
        RECT 345.000 183.000 351.000 183.600 ;
        RECT 445.800 183.000 454.800 183.600 ;
        RECT 325.200 181.800 328.200 183.000 ;
        RECT 346.200 182.400 352.200 183.000 ;
        RECT 447.600 182.400 456.600 183.000 ;
        RECT 347.400 181.800 353.400 182.400 ;
        RECT 449.400 181.800 457.800 182.400 ;
        RECT 528.600 181.800 531.600 183.600 ;
        RECT 324.600 180.600 327.600 181.800 ;
        RECT 348.600 181.200 356.400 181.800 ;
        RECT 450.600 181.200 459.000 181.800 ;
        RECT 349.800 180.600 357.000 181.200 ;
        RECT 452.400 180.600 460.200 181.200 ;
        RECT 182.400 178.800 184.800 180.600 ;
        RECT 324.000 180.000 327.600 180.600 ;
        RECT 352.200 180.000 357.000 180.600 ;
        RECT 454.200 180.000 461.400 180.600 ;
        RECT 528.000 180.000 531.000 181.800 ;
        RECT 324.000 178.800 327.000 180.000 ;
        RECT 182.400 171.000 185.400 178.800 ;
        RECT 323.400 177.600 326.400 178.800 ;
        RECT 354.600 177.600 357.600 180.000 ;
        RECT 455.400 179.400 462.000 180.000 ;
        RECT 527.400 179.400 531.000 180.000 ;
        RECT 585.600 180.000 588.600 185.400 ;
        RECT 585.600 179.400 588.000 180.000 ;
        RECT 457.200 178.800 463.200 179.400 ;
        RECT 458.400 178.200 463.800 178.800 ;
        RECT 527.400 178.200 530.400 179.400 ;
        RECT 459.600 177.600 464.400 178.200 ;
        RECT 526.800 177.600 530.400 178.200 ;
        RECT 322.800 177.000 326.400 177.600 ;
        RECT 322.800 176.400 325.800 177.000 ;
        RECT 322.200 175.800 325.800 176.400 ;
        RECT 322.200 174.600 325.200 175.800 ;
        RECT 355.200 174.600 358.200 177.600 ;
        RECT 460.800 177.000 465.000 177.600 ;
        RECT 461.400 176.400 465.600 177.000 ;
        RECT 526.800 176.400 529.800 177.600 ;
        RECT 462.000 175.800 466.200 176.400 ;
        RECT 462.600 175.200 466.800 175.800 ;
        RECT 526.200 175.200 529.200 176.400 ;
        RECT 585.000 175.800 588.000 179.400 ;
        RECT 463.200 174.600 467.400 175.200 ;
        RECT 525.600 174.600 529.200 175.200 ;
        RECT 584.400 175.200 588.000 175.800 ;
        RECT 321.600 173.400 324.600 174.600 ;
        RECT 321.000 172.800 324.600 173.400 ;
        RECT 321.000 172.200 324.000 172.800 ;
        RECT 355.800 172.200 358.800 174.600 ;
        RECT 463.800 174.000 468.000 174.600 ;
        RECT 464.400 173.400 468.600 174.000 ;
        RECT 525.600 173.400 528.600 174.600 ;
        RECT 465.000 172.800 468.600 173.400 ;
        RECT 465.600 172.200 469.200 172.800 ;
        RECT 525.000 172.200 528.000 173.400 ;
        RECT 584.400 172.800 587.400 175.200 ;
        RECT 320.400 171.600 324.000 172.200 ;
        RECT 320.400 171.000 323.400 171.600 ;
        RECT 183.000 169.800 185.400 171.000 ;
        RECT 319.800 170.400 323.400 171.000 ;
        RECT 356.400 170.400 359.400 172.200 ;
        RECT 466.200 171.000 469.800 172.200 ;
        RECT 524.400 171.600 528.000 172.200 ;
        RECT 583.800 172.200 587.400 172.800 ;
        RECT 524.400 171.000 527.400 171.600 ;
        RECT 466.800 170.400 470.400 171.000 ;
        RECT 319.800 169.800 322.800 170.400 ;
        RECT 183.000 164.400 186.000 169.800 ;
        RECT 319.200 169.200 322.800 169.800 ;
        RECT 357.000 169.200 360.000 170.400 ;
        RECT 467.400 169.800 470.400 170.400 ;
        RECT 523.800 170.400 527.400 171.000 ;
        RECT 583.800 170.400 586.800 172.200 ;
        RECT 523.800 169.800 526.800 170.400 ;
        RECT 467.400 169.200 471.000 169.800 ;
        RECT 318.600 168.600 322.200 169.200 ;
        RECT 357.000 168.600 360.600 169.200 ;
        RECT 318.600 168.000 321.600 168.600 ;
        RECT 318.000 167.400 321.600 168.000 ;
        RECT 357.600 168.000 360.600 168.600 ;
        RECT 468.000 168.000 471.000 169.200 ;
        RECT 523.200 169.200 526.800 169.800 ;
        RECT 583.200 169.800 586.800 170.400 ;
        RECT 523.200 168.600 526.200 169.200 ;
        RECT 583.200 168.600 586.200 169.800 ;
        RECT 522.600 168.000 526.200 168.600 ;
        RECT 582.600 168.000 586.200 168.600 ;
        RECT 357.600 167.400 361.200 168.000 ;
        RECT 465.600 167.400 471.600 168.000 ;
        RECT 522.600 167.400 525.600 168.000 ;
        RECT 318.000 166.800 321.000 167.400 ;
        RECT 317.400 166.200 321.000 166.800 ;
        RECT 358.200 166.800 361.200 167.400 ;
        RECT 453.600 166.800 456.600 167.400 ;
        RECT 358.200 166.200 361.800 166.800 ;
        RECT 317.400 165.600 320.400 166.200 ;
        RECT 316.800 165.000 320.400 165.600 ;
        RECT 358.800 165.600 361.800 166.200 ;
        RECT 453.600 166.200 459.000 166.800 ;
        RECT 464.400 166.200 471.600 167.400 ;
        RECT 522.000 166.800 525.600 167.400 ;
        RECT 453.600 165.600 460.800 166.200 ;
        RECT 358.800 165.000 362.400 165.600 ;
        RECT 453.600 165.000 462.000 165.600 ;
        RECT 463.800 165.000 471.600 166.200 ;
        RECT 521.400 166.200 525.000 166.800 ;
        RECT 582.600 166.200 585.600 168.000 ;
        RECT 521.400 165.600 524.400 166.200 ;
        RECT 183.600 163.800 186.000 164.400 ;
        RECT 316.200 163.800 319.800 165.000 ;
        RECT 359.400 164.400 363.000 165.000 ;
        RECT 454.800 164.400 471.600 165.000 ;
        RECT 520.800 165.000 524.400 165.600 ;
        RECT 582.000 165.600 585.600 166.200 ;
        RECT 582.000 165.000 585.000 165.600 ;
        RECT 520.800 164.400 523.800 165.000 ;
        RECT 359.400 163.800 363.600 164.400 ;
        RECT 456.600 163.800 466.800 164.400 ;
        RECT 468.000 163.800 471.600 164.400 ;
        RECT 520.200 163.800 523.800 164.400 ;
        RECT 581.400 163.800 585.000 165.000 ;
        RECT 183.600 159.000 186.600 163.800 ;
        RECT 315.600 163.200 320.400 163.800 ;
        RECT 360.000 163.200 364.200 163.800 ;
        RECT 459.000 163.200 466.800 163.800 ;
        RECT 468.600 163.200 472.200 163.800 ;
        RECT 519.600 163.200 523.200 163.800 ;
        RECT 581.400 163.200 584.400 163.800 ;
        RECT 315.000 162.600 321.000 163.200 ;
        RECT 360.600 162.600 364.800 163.200 ;
        RECT 460.200 162.600 466.800 163.200 ;
        RECT 469.200 162.600 472.800 163.200 ;
        RECT 519.600 162.600 522.600 163.200 ;
        RECT 315.000 162.000 321.600 162.600 ;
        RECT 361.200 162.000 365.400 162.600 ;
        RECT 461.400 162.000 466.800 162.600 ;
        RECT 314.400 161.400 322.200 162.000 ;
        RECT 361.800 161.400 366.600 162.000 ;
        RECT 462.000 161.400 466.800 162.000 ;
        RECT 469.800 162.000 472.800 162.600 ;
        RECT 519.000 162.000 522.600 162.600 ;
        RECT 580.800 162.000 584.400 163.200 ;
        RECT 469.800 161.400 473.400 162.000 ;
        RECT 313.800 160.200 317.400 161.400 ;
        RECT 318.600 160.800 322.800 161.400 ;
        RECT 362.400 160.800 367.200 161.400 ;
        RECT 463.200 160.800 467.400 161.400 ;
        RECT 319.200 160.200 323.400 160.800 ;
        RECT 363.000 160.200 368.400 160.800 ;
        RECT 463.800 160.200 467.400 160.800 ;
        RECT 470.400 160.800 473.400 161.400 ;
        RECT 518.400 161.400 522.000 162.000 ;
        RECT 580.800 161.400 583.800 162.000 ;
        RECT 518.400 160.800 521.400 161.400 ;
        RECT 470.400 160.200 474.000 160.800 ;
        RECT 517.800 160.200 521.400 160.800 ;
        RECT 580.200 160.800 583.800 161.400 ;
        RECT 313.200 159.600 316.800 160.200 ;
        RECT 319.800 159.600 324.000 160.200 ;
        RECT 363.600 159.600 369.600 160.200 ;
        RECT 184.200 158.400 186.600 159.000 ;
        RECT 312.600 158.400 316.200 159.600 ;
        RECT 320.400 159.000 324.600 159.600 ;
        RECT 364.800 159.000 370.800 159.600 ;
        RECT 464.400 159.000 468.000 160.200 ;
        RECT 471.000 159.000 474.000 160.200 ;
        RECT 517.200 159.600 520.800 160.200 ;
        RECT 580.200 159.600 583.200 160.800 ;
        RECT 321.000 158.400 325.200 159.000 ;
        RECT 365.400 158.400 372.600 159.000 ;
        RECT 465.000 158.400 468.600 159.000 ;
        RECT 184.200 154.200 187.200 158.400 ;
        RECT 312.000 157.800 315.600 158.400 ;
        RECT 321.600 157.800 325.800 158.400 ;
        RECT 366.600 157.800 374.400 158.400 ;
        RECT 465.600 157.800 468.600 158.400 ;
        RECT 311.400 157.200 315.000 157.800 ;
        RECT 322.200 157.200 326.400 157.800 ;
        RECT 367.800 157.200 376.800 157.800 ;
        RECT 465.600 157.200 469.200 157.800 ;
        RECT 471.600 157.200 474.600 159.000 ;
        RECT 516.600 158.400 520.200 159.600 ;
        RECT 579.600 159.000 583.200 159.600 ;
        RECT 579.600 158.400 582.600 159.000 ;
        RECT 516.000 157.800 519.600 158.400 ;
        RECT 579.000 157.800 582.600 158.400 ;
        RECT 515.400 157.200 519.000 157.800 ;
        RECT 310.800 156.600 314.400 157.200 ;
        RECT 322.800 156.600 327.600 157.200 ;
        RECT 369.000 156.600 379.200 157.200 ;
        RECT 438.000 156.600 440.400 157.200 ;
        RECT 456.000 156.600 458.400 157.200 ;
        RECT 465.600 156.600 469.800 157.200 ;
        RECT 310.200 156.000 314.400 156.600 ;
        RECT 323.400 156.000 328.200 156.600 ;
        RECT 370.800 156.000 381.600 156.600 ;
        RECT 438.000 156.000 441.600 156.600 ;
        RECT 454.800 156.000 459.600 156.600 ;
        RECT 466.200 156.000 470.400 156.600 ;
        RECT 310.200 155.400 313.800 156.000 ;
        RECT 324.000 155.400 328.800 156.000 ;
        RECT 372.000 155.400 384.600 156.000 ;
        RECT 438.000 155.400 442.200 156.000 ;
        RECT 454.200 155.400 460.200 156.000 ;
        RECT 309.600 154.800 313.200 155.400 ;
        RECT 325.200 154.800 329.400 155.400 ;
        RECT 374.400 154.800 388.200 155.400 ;
        RECT 438.600 154.800 442.800 155.400 ;
        RECT 454.200 154.800 460.800 155.400 ;
        RECT 466.200 154.800 471.000 156.000 ;
        RECT 472.200 154.800 475.200 157.200 ;
        RECT 514.800 156.600 518.400 157.200 ;
        RECT 579.000 156.600 582.000 157.800 ;
        RECT 514.200 156.000 518.400 156.600 ;
        RECT 578.400 156.000 582.000 156.600 ;
        RECT 513.600 155.400 517.800 156.000 ;
        RECT 513.600 154.800 517.200 155.400 ;
        RECT 578.400 154.800 581.400 156.000 ;
        RECT 309.000 154.200 312.600 154.800 ;
        RECT 325.800 154.200 330.000 154.800 ;
        RECT 376.200 154.200 393.000 154.800 ;
        RECT 439.200 154.200 444.000 154.800 ;
        RECT 454.200 154.200 461.400 154.800 ;
        RECT 466.200 154.200 475.200 154.800 ;
        RECT 513.000 154.200 516.600 154.800 ;
        RECT 184.800 153.600 187.200 154.200 ;
        RECT 308.400 153.600 312.000 154.200 ;
        RECT 326.400 153.600 330.600 154.200 ;
        RECT 378.600 153.600 397.200 154.200 ;
        RECT 439.800 153.600 444.600 154.200 ;
        RECT 184.800 150.000 187.800 153.600 ;
        RECT 307.800 153.000 311.400 153.600 ;
        RECT 327.000 153.000 331.200 153.600 ;
        RECT 381.600 153.000 399.000 153.600 ;
        RECT 441.000 153.000 444.600 153.600 ;
        RECT 307.200 152.400 311.400 153.000 ;
        RECT 327.600 152.400 332.400 153.000 ;
        RECT 385.200 152.400 400.800 153.000 ;
        RECT 441.600 152.400 445.200 153.000 ;
        RECT 306.600 151.800 310.800 152.400 ;
        RECT 328.200 151.800 333.000 152.400 ;
        RECT 388.800 151.800 402.600 152.400 ;
        RECT 442.200 151.800 445.800 152.400 ;
        RECT 306.000 151.200 310.200 151.800 ;
        RECT 328.800 151.200 333.600 151.800 ;
        RECT 393.600 151.200 404.400 151.800 ;
        RECT 305.400 150.600 309.600 151.200 ;
        RECT 330.000 150.600 334.200 151.200 ;
        RECT 396.600 150.600 405.600 151.200 ;
        RECT 442.800 150.600 446.400 151.800 ;
        RECT 453.600 150.600 456.600 154.200 ;
        RECT 457.800 153.600 462.000 154.200 ;
        RECT 458.400 153.000 462.600 153.600 ;
        RECT 459.000 152.400 462.600 153.000 ;
        RECT 459.600 151.800 463.200 152.400 ;
        RECT 460.200 151.200 463.200 151.800 ;
        RECT 466.200 151.200 475.800 154.200 ;
        RECT 512.400 153.600 516.000 154.200 ;
        RECT 577.800 153.600 580.800 154.800 ;
        RECT 511.800 153.000 515.400 153.600 ;
        RECT 511.200 152.400 515.400 153.000 ;
        RECT 577.200 153.000 580.800 153.600 ;
        RECT 577.200 152.400 580.200 153.000 ;
        RECT 510.600 151.800 514.800 152.400 ;
        RECT 576.600 151.800 580.200 152.400 ;
        RECT 510.000 151.200 514.200 151.800 ;
        RECT 460.200 150.600 463.800 151.200 ;
        RECT 304.200 150.000 309.000 150.600 ;
        RECT 330.600 150.000 335.400 150.600 ;
        RECT 398.400 150.000 408.000 150.600 ;
        RECT 443.400 150.000 447.000 150.600 ;
        RECT 185.400 149.400 187.800 150.000 ;
        RECT 303.600 149.400 308.400 150.000 ;
        RECT 331.200 149.400 336.000 150.000 ;
        RECT 400.800 149.400 409.800 150.000 ;
        RECT 444.000 149.400 447.600 150.000 ;
        RECT 185.400 145.800 188.400 149.400 ;
        RECT 303.000 148.800 307.800 149.400 ;
        RECT 331.800 148.800 336.600 149.400 ;
        RECT 402.000 148.800 411.000 149.400 ;
        RECT 444.600 148.800 447.600 149.400 ;
        RECT 454.200 148.800 457.200 150.600 ;
        RECT 460.800 150.000 463.800 150.600 ;
        RECT 460.800 149.400 464.400 150.000 ;
        RECT 302.400 148.200 306.600 148.800 ;
        RECT 332.400 148.200 337.200 148.800 ;
        RECT 402.000 148.200 412.800 148.800 ;
        RECT 444.600 148.200 448.200 148.800 ;
        RECT 454.200 148.200 457.800 148.800 ;
        RECT 461.400 148.200 464.400 149.400 ;
        RECT 466.200 148.200 469.200 151.200 ;
        RECT 470.400 150.000 475.800 151.200 ;
        RECT 509.400 150.600 513.600 151.200 ;
        RECT 576.600 150.600 579.600 151.800 ;
        RECT 508.800 150.000 513.000 150.600 ;
        RECT 471.000 148.800 475.800 150.000 ;
        RECT 508.200 149.400 512.400 150.000 ;
        RECT 576.000 149.400 579.000 150.600 ;
        RECT 507.600 148.800 511.800 149.400 ;
        RECT 575.400 148.800 579.000 149.400 ;
        RECT 471.000 148.200 475.200 148.800 ;
        RECT 507.000 148.200 511.200 148.800 ;
        RECT 575.400 148.200 578.400 148.800 ;
        RECT 301.200 147.600 306.600 148.200 ;
        RECT 333.600 147.600 338.400 148.200 ;
        RECT 402.600 147.600 414.600 148.200 ;
        RECT 445.200 147.600 448.200 148.200 ;
        RECT 300.600 147.000 306.600 147.600 ;
        RECT 334.200 147.000 339.000 147.600 ;
        RECT 403.200 147.000 415.800 147.600 ;
        RECT 445.200 147.000 448.800 147.600 ;
        RECT 299.400 146.400 306.600 147.000 ;
        RECT 334.800 146.400 339.600 147.000 ;
        RECT 404.400 146.400 417.600 147.000 ;
        RECT 445.800 146.400 448.800 147.000 ;
        RECT 454.800 147.000 457.800 148.200 ;
        RECT 462.000 147.000 469.200 148.200 ;
        RECT 454.800 146.400 458.400 147.000 ;
        RECT 462.000 146.400 468.600 147.000 ;
        RECT 471.600 146.400 475.200 148.200 ;
        RECT 505.800 147.600 510.600 148.200 ;
        RECT 574.800 147.600 578.400 148.200 ;
        RECT 505.200 147.000 510.000 147.600 ;
        RECT 574.800 147.000 577.800 147.600 ;
        RECT 504.600 146.400 509.400 147.000 ;
        RECT 574.200 146.400 577.800 147.000 ;
        RECT 298.800 145.800 306.600 146.400 ;
        RECT 336.000 145.800 340.800 146.400 ;
        RECT 405.000 145.800 418.800 146.400 ;
        RECT 438.000 145.800 439.200 146.400 ;
        RECT 445.800 145.800 449.400 146.400 ;
        RECT 186.000 145.200 188.400 145.800 ;
        RECT 186.000 142.200 189.000 145.200 ;
        RECT 297.600 144.600 306.000 145.800 ;
        RECT 336.600 145.200 341.400 145.800 ;
        RECT 405.600 145.200 419.400 145.800 ;
        RECT 436.200 145.200 441.000 145.800 ;
        RECT 446.400 145.200 449.400 145.800 ;
        RECT 455.400 145.800 458.400 146.400 ;
        RECT 462.600 145.800 468.600 146.400 ;
        RECT 472.200 145.800 474.600 146.400 ;
        RECT 504.000 145.800 508.200 146.400 ;
        RECT 455.400 145.200 459.000 145.800 ;
        RECT 337.200 144.600 342.000 145.200 ;
        RECT 406.800 144.600 412.800 145.200 ;
        RECT 414.000 144.600 420.000 145.200 ;
        RECT 435.600 144.600 441.600 145.200 ;
        RECT 446.400 144.600 450.000 145.200 ;
        RECT 297.000 144.000 301.200 144.600 ;
        RECT 297.000 143.400 300.000 144.000 ;
        RECT 303.000 142.800 306.000 144.600 ;
        RECT 337.800 144.000 343.200 144.600 ;
        RECT 407.400 144.000 412.800 144.600 ;
        RECT 415.200 144.000 420.600 144.600 ;
        RECT 435.000 144.000 442.200 144.600 ;
        RECT 339.000 143.400 343.800 144.000 ;
        RECT 408.600 143.400 413.400 144.000 ;
        RECT 416.400 143.400 420.600 144.000 ;
        RECT 434.400 143.400 442.800 144.000 ;
        RECT 447.000 143.400 450.000 144.600 ;
        RECT 456.000 144.600 459.000 145.200 ;
        RECT 462.600 145.200 468.000 145.800 ;
        RECT 472.800 145.200 474.000 145.800 ;
        RECT 503.400 145.200 507.600 145.800 ;
        RECT 574.200 145.200 577.200 146.400 ;
        RECT 456.000 144.000 459.600 144.600 ;
        RECT 456.600 143.400 459.600 144.000 ;
        RECT 462.600 144.000 467.400 145.200 ;
        RECT 502.200 144.600 507.000 145.200 ;
        RECT 501.600 144.000 506.400 144.600 ;
        RECT 573.600 144.000 576.600 145.200 ;
        RECT 462.600 143.400 466.800 144.000 ;
        RECT 501.000 143.400 505.800 144.000 ;
        RECT 573.000 143.400 576.600 144.000 ;
        RECT 339.600 142.800 345.000 143.400 ;
        RECT 409.200 142.800 414.600 143.400 ;
        RECT 186.600 141.600 189.000 142.200 ;
        RECT 186.600 138.600 189.600 141.600 ;
        RECT 302.400 141.000 305.400 142.800 ;
        RECT 340.800 142.200 345.600 142.800 ;
        RECT 410.400 142.200 415.200 142.800 ;
        RECT 417.600 142.200 421.200 143.400 ;
        RECT 434.400 142.800 443.400 143.400 ;
        RECT 433.800 142.200 437.400 142.800 ;
        RECT 341.400 141.600 346.800 142.200 ;
        RECT 411.000 141.600 415.800 142.200 ;
        RECT 418.200 141.600 421.800 142.200 ;
        RECT 342.000 141.000 347.400 141.600 ;
        RECT 411.600 141.000 417.000 141.600 ;
        RECT 418.800 141.000 421.800 141.600 ;
        RECT 301.800 140.400 305.400 141.000 ;
        RECT 343.200 140.400 348.600 141.000 ;
        RECT 412.800 140.400 417.600 141.000 ;
        RECT 418.800 140.400 422.400 141.000 ;
        RECT 301.800 138.600 304.800 140.400 ;
        RECT 343.800 139.800 349.200 140.400 ;
        RECT 413.400 139.800 423.000 140.400 ;
        RECT 345.000 139.200 350.400 139.800 ;
        RECT 414.600 139.200 423.000 139.800 ;
        RECT 345.600 138.600 351.600 139.200 ;
        RECT 415.200 138.600 423.600 139.200 ;
        RECT 187.200 135.000 190.200 138.600 ;
        RECT 301.200 136.800 304.200 138.600 ;
        RECT 346.800 138.000 352.200 138.600 ;
        RECT 415.800 138.000 424.200 138.600 ;
        RECT 433.800 138.000 436.800 142.200 ;
        RECT 440.400 141.600 444.000 142.800 ;
        RECT 447.600 141.600 450.600 143.400 ;
        RECT 456.600 142.800 460.200 143.400 ;
        RECT 457.200 142.200 460.800 142.800 ;
        RECT 462.600 142.200 466.200 143.400 ;
        RECT 499.800 142.800 504.600 143.400 ;
        RECT 573.000 142.800 576.000 143.400 ;
        RECT 499.200 142.200 504.000 142.800 ;
        RECT 572.400 142.200 576.000 142.800 ;
        RECT 457.200 141.600 461.400 142.200 ;
        RECT 441.000 141.000 444.000 141.600 ;
        RECT 448.200 141.000 452.400 141.600 ;
        RECT 457.800 141.000 461.400 141.600 ;
        RECT 441.600 139.200 444.600 141.000 ;
        RECT 448.200 140.400 453.600 141.000 ;
        RECT 457.800 140.400 462.000 141.000 ;
        RECT 448.200 139.800 462.000 140.400 ;
        RECT 463.200 139.800 465.600 142.200 ;
        RECT 498.000 141.600 503.400 142.200 ;
        RECT 572.400 141.600 575.400 142.200 ;
        RECT 497.400 141.000 502.200 141.600 ;
        RECT 571.800 141.000 575.400 141.600 ;
        RECT 496.200 140.400 501.600 141.000 ;
        RECT 571.800 140.400 574.800 141.000 ;
        RECT 495.600 139.800 501.000 140.400 ;
        RECT 571.200 139.800 574.800 140.400 ;
        RECT 448.200 139.200 465.600 139.800 ;
        RECT 494.400 139.200 499.800 139.800 ;
        RECT 571.200 139.200 574.200 139.800 ;
        RECT 348.000 137.400 353.400 138.000 ;
        RECT 416.400 137.400 424.200 138.000 ;
        RECT 348.600 136.800 354.600 137.400 ;
        RECT 417.600 136.800 424.800 137.400 ;
        RECT 434.400 136.800 437.400 138.000 ;
        RECT 442.200 136.800 445.200 139.200 ;
        RECT 448.800 138.000 465.600 139.200 ;
        RECT 493.800 138.600 499.200 139.200 ;
        RECT 570.600 138.600 574.200 139.200 ;
        RECT 492.600 138.000 498.000 138.600 ;
        RECT 570.600 138.000 573.600 138.600 ;
        RECT 448.800 136.800 451.800 138.000 ;
        RECT 453.600 137.400 458.400 138.000 ;
        RECT 300.600 135.000 303.600 136.800 ;
        RECT 349.800 136.200 355.200 136.800 ;
        RECT 418.200 136.200 425.400 136.800 ;
        RECT 434.400 136.200 438.000 136.800 ;
        RECT 350.400 135.600 356.400 136.200 ;
        RECT 418.800 135.600 426.000 136.200 ;
        RECT 435.000 135.600 438.000 136.200 ;
        RECT 442.800 136.200 445.200 136.800 ;
        RECT 448.200 136.200 451.800 136.800 ;
        RECT 460.200 136.200 465.600 138.000 ;
        RECT 491.400 137.400 497.400 138.000 ;
        RECT 570.000 137.400 573.600 138.000 ;
        RECT 490.800 136.800 496.200 137.400 ;
        RECT 570.000 136.800 573.000 137.400 ;
        RECT 489.600 136.200 495.000 136.800 ;
        RECT 569.400 136.200 573.000 136.800 ;
        RECT 351.600 135.000 357.600 135.600 ;
        RECT 419.400 135.000 426.600 135.600 ;
        RECT 435.000 135.000 438.600 135.600 ;
        RECT 187.800 132.000 190.800 135.000 ;
        RECT 263.400 134.400 264.000 135.000 ;
        RECT 262.800 133.800 264.600 134.400 ;
        RECT 262.800 132.600 265.200 133.800 ;
        RECT 300.000 133.200 303.000 135.000 ;
        RECT 352.800 134.400 358.800 135.000 ;
        RECT 420.000 134.400 427.200 135.000 ;
        RECT 435.600 134.400 438.600 135.000 ;
        RECT 442.800 134.400 445.800 136.200 ;
        RECT 448.200 135.600 451.200 136.200 ;
        RECT 447.600 135.000 451.200 135.600 ;
        RECT 447.000 134.400 450.600 135.000 ;
        RECT 460.800 134.400 465.600 136.200 ;
        RECT 488.400 135.600 494.400 136.200 ;
        RECT 569.400 135.600 572.400 136.200 ;
        RECT 487.200 135.000 493.200 135.600 ;
        RECT 568.800 135.000 572.400 135.600 ;
        RECT 486.000 134.400 492.000 135.000 ;
        RECT 568.800 134.400 571.800 135.000 ;
        RECT 354.000 133.800 360.000 134.400 ;
        RECT 420.600 133.800 427.800 134.400 ;
        RECT 435.600 133.800 439.200 134.400 ;
        RECT 354.600 133.200 361.200 133.800 ;
        RECT 421.800 133.200 429.000 133.800 ;
        RECT 436.200 133.200 439.800 133.800 ;
        RECT 442.800 133.200 450.000 134.400 ;
        RECT 188.400 129.000 191.400 132.000 ;
        RECT 262.800 131.400 265.800 132.600 ;
        RECT 299.400 131.400 302.400 133.200 ;
        RECT 355.800 132.600 362.400 133.200 ;
        RECT 422.400 132.600 430.800 133.200 ;
        RECT 436.200 132.600 440.400 133.200 ;
        RECT 357.000 132.000 363.600 132.600 ;
        RECT 423.000 132.000 440.400 132.600 ;
        RECT 442.800 132.600 449.400 133.200 ;
        RECT 461.400 132.600 465.600 134.400 ;
        RECT 484.800 133.800 491.400 134.400 ;
        RECT 568.200 133.800 571.800 134.400 ;
        RECT 483.600 133.200 490.200 133.800 ;
        RECT 568.200 133.200 571.200 133.800 ;
        RECT 482.400 132.600 489.000 133.200 ;
        RECT 567.600 132.600 571.200 133.200 ;
        RECT 442.800 132.000 448.800 132.600 ;
        RECT 462.000 132.000 465.600 132.600 ;
        RECT 481.200 132.000 487.800 132.600 ;
        RECT 567.000 132.000 570.600 132.600 ;
        RECT 358.200 131.400 364.800 132.000 ;
        RECT 423.600 131.400 441.000 132.000 ;
        RECT 442.800 131.400 447.600 132.000 ;
        RECT 462.000 131.400 465.000 132.000 ;
        RECT 479.400 131.400 486.600 132.000 ;
        RECT 567.000 131.400 570.000 132.000 ;
        RECT 263.400 130.200 266.400 131.400 ;
        RECT 298.800 130.200 301.800 131.400 ;
        RECT 359.400 130.800 366.000 131.400 ;
        RECT 424.200 130.800 441.600 131.400 ;
        RECT 442.800 130.800 447.000 131.400 ;
        RECT 462.600 130.800 465.000 131.400 ;
        RECT 478.200 130.800 485.400 131.400 ;
        RECT 566.400 130.800 570.000 131.400 ;
        RECT 360.600 130.200 367.200 130.800 ;
        RECT 424.800 130.200 445.800 130.800 ;
        RECT 477.000 130.200 484.200 130.800 ;
        RECT 566.400 130.200 569.400 130.800 ;
        RECT 264.000 129.600 267.000 130.200 ;
        RECT 298.200 129.600 301.800 130.200 ;
        RECT 361.800 129.600 369.000 130.200 ;
        RECT 425.400 129.600 436.800 130.200 ;
        RECT 438.600 129.600 445.800 130.200 ;
        RECT 475.200 129.600 483.000 130.200 ;
        RECT 565.800 129.600 569.400 130.200 ;
        RECT 264.000 129.000 267.600 129.600 ;
        RECT 189.000 126.000 192.000 129.000 ;
        RECT 264.600 128.400 267.600 129.000 ;
        RECT 298.200 128.400 301.200 129.600 ;
        RECT 363.000 129.000 370.200 129.600 ;
        RECT 426.000 129.000 430.200 129.600 ;
        RECT 364.200 128.400 371.400 129.000 ;
        RECT 426.600 128.400 430.200 129.000 ;
        RECT 439.200 128.400 445.800 129.600 ;
        RECT 474.000 129.000 481.200 129.600 ;
        RECT 565.800 129.000 568.800 129.600 ;
        RECT 472.200 128.400 480.000 129.000 ;
        RECT 565.200 128.400 568.800 129.000 ;
        RECT 264.600 127.200 268.200 128.400 ;
        RECT 297.600 127.200 300.600 128.400 ;
        RECT 365.400 127.800 373.200 128.400 ;
        RECT 367.200 127.200 375.000 127.800 ;
        RECT 427.200 127.200 430.800 128.400 ;
        RECT 439.800 127.200 445.800 128.400 ;
        RECT 470.400 127.800 478.800 128.400 ;
        RECT 468.600 127.200 477.000 127.800 ;
        RECT 564.600 127.200 568.200 128.400 ;
        RECT 265.200 126.600 268.800 127.200 ;
        RECT 265.800 126.000 268.800 126.600 ;
        RECT 297.000 126.600 300.600 127.200 ;
        RECT 368.400 126.600 376.200 127.200 ;
        RECT 427.800 126.600 431.400 127.200 ;
        RECT 439.800 126.600 445.200 127.200 ;
        RECT 467.400 126.600 475.800 127.200 ;
        RECT 564.000 126.600 567.600 127.200 ;
        RECT 189.600 123.600 192.600 126.000 ;
        RECT 265.800 125.400 269.400 126.000 ;
        RECT 297.000 125.400 300.000 126.600 ;
        RECT 369.600 126.000 378.000 126.600 ;
        RECT 428.400 126.000 431.400 126.600 ;
        RECT 371.400 125.400 379.800 126.000 ;
        RECT 266.400 124.800 269.400 125.400 ;
        RECT 247.800 124.200 249.600 124.800 ;
        RECT 266.400 124.200 270.000 124.800 ;
        RECT 296.400 124.200 299.400 125.400 ;
        RECT 372.600 124.800 381.600 125.400 ;
        RECT 428.400 124.800 432.000 126.000 ;
        RECT 374.400 124.200 384.000 124.800 ;
        RECT 429.000 124.200 432.000 124.800 ;
        RECT 440.400 125.400 445.200 126.600 ;
        RECT 465.600 126.000 474.000 126.600 ;
        RECT 564.000 126.000 567.000 126.600 ;
        RECT 463.200 125.400 472.800 126.000 ;
        RECT 563.400 125.400 567.000 126.000 ;
        RECT 440.400 124.200 444.600 125.400 ;
        RECT 461.400 124.800 471.000 125.400 ;
        RECT 459.000 124.200 469.200 124.800 ;
        RECT 562.800 124.200 566.400 125.400 ;
        RECT 190.200 120.600 193.200 123.600 ;
        RECT 247.200 120.600 250.200 124.200 ;
        RECT 267.000 123.000 270.600 124.200 ;
        RECT 295.800 123.600 299.400 124.200 ;
        RECT 376.200 123.600 385.800 124.200 ;
        RECT 295.800 123.000 298.800 123.600 ;
        RECT 378.000 123.000 388.200 123.600 ;
        RECT 267.600 121.800 271.200 123.000 ;
        RECT 295.200 122.400 298.800 123.000 ;
        RECT 379.800 122.400 391.200 123.000 ;
        RECT 429.000 122.400 432.600 124.200 ;
        RECT 441.000 123.600 444.600 124.200 ;
        RECT 456.600 123.600 467.400 124.200 ;
        RECT 562.200 123.600 565.800 124.200 ;
        RECT 441.600 123.000 444.000 123.600 ;
        RECT 453.600 123.000 465.600 123.600 ;
        RECT 562.200 123.000 565.200 123.600 ;
        RECT 441.600 122.400 443.400 123.000 ;
        RECT 450.600 122.400 463.200 123.000 ;
        RECT 561.600 122.400 565.200 123.000 ;
        RECT 268.200 121.200 271.800 121.800 ;
        RECT 295.200 121.200 298.200 122.400 ;
        RECT 381.600 121.800 393.600 122.400 ;
        RECT 384.000 121.200 396.600 121.800 ;
        RECT 429.600 121.200 432.600 122.400 ;
        RECT 447.600 121.800 461.400 122.400 ;
        RECT 561.000 121.800 564.600 122.400 ;
        RECT 444.000 121.200 459.000 121.800 ;
        RECT 561.000 121.200 564.000 121.800 ;
        RECT 268.200 120.600 272.400 121.200 ;
        RECT 190.800 118.200 193.800 120.600 ;
        RECT 247.800 118.200 250.800 120.600 ;
        RECT 268.800 120.000 272.400 120.600 ;
        RECT 294.600 120.000 297.600 121.200 ;
        RECT 385.800 120.600 400.800 121.200 ;
        RECT 388.200 120.000 405.000 120.600 ;
        RECT 430.200 120.000 433.200 121.200 ;
        RECT 440.400 120.600 456.600 121.200 ;
        RECT 560.400 120.600 564.000 121.200 ;
        RECT 435.000 120.000 453.600 120.600 ;
        RECT 269.400 118.800 273.000 120.000 ;
        RECT 294.000 118.800 297.000 120.000 ;
        RECT 391.200 119.400 412.800 120.000 ;
        RECT 427.800 119.400 450.600 120.000 ;
        RECT 559.800 119.400 563.400 120.600 ;
        RECT 393.600 118.800 447.600 119.400 ;
        RECT 559.200 118.800 562.800 119.400 ;
        RECT 270.000 118.200 273.600 118.800 ;
        RECT 293.400 118.200 296.400 118.800 ;
        RECT 397.200 118.200 444.000 118.800 ;
        RECT 191.400 115.800 194.400 118.200 ;
        RECT 248.400 117.000 251.400 118.200 ;
        RECT 270.600 117.000 274.200 118.200 ;
        RECT 292.800 117.600 296.400 118.200 ;
        RECT 400.800 117.600 439.800 118.200 ;
        RECT 558.600 117.600 562.200 118.800 ;
        RECT 292.800 117.000 295.800 117.600 ;
        RECT 405.600 117.000 434.400 117.600 ;
        RECT 558.000 117.000 561.600 117.600 ;
        RECT 248.400 116.400 252.000 117.000 ;
        RECT 192.000 113.400 195.000 115.800 ;
        RECT 249.000 115.200 252.000 116.400 ;
        RECT 271.200 116.400 274.800 117.000 ;
        RECT 292.200 116.400 295.800 117.000 ;
        RECT 414.000 116.400 426.000 117.000 ;
        RECT 557.400 116.400 561.000 117.000 ;
        RECT 271.200 115.200 275.400 116.400 ;
        RECT 292.200 115.800 295.200 116.400 ;
        RECT 291.600 115.200 295.200 115.800 ;
        RECT 556.800 115.200 560.400 116.400 ;
        RECT 249.000 114.600 252.600 115.200 ;
        RECT 249.600 114.000 252.600 114.600 ;
        RECT 271.200 114.600 276.000 115.200 ;
        RECT 291.600 114.600 294.600 115.200 ;
        RECT 556.200 114.600 559.800 115.200 ;
        RECT 271.200 114.000 276.600 114.600 ;
        RECT 291.000 114.000 294.600 114.600 ;
        RECT 555.600 114.000 559.200 114.600 ;
        RECT 249.600 113.400 253.200 114.000 ;
        RECT 192.600 111.000 195.600 113.400 ;
        RECT 250.200 112.800 253.200 113.400 ;
        RECT 271.200 112.800 277.200 114.000 ;
        RECT 290.400 113.400 294.000 114.000 ;
        RECT 555.000 113.400 559.200 114.000 ;
        RECT 290.400 112.800 293.400 113.400 ;
        RECT 555.000 112.800 558.600 113.400 ;
        RECT 229.800 112.200 231.000 112.800 ;
        RECT 250.200 112.200 253.800 112.800 ;
        RECT 229.200 111.600 231.600 112.200 ;
        RECT 250.800 111.600 253.800 112.200 ;
        RECT 271.200 112.200 277.800 112.800 ;
        RECT 289.800 112.200 293.400 112.800 ;
        RECT 554.400 112.200 558.000 112.800 ;
        RECT 271.200 111.600 278.400 112.200 ;
        RECT 289.200 111.600 292.800 112.200 ;
        RECT 553.800 111.600 557.400 112.200 ;
        RECT 193.200 109.200 196.200 111.000 ;
        RECT 229.200 110.400 232.200 111.600 ;
        RECT 250.800 111.000 254.400 111.600 ;
        RECT 251.400 110.400 254.400 111.000 ;
        RECT 271.800 111.000 279.000 111.600 ;
        RECT 271.800 110.400 279.600 111.000 ;
        RECT 288.600 110.400 292.200 111.600 ;
        RECT 553.200 111.000 557.400 111.600 ;
        RECT 553.200 110.400 556.800 111.000 ;
        RECT 193.800 107.400 196.800 109.200 ;
        RECT 229.800 108.600 232.800 110.400 ;
        RECT 251.400 109.800 255.000 110.400 ;
        RECT 252.000 109.200 255.000 109.800 ;
        RECT 252.000 108.600 255.600 109.200 ;
        RECT 230.400 107.400 233.400 108.600 ;
        RECT 252.600 108.000 256.200 108.600 ;
        RECT 253.200 107.400 256.200 108.000 ;
        RECT 193.800 106.800 197.400 107.400 ;
        RECT 194.400 105.600 197.400 106.800 ;
        RECT 231.000 106.200 234.000 107.400 ;
        RECT 253.200 106.800 256.800 107.400 ;
        RECT 253.800 106.200 257.400 106.800 ;
        RECT 231.000 105.600 234.600 106.200 ;
        RECT 194.400 105.000 198.000 105.600 ;
        RECT 195.000 104.400 198.000 105.000 ;
        RECT 231.600 105.000 234.600 105.600 ;
        RECT 254.400 105.600 258.000 106.200 ;
        RECT 231.600 104.400 235.200 105.000 ;
        RECT 254.400 104.400 258.600 105.600 ;
        RECT 195.000 103.200 198.600 104.400 ;
        RECT 232.200 103.200 235.800 104.400 ;
        RECT 254.400 103.800 259.200 104.400 ;
        RECT 254.400 103.200 259.800 103.800 ;
        RECT 195.600 102.000 198.600 103.200 ;
        RECT 232.800 102.000 236.400 103.200 ;
        RECT 254.400 102.600 260.400 103.200 ;
        RECT 254.400 102.000 261.600 102.600 ;
        RECT 271.800 102.000 274.800 110.400 ;
        RECT 276.000 109.800 280.200 110.400 ;
        RECT 288.000 109.800 291.600 110.400 ;
        RECT 552.600 109.800 556.200 110.400 ;
        RECT 276.600 109.200 280.800 109.800 ;
        RECT 287.400 109.200 291.000 109.800 ;
        RECT 552.000 109.200 555.600 109.800 ;
        RECT 277.200 108.600 281.400 109.200 ;
        RECT 286.800 108.600 290.400 109.200 ;
        RECT 551.400 108.600 555.000 109.200 ;
        RECT 277.800 108.000 282.000 108.600 ;
        RECT 286.200 108.000 290.400 108.600 ;
        RECT 550.800 108.000 555.000 108.600 ;
        RECT 278.400 107.400 282.600 108.000 ;
        RECT 285.600 107.400 289.800 108.000 ;
        RECT 550.200 107.400 554.400 108.000 ;
        RECT 279.000 106.800 283.200 107.400 ;
        RECT 284.400 106.800 289.200 107.400 ;
        RECT 549.600 106.800 553.800 107.400 ;
        RECT 279.600 106.200 288.600 106.800 ;
        RECT 549.600 106.200 553.200 106.800 ;
        RECT 280.200 105.600 288.000 106.200 ;
        RECT 549.000 105.600 552.600 106.200 ;
        RECT 280.800 105.000 287.400 105.600 ;
        RECT 548.400 105.000 552.000 105.600 ;
        RECT 281.400 104.400 286.800 105.000 ;
        RECT 547.800 104.400 551.400 105.000 ;
        RECT 282.000 103.800 285.600 104.400 ;
        RECT 547.200 103.800 551.400 104.400 ;
        RECT 282.600 103.200 284.400 103.800 ;
        RECT 546.600 103.200 550.800 103.800 ;
        RECT 546.000 102.600 550.200 103.200 ;
        RECT 545.400 102.000 549.600 102.600 ;
        RECT 195.600 100.800 199.200 102.000 ;
        RECT 196.200 100.200 199.200 100.800 ;
        RECT 232.200 100.800 237.000 102.000 ;
        RECT 253.800 101.400 262.200 102.000 ;
        RECT 253.800 100.800 262.800 101.400 ;
        RECT 232.200 100.200 237.600 100.800 ;
        RECT 196.200 99.000 199.800 100.200 ;
        RECT 232.200 99.000 238.200 100.200 ;
        RECT 196.800 98.400 199.800 99.000 ;
        RECT 231.600 98.400 238.800 99.000 ;
        RECT 253.800 98.400 256.800 100.800 ;
        RECT 258.600 100.200 264.000 100.800 ;
        RECT 259.200 99.600 265.200 100.200 ;
        RECT 259.800 99.000 267.600 99.600 ;
        RECT 271.200 99.000 274.800 102.000 ;
        RECT 544.800 101.400 549.000 102.000 ;
        RECT 544.200 100.800 548.400 101.400 ;
        RECT 543.600 100.200 547.800 100.800 ;
        RECT 543.000 99.600 547.200 100.200 ;
        RECT 542.400 99.000 546.600 99.600 ;
        RECT 260.400 98.400 274.200 99.000 ;
        RECT 541.800 98.400 546.000 99.000 ;
        RECT 196.800 97.200 200.400 98.400 ;
        RECT 197.400 96.600 200.400 97.200 ;
        RECT 231.600 96.600 234.600 98.400 ;
        RECT 235.800 97.200 239.400 98.400 ;
        RECT 236.400 96.600 240.000 97.200 ;
        RECT 197.400 96.000 201.000 96.600 ;
        RECT 198.000 95.400 201.000 96.000 ;
        RECT 198.000 94.200 201.600 95.400 ;
        RECT 231.000 94.800 234.000 96.600 ;
        RECT 237.000 96.000 240.600 96.600 ;
        RECT 237.000 95.400 241.200 96.000 ;
        RECT 253.200 95.400 256.200 98.400 ;
        RECT 261.600 97.800 274.200 98.400 ;
        RECT 540.600 97.800 545.400 98.400 ;
        RECT 262.200 97.200 274.200 97.800 ;
        RECT 540.000 97.200 544.800 97.800 ;
        RECT 263.400 96.600 273.600 97.200 ;
        RECT 539.400 96.600 544.200 97.200 ;
        RECT 264.000 96.000 273.000 96.600 ;
        RECT 538.800 96.000 543.000 96.600 ;
        RECT 265.200 95.400 271.800 96.000 ;
        RECT 538.200 95.400 542.400 96.000 ;
        RECT 237.600 94.800 241.200 95.400 ;
        RECT 198.600 93.600 201.600 94.200 ;
        RECT 198.600 92.400 202.200 93.600 ;
        RECT 230.400 93.000 233.400 94.800 ;
        RECT 238.200 94.200 241.800 94.800 ;
        RECT 238.800 93.600 242.400 94.200 ;
        RECT 238.800 93.000 243.000 93.600 ;
        RECT 199.200 91.200 202.800 92.400 ;
        RECT 229.800 91.200 232.800 93.000 ;
        RECT 239.400 92.400 243.600 93.000 ;
        RECT 252.600 92.400 255.600 95.400 ;
        RECT 265.800 94.800 271.800 95.400 ;
        RECT 537.600 94.800 541.800 95.400 ;
        RECT 267.000 94.200 272.400 94.800 ;
        RECT 537.000 94.200 541.200 94.800 ;
        RECT 268.200 93.600 273.600 94.200 ;
        RECT 536.400 93.600 540.600 94.200 ;
        RECT 268.800 93.000 274.800 93.600 ;
        RECT 535.800 93.000 540.000 93.600 ;
        RECT 270.000 92.400 275.400 93.000 ;
        RECT 535.200 92.400 539.400 93.000 ;
        RECT 240.000 91.800 244.200 92.400 ;
        RECT 240.600 91.200 244.200 91.800 ;
        RECT 199.800 90.000 203.400 91.200 ;
        RECT 229.200 90.000 232.200 91.200 ;
        RECT 241.200 90.600 244.800 91.200 ;
        RECT 241.800 90.000 245.400 90.600 ;
        RECT 200.400 89.400 203.400 90.000 ;
        RECT 228.600 89.400 232.200 90.000 ;
        RECT 242.400 89.400 246.000 90.000 ;
        RECT 252.000 89.400 255.000 92.400 ;
        RECT 271.200 91.800 276.600 92.400 ;
        RECT 534.600 91.800 538.800 92.400 ;
        RECT 271.800 91.200 277.800 91.800 ;
        RECT 534.000 91.200 538.200 91.800 ;
        RECT 273.000 90.600 279.000 91.200 ;
        RECT 533.400 90.600 537.600 91.200 ;
        RECT 274.200 90.000 279.600 90.600 ;
        RECT 532.800 90.000 537.000 90.600 ;
        RECT 274.800 89.400 280.800 90.000 ;
        RECT 531.600 89.400 536.400 90.000 ;
        RECT 200.400 88.800 204.000 89.400 ;
        RECT 201.000 88.200 204.000 88.800 ;
        RECT 228.600 88.200 231.600 89.400 ;
        RECT 243.000 88.800 246.600 89.400 ;
        RECT 243.000 88.200 247.800 88.800 ;
        RECT 201.000 87.600 204.600 88.200 ;
        RECT 201.600 87.000 204.600 87.600 ;
        RECT 228.000 87.600 231.600 88.200 ;
        RECT 243.600 87.600 248.400 88.200 ;
        RECT 228.000 87.000 231.000 87.600 ;
        RECT 244.800 87.000 249.000 87.600 ;
        RECT 201.600 86.400 205.200 87.000 ;
        RECT 227.400 86.400 231.000 87.000 ;
        RECT 245.400 86.400 249.600 87.000 ;
        RECT 251.400 86.400 254.400 89.400 ;
        RECT 276.000 88.800 282.000 89.400 ;
        RECT 531.000 88.800 535.800 89.400 ;
        RECT 277.200 88.200 283.200 88.800 ;
        RECT 530.400 88.200 535.200 88.800 ;
        RECT 278.400 87.600 284.400 88.200 ;
        RECT 529.800 87.600 534.000 88.200 ;
        RECT 279.000 87.000 285.000 87.600 ;
        RECT 529.200 87.000 533.400 87.600 ;
        RECT 280.200 86.400 286.200 87.000 ;
        RECT 528.000 86.400 532.800 87.000 ;
        RECT 202.200 85.200 205.800 86.400 ;
        RECT 227.400 85.200 230.400 86.400 ;
        RECT 246.000 85.800 250.200 86.400 ;
        RECT 251.400 85.800 253.800 86.400 ;
        RECT 281.400 85.800 287.400 86.400 ;
        RECT 527.400 85.800 532.200 86.400 ;
        RECT 246.600 85.200 253.800 85.800 ;
        RECT 282.600 85.200 288.600 85.800 ;
        RECT 526.800 85.200 531.600 85.800 ;
        RECT 202.800 84.000 206.400 85.200 ;
        RECT 226.800 84.000 229.800 85.200 ;
        RECT 247.200 84.600 253.800 85.200 ;
        RECT 283.800 84.600 289.800 85.200 ;
        RECT 526.200 84.600 531.000 85.200 ;
        RECT 248.400 84.000 253.800 84.600 ;
        RECT 284.400 84.000 291.000 84.600 ;
        RECT 525.000 84.000 529.800 84.600 ;
        RECT 203.400 82.800 207.000 84.000 ;
        RECT 226.200 83.400 229.800 84.000 ;
        RECT 249.000 83.400 253.800 84.000 ;
        RECT 285.600 83.400 292.200 84.000 ;
        RECT 524.400 83.400 529.200 84.000 ;
        RECT 226.200 82.800 229.200 83.400 ;
        RECT 250.800 82.800 253.800 83.400 ;
        RECT 286.800 82.800 293.400 83.400 ;
        RECT 523.800 82.800 528.600 83.400 ;
        RECT 204.000 82.200 207.600 82.800 ;
        RECT 204.600 81.600 207.600 82.200 ;
        RECT 225.600 82.200 229.200 82.800 ;
        RECT 251.400 82.200 253.200 82.800 ;
        RECT 288.000 82.200 294.600 82.800 ;
        RECT 522.600 82.200 528.000 82.800 ;
        RECT 225.600 81.600 228.600 82.200 ;
        RECT 289.200 81.600 295.800 82.200 ;
        RECT 522.000 81.600 526.800 82.200 ;
        RECT 204.600 81.000 208.200 81.600 ;
        RECT 225.000 81.000 228.600 81.600 ;
        RECT 290.400 81.000 297.000 81.600 ;
        RECT 521.400 81.000 526.200 81.600 ;
        RECT 205.200 80.400 208.800 81.000 ;
        RECT 225.000 80.400 228.000 81.000 ;
        RECT 291.600 80.400 298.200 81.000 ;
        RECT 520.200 80.400 525.600 81.000 ;
        RECT 205.800 79.800 208.800 80.400 ;
        RECT 224.400 79.800 228.000 80.400 ;
        RECT 292.800 79.800 299.400 80.400 ;
        RECT 519.600 79.800 524.400 80.400 ;
        RECT 205.800 79.200 209.400 79.800 ;
        RECT 224.400 79.200 227.400 79.800 ;
        RECT 294.000 79.200 300.600 79.800 ;
        RECT 518.400 79.200 523.800 79.800 ;
        RECT 206.400 78.600 209.400 79.200 ;
        RECT 223.800 78.600 227.400 79.200 ;
        RECT 295.200 78.600 301.800 79.200 ;
        RECT 517.800 78.600 522.600 79.200 ;
        RECT 206.400 78.000 210.000 78.600 ;
        RECT 223.800 78.000 226.800 78.600 ;
        RECT 296.400 78.000 303.600 78.600 ;
        RECT 516.600 78.000 522.000 78.600 ;
        RECT 207.000 77.400 210.600 78.000 ;
        RECT 223.200 77.400 226.800 78.000 ;
        RECT 297.600 77.400 304.800 78.000 ;
        RECT 516.000 77.400 521.400 78.000 ;
        RECT 207.600 76.200 211.200 77.400 ;
        RECT 223.200 76.800 226.200 77.400 ;
        RECT 298.800 76.800 306.000 77.400 ;
        RECT 514.800 76.800 520.200 77.400 ;
        RECT 222.600 76.200 226.200 76.800 ;
        RECT 300.000 76.200 307.200 76.800 ;
        RECT 514.200 76.200 519.600 76.800 ;
        RECT 208.200 75.600 211.800 76.200 ;
        RECT 222.000 75.600 225.600 76.200 ;
        RECT 301.800 75.600 309.000 76.200 ;
        RECT 513.000 75.600 518.400 76.200 ;
        RECT 208.800 75.000 212.400 75.600 ;
        RECT 209.400 74.400 213.000 75.000 ;
        RECT 221.400 74.400 225.000 75.600 ;
        RECT 303.000 75.000 310.200 75.600 ;
        RECT 511.800 75.000 517.800 75.600 ;
        RECT 304.200 74.400 311.400 75.000 ;
        RECT 511.200 74.400 516.600 75.000 ;
        RECT 209.400 73.800 213.600 74.400 ;
        RECT 220.800 73.800 224.400 74.400 ;
        RECT 305.400 73.800 313.200 74.400 ;
        RECT 510.000 73.800 515.400 74.400 ;
        RECT 210.000 73.200 214.200 73.800 ;
        RECT 220.200 73.200 223.800 73.800 ;
        RECT 307.200 73.200 314.400 73.800 ;
        RECT 508.800 73.200 514.800 73.800 ;
        RECT 210.600 72.600 215.400 73.200 ;
        RECT 219.600 72.600 223.800 73.200 ;
        RECT 308.400 72.600 316.200 73.200 ;
        RECT 507.600 72.600 513.600 73.200 ;
        RECT 211.200 72.000 216.000 72.600 ;
        RECT 219.000 72.000 223.200 72.600 ;
        RECT 309.600 72.000 317.400 72.600 ;
        RECT 507.000 72.000 512.400 72.600 ;
        RECT 211.800 71.400 216.600 72.000 ;
        RECT 218.400 71.400 222.600 72.000 ;
        RECT 311.400 71.400 319.200 72.000 ;
        RECT 505.800 71.400 511.800 72.000 ;
        RECT 212.400 70.800 222.000 71.400 ;
        RECT 312.600 70.800 320.400 71.400 ;
        RECT 504.600 70.800 510.600 71.400 ;
        RECT 213.000 70.200 221.400 70.800 ;
        RECT 314.400 70.200 322.200 70.800 ;
        RECT 503.400 70.200 509.400 70.800 ;
        RECT 213.600 69.600 220.800 70.200 ;
        RECT 315.600 69.600 324.000 70.200 ;
        RECT 502.200 69.600 508.200 70.200 ;
        RECT 214.200 69.000 219.600 69.600 ;
        RECT 317.400 69.000 325.800 69.600 ;
        RECT 501.000 69.000 507.000 69.600 ;
        RECT 214.800 68.400 219.000 69.000 ;
        RECT 318.600 68.400 327.000 69.000 ;
        RECT 499.200 68.400 506.400 69.000 ;
        RECT 216.000 67.800 218.400 68.400 ;
        RECT 320.400 67.800 328.800 68.400 ;
        RECT 498.000 67.800 505.200 68.400 ;
        RECT 322.200 67.200 330.600 67.800 ;
        RECT 496.800 67.200 504.000 67.800 ;
        RECT 323.400 66.600 332.400 67.200 ;
        RECT 495.600 66.600 502.800 67.200 ;
        RECT 325.200 66.000 334.200 66.600 ;
        RECT 493.800 66.000 501.000 66.600 ;
        RECT 327.000 65.400 336.600 66.000 ;
        RECT 492.600 65.400 499.800 66.000 ;
        RECT 328.800 64.800 338.400 65.400 ;
        RECT 490.800 64.800 498.600 65.400 ;
        RECT 330.600 64.200 340.200 64.800 ;
        RECT 489.000 64.200 497.400 64.800 ;
        RECT 332.400 63.600 342.600 64.200 ;
        RECT 487.200 63.600 495.600 64.200 ;
        RECT 334.200 63.000 344.400 63.600 ;
        RECT 485.400 63.000 494.400 63.600 ;
        RECT 336.000 62.400 346.800 63.000 ;
        RECT 483.600 62.400 492.600 63.000 ;
        RECT 338.400 61.800 349.200 62.400 ;
        RECT 481.800 61.800 491.400 62.400 ;
        RECT 340.200 61.200 351.600 61.800 ;
        RECT 479.400 61.200 491.400 61.800 ;
        RECT 342.000 60.600 354.000 61.200 ;
        RECT 477.600 60.600 491.400 61.200 ;
        RECT 344.400 60.000 356.400 60.600 ;
        RECT 474.600 60.000 493.200 60.600 ;
        RECT 346.800 59.400 359.400 60.000 ;
        RECT 472.200 59.400 484.200 60.000 ;
        RECT 487.200 59.400 495.600 60.000 ;
        RECT 349.200 58.800 362.400 59.400 ;
        RECT 469.200 58.800 481.800 59.400 ;
        RECT 488.400 58.800 499.800 59.400 ;
        RECT 351.600 58.200 365.400 58.800 ;
        RECT 465.600 58.200 480.000 58.800 ;
        RECT 489.600 58.200 505.800 58.800 ;
        RECT 354.000 57.600 368.400 58.200 ;
        RECT 462.600 57.600 477.600 58.200 ;
        RECT 490.800 57.600 517.800 58.200 ;
        RECT 356.400 57.000 372.000 57.600 ;
        RECT 458.400 57.000 475.200 57.600 ;
        RECT 493.200 57.000 525.000 57.600 ;
        RECT 359.400 56.400 376.200 57.000 ;
        RECT 454.800 56.400 472.200 57.000 ;
        RECT 495.600 56.400 528.600 57.000 ;
        RECT 362.400 55.800 380.400 56.400 ;
        RECT 450.000 55.800 469.200 56.400 ;
        RECT 500.400 55.800 531.000 56.400 ;
        RECT 365.400 55.200 385.200 55.800 ;
        RECT 444.600 55.200 465.600 55.800 ;
        RECT 506.400 55.200 532.800 55.800 ;
        RECT 368.400 54.600 391.200 55.200 ;
        RECT 438.000 54.600 462.000 55.200 ;
        RECT 519.600 54.600 534.000 55.200 ;
        RECT 372.000 54.000 399.600 54.600 ;
        RECT 430.200 54.000 458.400 54.600 ;
        RECT 525.600 54.000 534.600 54.600 ;
        RECT 376.200 53.400 454.200 54.000 ;
        RECT 528.600 53.400 535.200 54.000 ;
        RECT 380.400 52.800 449.400 53.400 ;
        RECT 530.400 52.800 535.200 53.400 ;
        RECT 385.800 52.200 444.600 52.800 ;
        RECT 532.200 52.200 535.800 52.800 ;
        RECT 391.800 51.600 441.600 52.200 ;
        RECT 533.400 51.600 535.800 52.200 ;
        RECT 400.800 51.000 441.600 51.600 ;
        RECT 534.000 51.000 537.000 51.600 ;
        RECT 411.600 49.800 415.200 51.000 ;
        RECT 425.400 50.400 442.200 51.000 ;
        RECT 534.600 50.400 537.600 51.000 ;
        RECT 426.000 49.800 436.200 50.400 ;
        RECT 412.200 48.600 415.800 49.800 ;
        RECT 427.800 49.200 436.200 49.800 ;
        RECT 439.200 49.800 442.800 50.400 ;
        RECT 535.200 49.800 538.200 50.400 ;
        RECT 439.200 49.200 443.400 49.800 ;
        RECT 535.800 49.200 538.800 49.800 ;
        RECT 430.200 48.600 436.800 49.200 ;
        RECT 439.800 48.600 443.400 49.200 ;
        RECT 518.400 48.600 525.000 49.200 ;
        RECT 536.400 48.600 539.400 49.200 ;
        RECT 412.800 48.000 416.400 48.600 ;
        RECT 431.400 48.000 438.600 48.600 ;
        RECT 439.800 48.000 444.000 48.600 ;
        RECT 516.600 48.000 526.200 48.600 ;
        RECT 536.400 48.000 540.000 48.600 ;
        RECT 413.400 46.800 417.000 48.000 ;
        RECT 432.000 47.400 445.200 48.000 ;
        RECT 515.400 47.400 527.400 48.000 ;
        RECT 537.000 47.400 540.000 48.000 ;
        RECT 433.200 46.800 445.800 47.400 ;
        RECT 514.200 46.800 528.600 47.400 ;
        RECT 537.000 46.800 540.600 47.400 ;
        RECT 414.000 46.200 417.600 46.800 ;
        RECT 434.400 46.200 445.800 46.800 ;
        RECT 513.600 46.200 529.200 46.800 ;
        RECT 414.600 45.600 418.200 46.200 ;
        RECT 436.200 45.600 445.200 46.200 ;
        RECT 513.000 45.600 518.400 46.200 ;
        RECT 524.400 45.600 529.800 46.200 ;
        RECT 415.200 45.000 418.800 45.600 ;
        RECT 438.600 45.000 444.600 45.600 ;
        RECT 513.000 45.000 517.200 45.600 ;
        RECT 526.200 45.000 530.400 45.600 ;
        RECT 537.600 45.000 540.600 46.800 ;
        RECT 415.200 44.400 419.400 45.000 ;
        RECT 513.000 44.400 516.000 45.000 ;
        RECT 526.800 44.400 531.000 45.000 ;
        RECT 537.600 44.400 541.200 45.000 ;
        RECT 415.800 43.800 419.400 44.400 ;
        RECT 498.000 43.800 499.200 44.400 ;
        RECT 513.000 43.800 515.400 44.400 ;
        RECT 527.400 43.800 531.600 44.400 ;
        RECT 536.400 43.800 541.800 44.400 ;
        RECT 416.400 43.200 420.000 43.800 ;
        RECT 493.200 43.200 502.800 43.800 ;
        RECT 513.000 43.200 514.800 43.800 ;
        RECT 528.000 43.200 531.600 43.800 ;
        RECT 535.800 43.200 543.000 43.800 ;
        RECT 417.000 42.600 420.600 43.200 ;
        RECT 490.800 42.600 504.600 43.200 ;
        RECT 528.600 42.600 532.200 43.200 ;
        RECT 535.200 42.600 543.600 43.200 ;
        RECT 417.600 42.000 421.200 42.600 ;
        RECT 489.000 42.000 505.800 42.600 ;
        RECT 529.200 42.000 532.200 42.600 ;
        RECT 534.600 42.000 543.600 42.600 ;
        RECT 417.600 41.400 421.800 42.000 ;
        RECT 487.200 41.400 507.000 42.000 ;
        RECT 529.200 41.400 532.800 42.000 ;
        RECT 418.200 40.800 422.400 41.400 ;
        RECT 486.600 40.800 496.800 41.400 ;
        RECT 500.400 40.800 507.600 41.400 ;
        RECT 418.800 40.200 423.000 40.800 ;
        RECT 486.000 40.200 493.200 40.800 ;
        RECT 502.800 40.200 508.800 40.800 ;
        RECT 529.800 40.200 532.800 41.400 ;
        RECT 534.600 41.400 538.200 42.000 ;
        RECT 540.600 41.400 544.200 42.000 ;
        RECT 534.600 40.800 537.600 41.400 ;
        RECT 541.200 40.800 544.200 41.400 ;
        RECT 419.400 39.600 424.200 40.200 ;
        RECT 486.600 39.600 490.800 40.200 ;
        RECT 504.000 39.600 509.400 40.200 ;
        RECT 420.000 39.000 424.800 39.600 ;
        RECT 487.200 39.000 488.400 39.600 ;
        RECT 505.200 39.000 510.000 39.600 ;
        RECT 420.600 38.400 425.400 39.000 ;
        RECT 506.400 38.400 510.600 39.000 ;
        RECT 421.800 37.800 426.000 38.400 ;
        RECT 507.000 37.800 510.600 38.400 ;
        RECT 530.400 37.800 533.400 40.200 ;
        RECT 534.600 37.800 537.000 40.800 ;
        RECT 541.200 40.200 544.800 40.800 ;
        RECT 422.400 37.200 427.200 37.800 ;
        RECT 507.600 37.200 511.200 37.800 ;
        RECT 531.000 37.200 537.000 37.800 ;
        RECT 423.000 36.600 427.800 37.200 ;
        RECT 423.600 36.000 429.000 36.600 ;
        RECT 508.200 36.000 511.800 37.200 ;
        RECT 522.600 36.000 525.600 36.600 ;
        RECT 424.200 35.400 429.600 36.000 ;
        RECT 508.800 35.400 511.800 36.000 ;
        RECT 522.000 35.400 526.200 36.000 ;
        RECT 425.400 34.800 430.800 35.400 ;
        RECT 426.000 34.200 432.000 34.800 ;
        RECT 427.200 33.600 433.800 34.200 ;
        RECT 427.800 33.000 435.600 33.600 ;
        RECT 509.400 33.000 512.400 35.400 ;
        RECT 521.400 34.200 526.800 35.400 ;
        RECT 521.400 33.600 527.400 34.200 ;
        RECT 520.800 33.000 527.400 33.600 ;
        RECT 429.000 32.400 437.400 33.000 ;
        RECT 430.200 31.800 439.800 32.400 ;
        RECT 504.000 31.800 506.400 32.400 ;
        RECT 432.000 31.200 442.200 31.800 ;
        RECT 502.800 31.200 507.600 31.800 ;
        RECT 433.800 30.600 444.600 31.200 ;
        RECT 502.200 30.600 508.200 31.200 ;
        RECT 435.600 30.000 447.600 30.600 ;
        RECT 502.200 30.000 508.800 30.600 ;
        RECT 437.400 29.400 451.200 30.000 ;
        RECT 501.600 29.400 508.800 30.000 ;
        RECT 510.000 29.400 513.000 33.000 ;
        RECT 520.800 32.400 528.000 33.000 ;
        RECT 520.800 30.600 523.800 32.400 ;
        RECT 525.000 30.600 528.000 32.400 ;
        RECT 531.000 31.800 537.600 37.200 ;
        RECT 541.800 34.800 544.800 40.200 ;
        RECT 541.200 33.000 544.200 34.800 ;
        RECT 531.000 31.200 533.400 31.800 ;
        RECT 520.800 30.000 523.200 30.600 ;
        RECT 439.800 28.800 453.600 29.400 ;
        RECT 501.000 28.800 504.600 29.400 ;
        RECT 505.800 28.800 513.000 29.400 ;
        RECT 442.200 28.200 456.000 28.800 ;
        RECT 444.600 27.600 457.800 28.200 ;
        RECT 447.600 27.000 459.600 27.600 ;
        RECT 501.000 27.000 504.000 28.800 ;
        RECT 506.400 27.600 512.400 28.800 ;
        RECT 450.000 26.400 461.400 27.000 ;
        RECT 453.000 25.800 462.600 26.400 ;
        RECT 456.000 25.200 464.400 25.800 ;
        RECT 457.800 24.600 465.600 25.200 ;
        RECT 459.600 24.000 466.800 24.600 ;
        RECT 460.800 23.400 468.600 24.000 ;
        RECT 462.600 22.800 469.800 23.400 ;
        RECT 463.800 22.200 471.000 22.800 ;
        RECT 465.000 21.600 472.200 22.200 ;
        RECT 466.800 21.000 473.400 21.600 ;
        RECT 500.400 21.000 503.400 27.000 ;
        RECT 507.000 25.800 512.400 27.600 ;
        RECT 507.600 23.400 511.800 25.800 ;
        RECT 520.200 23.400 523.200 30.000 ;
        RECT 525.600 30.000 528.000 30.600 ;
        RECT 525.600 25.200 528.600 30.000 ;
        RECT 530.400 27.600 533.400 31.200 ;
        RECT 534.600 28.200 537.600 31.800 ;
        RECT 540.600 32.400 544.200 33.000 ;
        RECT 540.600 31.200 543.600 32.400 ;
        RECT 540.000 30.000 543.000 31.200 ;
        RECT 539.400 29.400 543.000 30.000 ;
        RECT 539.400 28.800 542.400 29.400 ;
        RECT 535.200 27.600 537.600 28.200 ;
        RECT 538.800 28.200 542.400 28.800 ;
        RECT 538.800 27.600 541.800 28.200 ;
        RECT 529.800 25.200 532.800 27.600 ;
        RECT 535.200 27.000 541.800 27.600 ;
        RECT 535.200 25.800 541.200 27.000 ;
        RECT 534.600 25.200 540.600 25.800 ;
        RECT 525.600 24.600 540.600 25.200 ;
        RECT 507.600 21.600 511.200 23.400 ;
        RECT 468.000 20.400 474.600 21.000 ;
        RECT 501.000 20.400 503.400 21.000 ;
        RECT 507.000 20.400 510.600 21.600 ;
        RECT 519.600 20.400 523.200 23.400 ;
        RECT 525.000 23.400 528.000 24.600 ;
        RECT 529.200 23.400 540.000 24.600 ;
        RECT 525.000 22.800 539.400 23.400 ;
        RECT 525.000 22.200 538.800 22.800 ;
        RECT 525.000 21.600 538.200 22.200 ;
        RECT 525.000 21.000 532.800 21.600 ;
        RECT 535.200 21.000 537.600 21.600 ;
        RECT 469.200 19.800 475.800 20.400 ;
        RECT 470.400 19.200 477.000 19.800 ;
        RECT 471.600 18.600 478.200 19.200 ;
        RECT 472.800 18.000 479.400 18.600 ;
        RECT 474.000 17.400 480.600 18.000 ;
        RECT 501.000 17.400 504.000 20.400 ;
        RECT 507.000 19.800 511.200 20.400 ;
        RECT 520.200 19.800 523.200 20.400 ;
        RECT 524.400 20.400 531.000 21.000 ;
        RECT 507.000 19.200 511.800 19.800 ;
        RECT 506.400 18.600 511.800 19.200 ;
        RECT 520.200 18.600 522.600 19.800 ;
        RECT 524.400 19.200 530.400 20.400 ;
        RECT 506.400 18.000 512.400 18.600 ;
        RECT 506.400 17.400 513.000 18.000 ;
        RECT 519.600 17.400 522.600 18.600 ;
        RECT 523.800 18.000 529.800 19.200 ;
        RECT 523.800 17.400 529.200 18.000 ;
        RECT 475.200 16.800 481.800 17.400 ;
        RECT 476.400 16.200 483.600 16.800 ;
        RECT 477.600 15.600 484.800 16.200 ;
        RECT 478.800 15.000 486.000 15.600 ;
        RECT 501.600 15.000 504.600 17.400 ;
        RECT 506.400 16.800 513.600 17.400 ;
        RECT 519.600 16.800 528.600 17.400 ;
        RECT 505.800 15.000 508.800 16.800 ;
        RECT 510.000 16.200 514.800 16.800 ;
        RECT 519.600 16.200 528.000 16.800 ;
        RECT 510.600 15.600 528.000 16.200 ;
        RECT 511.200 15.000 527.400 15.600 ;
        RECT 480.600 14.400 487.200 15.000 ;
        RECT 481.800 13.800 489.000 14.400 ;
        RECT 501.600 13.800 508.200 15.000 ;
        RECT 511.800 14.400 526.200 15.000 ;
        RECT 513.000 13.800 525.600 14.400 ;
        RECT 483.000 13.200 490.800 13.800 ;
        RECT 500.400 13.200 508.200 13.800 ;
        RECT 514.200 13.200 525.000 13.800 ;
        RECT 484.200 12.600 507.600 13.200 ;
        RECT 485.400 12.000 507.600 12.600 ;
        RECT 519.000 12.000 524.400 13.200 ;
        RECT 487.200 11.400 507.600 12.000 ;
        RECT 518.400 11.400 523.800 12.000 ;
        RECT 488.400 10.800 507.000 11.400 ;
        RECT 490.800 10.200 500.400 10.800 ;
        RECT 502.200 10.200 507.000 10.800 ;
        RECT 518.400 10.200 523.200 11.400 ;
        RECT 502.200 8.400 506.400 10.200 ;
        RECT 517.800 9.600 522.600 10.200 ;
        RECT 517.800 9.000 521.400 9.600 ;
        RECT 518.400 8.400 520.800 9.000 ;
        RECT 502.200 7.200 505.800 8.400 ;
        RECT 501.600 6.600 505.200 7.200 ;
        RECT 501.600 6.000 504.600 6.600 ;
        RECT 502.200 5.400 504.600 6.000 ;
        RECT 502.200 4.800 504.000 5.400 ;
      LAYER Metal5 ;
        RECT 103.800 577.200 105.000 577.800 ;
        RECT 103.200 576.600 106.200 577.200 ;
        RECT 103.200 576.000 106.800 576.600 ;
        RECT 103.800 575.400 107.400 576.000 ;
        RECT 103.800 574.800 108.000 575.400 ;
        RECT 104.400 574.200 109.200 574.800 ;
        RECT 104.400 573.600 109.800 574.200 ;
        RECT 104.400 573.000 110.400 573.600 ;
        RECT 104.400 572.400 111.000 573.000 ;
        RECT 104.400 571.800 112.200 572.400 ;
        RECT 105.000 571.200 112.800 571.800 ;
        RECT 105.000 568.800 108.000 571.200 ;
        RECT 109.200 570.600 113.400 571.200 ;
        RECT 109.800 570.000 114.000 570.600 ;
        RECT 110.400 569.400 115.200 570.000 ;
        RECT 111.000 568.800 115.800 569.400 ;
        RECT 105.600 565.800 108.600 568.800 ;
        RECT 112.200 568.200 116.400 568.800 ;
        RECT 112.800 567.600 117.000 568.200 ;
        RECT 113.400 567.000 117.600 567.600 ;
        RECT 114.000 566.400 118.200 567.000 ;
        RECT 114.600 565.800 119.400 566.400 ;
        RECT 106.200 562.800 109.200 565.800 ;
        RECT 115.200 565.200 120.000 565.800 ;
        RECT 116.400 564.600 120.600 565.200 ;
        RECT 117.000 564.000 121.200 564.600 ;
        RECT 117.600 563.400 121.800 564.000 ;
        RECT 118.200 562.800 122.400 563.400 ;
        RECT 106.800 562.200 109.200 562.800 ;
        RECT 118.800 562.200 123.000 562.800 ;
        RECT 106.800 558.000 109.800 562.200 ;
        RECT 119.400 561.600 123.600 562.200 ;
        RECT 120.000 561.000 124.200 561.600 ;
        RECT 120.600 560.400 125.400 561.000 ;
        RECT 121.200 559.800 126.000 560.400 ;
        RECT 122.400 559.200 126.600 559.800 ;
        RECT 123.000 558.600 127.200 559.200 ;
        RECT 123.600 558.000 127.800 558.600 ;
        RECT 107.400 557.400 109.800 558.000 ;
        RECT 124.200 557.400 128.400 558.000 ;
        RECT 107.400 550.200 110.400 557.400 ;
        RECT 124.800 556.800 129.000 557.400 ;
        RECT 125.400 556.200 129.600 556.800 ;
        RECT 126.000 555.600 130.200 556.200 ;
        RECT 126.600 555.000 130.800 555.600 ;
        RECT 127.200 554.400 131.400 555.000 ;
        RECT 127.800 553.800 132.000 554.400 ;
        RECT 128.400 553.200 132.600 553.800 ;
        RECT 129.000 552.600 133.200 553.200 ;
        RECT 129.600 552.000 133.800 552.600 ;
        RECT 130.200 551.400 134.400 552.000 ;
        RECT 130.800 550.800 135.000 551.400 ;
        RECT 131.400 550.200 135.000 550.800 ;
        RECT 108.000 549.000 110.400 550.200 ;
        RECT 132.000 549.600 135.600 550.200 ;
        RECT 132.600 549.000 136.200 549.600 ;
        RECT 7.200 546.000 9.000 546.600 ;
        RECT 6.000 545.400 9.600 546.000 ;
        RECT 6.600 544.800 10.800 545.400 ;
        RECT 6.600 544.200 12.000 544.800 ;
        RECT 7.200 543.600 13.200 544.200 ;
        RECT 7.200 543.000 13.800 543.600 ;
        RECT 7.200 542.400 15.000 543.000 ;
        RECT 7.800 541.800 16.200 542.400 ;
        RECT 7.800 541.200 17.400 541.800 ;
        RECT 8.400 540.600 18.600 541.200 ;
        RECT 8.400 540.000 19.800 540.600 ;
        RECT 9.000 538.800 12.600 540.000 ;
        RECT 14.400 539.400 20.400 540.000 ;
        RECT 15.600 538.800 21.600 539.400 ;
        RECT 9.600 538.200 13.200 538.800 ;
        RECT 16.200 538.200 22.800 538.800 ;
        RECT 10.200 537.000 13.800 538.200 ;
        RECT 17.400 537.600 23.400 538.200 ;
        RECT 18.600 537.000 24.600 537.600 ;
        RECT 10.800 536.400 14.400 537.000 ;
        RECT 19.800 536.400 25.800 537.000 ;
        RECT 10.800 535.800 15.000 536.400 ;
        RECT 21.000 535.800 26.400 536.400 ;
        RECT 11.400 535.200 15.000 535.800 ;
        RECT 21.600 535.200 27.600 535.800 ;
        RECT 12.000 534.000 15.600 535.200 ;
        RECT 22.800 534.600 28.800 535.200 ;
        RECT 24.000 534.000 30.000 534.600 ;
        RECT 108.000 534.000 111.000 549.000 ;
        RECT 133.200 548.400 136.800 549.000 ;
        RECT 133.800 547.800 137.400 548.400 ;
        RECT 133.800 547.200 138.000 547.800 ;
        RECT 134.400 546.600 138.600 547.200 ;
        RECT 135.000 546.000 139.200 546.600 ;
        RECT 135.600 545.400 139.800 546.000 ;
        RECT 136.200 544.800 140.400 545.400 ;
        RECT 136.800 544.200 140.400 544.800 ;
        RECT 137.400 543.600 141.000 544.200 ;
        RECT 138.000 543.000 141.600 543.600 ;
        RECT 138.600 542.400 142.200 543.000 ;
        RECT 138.600 541.800 142.800 542.400 ;
        RECT 139.200 541.200 143.400 541.800 ;
        RECT 139.800 540.600 144.000 541.200 ;
        RECT 140.400 540.000 144.600 540.600 ;
        RECT 141.000 539.400 144.600 540.000 ;
        RECT 141.600 538.800 145.200 539.400 ;
        RECT 142.200 538.200 145.800 538.800 ;
        RECT 142.800 537.600 146.400 538.200 ;
        RECT 142.800 537.000 147.000 537.600 ;
        RECT 143.400 536.400 147.600 537.000 ;
        RECT 144.000 535.800 147.600 536.400 ;
        RECT 144.600 535.200 148.200 535.800 ;
        RECT 145.200 534.600 148.800 535.200 ;
        RECT 12.600 533.400 16.200 534.000 ;
        RECT 24.600 533.400 30.600 534.000 ;
        RECT 13.200 532.200 16.800 533.400 ;
        RECT 25.800 532.800 31.800 533.400 ;
        RECT 27.000 532.200 33.000 532.800 ;
        RECT 108.600 532.200 111.000 534.000 ;
        RECT 145.800 534.000 149.400 534.600 ;
        RECT 145.800 533.400 150.000 534.000 ;
        RECT 146.400 532.800 150.000 533.400 ;
        RECT 147.000 532.200 150.600 532.800 ;
        RECT 271.200 532.200 315.600 537.600 ;
        RECT 13.800 531.600 17.400 532.200 ;
        RECT 27.600 531.600 33.600 532.200 ;
        RECT 14.400 531.000 17.400 531.600 ;
        RECT 28.800 531.000 34.800 531.600 ;
        RECT 14.400 530.400 18.000 531.000 ;
        RECT 29.400 530.400 36.000 531.000 ;
        RECT 15.000 529.200 18.600 530.400 ;
        RECT 30.600 529.800 36.600 530.400 ;
        RECT 31.800 529.200 37.800 529.800 ;
        RECT 15.600 528.600 19.200 529.200 ;
        RECT 33.000 528.600 39.000 529.200 ;
        RECT 16.200 528.000 19.200 528.600 ;
        RECT 34.200 528.000 39.600 528.600 ;
        RECT 16.200 527.400 19.800 528.000 ;
        RECT 35.400 527.400 40.800 528.000 ;
        RECT 16.800 526.200 20.400 527.400 ;
        RECT 36.000 526.800 42.000 527.400 ;
        RECT 37.200 526.200 42.600 526.800 ;
        RECT 17.400 525.600 21.000 526.200 ;
        RECT 38.400 525.600 43.800 526.200 ;
        RECT 18.000 525.000 21.000 525.600 ;
        RECT 39.000 525.000 44.400 525.600 ;
        RECT 18.000 524.400 21.600 525.000 ;
        RECT 40.200 524.400 45.600 525.000 ;
        RECT 18.600 523.800 21.600 524.400 ;
        RECT 40.800 523.800 46.800 524.400 ;
        RECT 18.600 523.200 22.200 523.800 ;
        RECT 42.000 523.200 47.400 523.800 ;
        RECT 19.200 522.600 22.800 523.200 ;
        RECT 43.200 522.600 48.600 523.200 ;
        RECT 108.600 522.600 111.600 532.200 ;
        RECT 147.600 531.600 151.200 532.200 ;
        RECT 148.200 531.000 151.800 531.600 ;
        RECT 148.200 530.400 152.400 531.000 ;
        RECT 148.800 529.800 152.400 530.400 ;
        RECT 149.400 529.200 153.000 529.800 ;
        RECT 150.000 528.600 153.600 529.200 ;
        RECT 150.600 528.000 154.200 528.600 ;
        RECT 150.600 527.400 154.800 528.000 ;
        RECT 151.200 526.800 154.800 527.400 ;
        RECT 151.800 526.200 155.400 526.800 ;
        RECT 152.400 525.600 156.000 526.200 ;
        RECT 153.000 524.400 156.600 525.600 ;
        RECT 153.600 523.800 157.200 524.400 ;
        RECT 154.200 523.200 157.800 523.800 ;
        RECT 19.800 522.000 22.800 522.600 ;
        RECT 43.800 522.000 49.800 522.600 ;
        RECT 109.200 522.000 111.600 522.600 ;
        RECT 154.800 522.000 158.400 523.200 ;
        RECT 19.800 521.400 23.400 522.000 ;
        RECT 45.000 521.400 50.400 522.000 ;
        RECT 20.400 520.800 23.400 521.400 ;
        RECT 46.200 520.800 51.600 521.400 ;
        RECT 20.400 520.200 24.000 520.800 ;
        RECT 46.800 520.200 52.200 520.800 ;
        RECT 21.000 519.600 24.000 520.200 ;
        RECT 48.000 519.600 53.400 520.200 ;
        RECT 21.000 519.000 24.600 519.600 ;
        RECT 48.600 519.000 54.000 519.600 ;
        RECT 21.600 518.400 24.600 519.000 ;
        RECT 49.800 518.400 55.200 519.000 ;
        RECT 21.600 517.800 25.200 518.400 ;
        RECT 51.000 517.800 56.400 518.400 ;
        RECT 22.200 517.200 25.200 517.800 ;
        RECT 51.600 517.200 57.000 517.800 ;
        RECT 22.200 516.600 25.800 517.200 ;
        RECT 52.800 516.600 58.200 517.200 ;
        RECT 22.800 516.000 25.800 516.600 ;
        RECT 53.400 516.000 58.800 516.600 ;
        RECT 109.200 516.000 112.200 522.000 ;
        RECT 155.400 521.400 159.000 522.000 ;
        RECT 156.000 520.800 159.600 521.400 ;
        RECT 156.600 519.600 160.200 520.800 ;
        RECT 157.200 519.000 160.800 519.600 ;
        RECT 157.800 518.400 161.400 519.000 ;
        RECT 158.400 517.200 162.000 518.400 ;
        RECT 159.000 516.600 162.600 517.200 ;
        RECT 159.600 516.000 163.200 516.600 ;
        RECT 22.800 515.400 26.400 516.000 ;
        RECT 54.600 515.400 60.000 516.000 ;
        RECT 109.800 515.400 112.200 516.000 ;
        RECT 23.400 514.200 26.400 515.400 ;
        RECT 55.200 514.800 60.600 515.400 ;
        RECT 56.400 514.200 61.800 514.800 ;
        RECT 24.000 513.000 27.000 514.200 ;
        RECT 57.600 513.600 63.000 514.200 ;
        RECT 58.200 513.000 63.600 513.600 ;
        RECT 24.000 512.400 27.600 513.000 ;
        RECT 59.400 512.400 64.800 513.000 ;
        RECT 24.600 511.800 27.600 512.400 ;
        RECT 60.000 511.800 65.400 512.400 ;
        RECT 24.600 511.200 28.200 511.800 ;
        RECT 61.200 511.200 66.600 511.800 ;
        RECT 25.200 510.600 28.200 511.200 ;
        RECT 61.800 510.600 67.200 511.200 ;
        RECT 109.800 510.600 112.800 515.400 ;
        RECT 160.200 514.800 163.800 516.000 ;
        RECT 160.800 514.200 164.400 514.800 ;
        RECT 161.400 513.600 165.000 514.200 ;
        RECT 162.000 512.400 165.600 513.600 ;
        RECT 162.600 511.800 166.200 512.400 ;
        RECT 163.200 510.600 166.800 511.800 ;
        RECT 25.200 510.000 28.800 510.600 ;
        RECT 63.000 510.000 68.400 510.600 ;
        RECT 25.800 508.800 28.800 510.000 ;
        RECT 63.600 509.400 69.000 510.000 ;
        RECT 64.800 508.800 70.200 509.400 ;
        RECT 26.400 507.600 29.400 508.800 ;
        RECT 65.400 508.200 70.800 508.800 ;
        RECT 66.600 507.600 72.000 508.200 ;
        RECT 26.400 507.000 30.000 507.600 ;
        RECT 67.200 507.000 72.600 507.600 ;
        RECT 110.400 507.000 113.400 510.600 ;
        RECT 163.800 510.000 167.400 510.600 ;
        RECT 164.400 509.400 168.000 510.000 ;
        RECT 164.400 508.800 168.600 509.400 ;
        RECT 165.000 508.200 168.600 508.800 ;
        RECT 165.600 507.600 169.200 508.200 ;
        RECT 165.600 507.000 169.800 507.600 ;
        RECT 27.000 506.400 30.000 507.000 ;
        RECT 68.400 506.400 73.800 507.000 ;
        RECT 27.000 505.800 30.600 506.400 ;
        RECT 69.000 505.800 74.400 506.400 ;
        RECT 27.600 505.200 30.600 505.800 ;
        RECT 70.200 505.200 75.600 505.800 ;
        RECT 27.600 504.600 31.200 505.200 ;
        RECT 70.800 504.600 76.200 505.200 ;
        RECT 111.000 504.600 114.000 507.000 ;
        RECT 166.200 506.400 170.400 507.000 ;
        RECT 166.800 505.800 170.400 506.400 ;
        RECT 167.400 505.200 171.000 505.800 ;
        RECT 168.000 504.600 171.600 505.200 ;
        RECT 28.200 503.400 31.200 504.600 ;
        RECT 72.000 504.000 77.400 504.600 ;
        RECT 72.600 503.400 78.000 504.000 ;
        RECT 28.800 502.200 31.800 503.400 ;
        RECT 73.800 502.800 79.200 503.400 ;
        RECT 75.000 502.200 79.800 502.800 ;
        RECT 28.800 501.600 32.400 502.200 ;
        RECT 75.600 501.600 81.000 502.200 ;
        RECT 111.600 501.600 114.600 504.600 ;
        RECT 168.000 504.000 172.200 504.600 ;
        RECT 168.600 503.400 172.200 504.000 ;
        RECT 169.200 502.800 172.800 503.400 ;
        RECT 169.800 502.200 173.400 502.800 ;
        RECT 169.800 501.600 174.000 502.200 ;
        RECT 29.400 501.000 32.400 501.600 ;
        RECT 76.800 501.000 81.600 501.600 ;
        RECT 29.400 500.400 33.000 501.000 ;
        RECT 77.400 500.400 82.800 501.000 ;
        RECT 30.000 499.800 33.000 500.400 ;
        RECT 78.600 499.800 83.400 500.400 ;
        RECT 30.000 499.200 33.600 499.800 ;
        RECT 79.200 499.200 84.600 499.800 ;
        RECT 112.200 499.200 115.200 501.600 ;
        RECT 170.400 501.000 174.000 501.600 ;
        RECT 171.000 500.400 174.600 501.000 ;
        RECT 178.800 500.400 180.600 501.000 ;
        RECT 171.600 499.200 175.200 500.400 ;
        RECT 177.000 499.800 181.800 500.400 ;
        RECT 176.400 499.200 183.000 499.800 ;
        RECT 30.600 498.000 33.600 499.200 ;
        RECT 80.400 498.600 85.200 499.200 ;
        RECT 81.000 498.000 86.400 498.600 ;
        RECT 31.200 496.800 34.200 498.000 ;
        RECT 82.200 497.400 87.000 498.000 ;
        RECT 112.800 497.400 115.800 499.200 ;
        RECT 172.200 498.600 184.200 499.200 ;
        RECT 172.800 498.000 184.800 498.600 ;
        RECT 82.800 496.800 88.200 497.400 ;
        RECT 113.400 496.800 115.800 497.400 ;
        RECT 173.400 497.400 178.800 498.000 ;
        RECT 180.000 497.400 185.400 498.000 ;
        RECT 173.400 496.800 178.200 497.400 ;
        RECT 181.200 496.800 186.000 497.400 ;
        RECT 31.200 496.200 34.800 496.800 ;
        RECT 84.000 496.200 88.800 496.800 ;
        RECT 31.800 495.600 34.800 496.200 ;
        RECT 84.600 495.600 90.000 496.200 ;
        RECT 113.400 495.600 116.400 496.800 ;
        RECT 174.000 496.200 178.200 496.800 ;
        RECT 182.400 496.200 186.600 496.800 ;
        RECT 174.600 495.600 178.200 496.200 ;
        RECT 183.000 495.600 187.200 496.200 ;
        RECT 31.800 495.000 35.400 495.600 ;
        RECT 85.800 495.000 90.600 495.600 ;
        RECT 114.000 495.000 116.400 495.600 ;
        RECT 32.400 494.400 35.400 495.000 ;
        RECT 86.400 494.400 91.800 495.000 ;
        RECT 32.400 493.800 36.000 494.400 ;
        RECT 87.600 493.800 92.400 494.400 ;
        RECT 114.000 493.800 117.000 495.000 ;
        RECT 33.000 492.600 36.000 493.800 ;
        RECT 88.200 493.200 93.600 493.800 ;
        RECT 114.600 493.200 117.000 493.800 ;
        RECT 89.400 492.600 94.200 493.200 ;
        RECT 33.600 491.400 36.600 492.600 ;
        RECT 90.000 492.000 95.400 492.600 ;
        RECT 114.600 492.000 117.600 493.200 ;
        RECT 91.200 491.400 96.000 492.000 ;
        RECT 33.600 490.800 37.200 491.400 ;
        RECT 91.800 490.800 97.200 491.400 ;
        RECT 115.200 490.800 117.600 492.000 ;
        RECT 155.400 491.400 157.800 492.000 ;
        RECT 154.200 490.800 158.400 491.400 ;
        RECT 175.200 490.800 178.200 495.600 ;
        RECT 183.600 495.000 187.200 495.600 ;
        RECT 184.200 494.400 187.800 495.000 ;
        RECT 184.800 493.800 187.800 494.400 ;
        RECT 184.800 493.200 188.400 493.800 ;
        RECT 185.400 492.600 188.400 493.200 ;
        RECT 185.400 492.000 189.000 492.600 ;
        RECT 186.000 490.800 189.000 492.000 ;
        RECT 34.200 490.200 37.200 490.800 ;
        RECT 93.000 490.200 97.800 490.800 ;
        RECT 113.400 490.200 118.200 490.800 ;
        RECT 153.600 490.200 159.000 490.800 ;
        RECT 34.200 489.600 37.800 490.200 ;
        RECT 93.600 489.600 99.000 490.200 ;
        RECT 111.000 489.600 121.800 490.200 ;
        RECT 132.000 489.600 138.600 490.200 ;
        RECT 153.600 489.600 159.600 490.200 ;
        RECT 34.800 489.000 37.800 489.600 ;
        RECT 94.800 489.000 100.200 489.600 ;
        RECT 109.800 489.000 123.600 489.600 ;
        RECT 131.400 489.000 140.400 489.600 ;
        RECT 34.800 488.400 38.400 489.000 ;
        RECT 95.400 488.400 100.800 489.000 ;
        RECT 109.200 488.400 125.400 489.000 ;
        RECT 130.800 488.400 142.800 489.000 ;
        RECT 153.000 488.400 160.200 489.600 ;
        RECT 175.800 489.000 178.800 490.800 ;
        RECT 175.800 488.400 179.400 489.000 ;
        RECT 35.400 487.800 38.400 488.400 ;
        RECT 96.600 487.800 102.000 488.400 ;
        RECT 108.600 487.800 127.200 488.400 ;
        RECT 130.800 487.800 144.600 488.400 ;
        RECT 152.400 487.800 156.000 488.400 ;
        RECT 157.200 487.800 160.800 488.400 ;
        RECT 35.400 487.200 39.000 487.800 ;
        RECT 97.200 487.200 102.600 487.800 ;
        RECT 108.600 487.200 113.400 487.800 ;
        RECT 120.000 487.200 128.400 487.800 ;
        RECT 130.800 487.200 145.800 487.800 ;
        RECT 36.000 486.000 39.000 487.200 ;
        RECT 98.400 486.600 103.800 487.200 ;
        RECT 99.000 486.000 104.400 486.600 ;
        RECT 108.600 486.000 111.600 487.200 ;
        RECT 121.800 486.600 129.600 487.200 ;
        RECT 130.800 486.600 134.400 487.200 ;
        RECT 138.600 486.600 147.600 487.200 ;
        RECT 152.400 486.600 155.400 487.800 ;
        RECT 157.800 487.200 160.800 487.800 ;
        RECT 176.400 487.200 179.400 488.400 ;
        RECT 157.800 486.600 161.400 487.200 ;
        RECT 123.600 486.000 134.400 486.600 ;
        RECT 140.400 486.000 148.800 486.600 ;
        RECT 151.800 486.000 155.400 486.600 ;
        RECT 36.600 484.800 39.600 486.000 ;
        RECT 100.200 485.400 105.600 486.000 ;
        RECT 108.600 485.400 112.200 486.000 ;
        RECT 125.400 485.400 135.000 486.000 ;
        RECT 142.200 485.400 150.600 486.000 ;
        RECT 151.800 485.400 154.800 486.000 ;
        RECT 158.400 485.400 161.400 486.600 ;
        RECT 177.000 486.000 180.000 487.200 ;
        RECT 186.600 486.000 189.600 490.800 ;
        RECT 194.400 489.000 198.600 489.600 ;
        RECT 193.200 488.400 199.800 489.000 ;
        RECT 192.600 487.800 200.400 488.400 ;
        RECT 192.000 487.200 201.000 487.800 ;
        RECT 191.400 486.600 201.000 487.200 ;
        RECT 190.800 486.000 195.000 486.600 ;
        RECT 198.000 486.000 201.600 486.600 ;
        RECT 289.800 486.000 297.000 532.200 ;
        RECT 321.000 520.800 328.200 540.000 ;
        RECT 336.600 525.600 344.400 526.200 ;
        RECT 377.400 525.600 386.400 526.200 ;
        RECT 334.800 525.000 346.200 525.600 ;
        RECT 375.000 525.000 388.200 525.600 ;
        RECT 333.600 524.400 347.400 525.000 ;
        RECT 373.800 524.400 389.400 525.000 ;
        RECT 332.400 523.800 348.600 524.400 ;
        RECT 372.600 523.800 390.600 524.400 ;
        RECT 331.800 523.200 349.200 523.800 ;
        RECT 371.400 523.200 391.800 523.800 ;
        RECT 331.200 522.600 349.800 523.200 ;
        RECT 370.800 522.600 392.400 523.200 ;
        RECT 330.000 522.000 350.400 522.600 ;
        RECT 370.200 522.000 393.600 522.600 ;
        RECT 329.400 520.800 351.000 522.000 ;
        RECT 369.600 521.400 394.200 522.000 ;
        RECT 369.000 520.800 394.800 521.400 ;
        RECT 321.000 520.200 337.200 520.800 ;
        RECT 340.800 520.200 351.600 520.800 ;
        RECT 368.400 520.200 379.800 520.800 ;
        RECT 383.400 520.200 394.800 520.800 ;
        RECT 321.000 519.600 334.800 520.200 ;
        RECT 342.600 519.600 352.200 520.200 ;
        RECT 367.800 519.600 378.000 520.200 ;
        RECT 385.800 519.600 395.400 520.200 ;
        RECT 321.000 519.000 333.600 519.600 ;
        RECT 343.800 519.000 352.200 519.600 ;
        RECT 367.200 519.000 376.800 519.600 ;
        RECT 387.000 519.000 396.000 519.600 ;
        RECT 321.000 518.400 332.400 519.000 ;
        RECT 344.400 518.400 352.800 519.000 ;
        RECT 367.200 518.400 375.600 519.000 ;
        RECT 387.600 518.400 396.600 519.000 ;
        RECT 321.000 517.800 331.800 518.400 ;
        RECT 345.000 517.800 352.800 518.400 ;
        RECT 366.600 517.800 375.000 518.400 ;
        RECT 388.200 517.800 396.600 518.400 ;
        RECT 321.000 517.200 331.200 517.800 ;
        RECT 345.600 517.200 352.800 517.800 ;
        RECT 366.000 517.200 374.400 517.800 ;
        RECT 388.800 517.200 397.200 517.800 ;
        RECT 321.000 516.600 330.600 517.200 ;
        RECT 345.600 516.600 353.400 517.200 ;
        RECT 321.000 515.400 330.000 516.600 ;
        RECT 346.200 515.400 353.400 516.600 ;
        RECT 366.000 516.000 373.800 517.200 ;
        RECT 389.400 516.600 397.200 517.200 ;
        RECT 321.000 514.200 329.400 515.400 ;
        RECT 346.800 514.200 353.400 515.400 ;
        RECT 365.400 515.400 373.200 516.000 ;
        RECT 390.000 515.400 397.800 516.600 ;
        RECT 365.400 514.800 372.600 515.400 ;
        RECT 364.800 514.200 372.600 514.800 ;
        RECT 390.600 514.800 397.800 515.400 ;
        RECT 390.600 514.200 398.400 514.800 ;
        RECT 321.000 512.400 328.800 514.200 ;
        RECT 346.800 512.400 354.000 514.200 ;
        RECT 364.800 512.400 372.000 514.200 ;
        RECT 391.200 513.000 398.400 514.200 ;
        RECT 321.000 486.000 328.200 512.400 ;
        RECT 347.400 486.000 354.000 512.400 ;
        RECT 364.200 510.000 371.400 512.400 ;
        RECT 391.800 510.600 399.000 513.000 ;
        RECT 392.400 510.000 399.000 510.600 ;
        RECT 364.200 508.800 370.800 510.000 ;
        RECT 363.600 502.200 370.800 508.800 ;
        RECT 364.200 501.000 370.800 502.200 ;
        RECT 392.400 501.000 399.600 510.000 ;
        RECT 364.200 498.600 371.400 501.000 ;
        RECT 392.400 500.400 399.000 501.000 ;
        RECT 364.800 496.800 372.000 498.600 ;
        RECT 391.800 498.000 399.000 500.400 ;
        RECT 391.200 496.800 398.400 498.000 ;
        RECT 364.800 496.200 372.600 496.800 ;
        RECT 365.400 495.600 372.600 496.200 ;
        RECT 390.600 496.200 398.400 496.800 ;
        RECT 390.600 495.600 397.800 496.200 ;
        RECT 365.400 495.000 373.200 495.600 ;
        RECT 366.000 494.400 373.200 495.000 ;
        RECT 390.000 494.400 397.800 495.600 ;
        RECT 366.000 493.800 373.800 494.400 ;
        RECT 389.400 493.800 397.200 494.400 ;
        RECT 366.000 493.200 374.400 493.800 ;
        RECT 388.800 493.200 397.200 493.800 ;
        RECT 366.600 492.600 375.000 493.200 ;
        RECT 388.200 492.600 396.600 493.200 ;
        RECT 367.200 492.000 375.600 492.600 ;
        RECT 387.600 492.000 396.600 492.600 ;
        RECT 367.200 491.400 376.800 492.000 ;
        RECT 387.000 491.400 396.000 492.000 ;
        RECT 367.800 490.800 378.000 491.400 ;
        RECT 385.800 490.800 395.400 491.400 ;
        RECT 368.400 490.200 379.800 490.800 ;
        RECT 383.400 490.200 394.800 490.800 ;
        RECT 369.000 489.600 394.800 490.200 ;
        RECT 369.600 489.000 394.200 489.600 ;
        RECT 370.200 488.400 393.600 489.000 ;
        RECT 370.800 487.800 392.400 488.400 ;
        RECT 371.400 487.200 391.800 487.800 ;
        RECT 372.600 486.600 390.600 487.200 ;
        RECT 373.800 486.000 389.400 486.600 ;
        RECT 409.800 486.000 416.400 540.000 ;
        RECT 429.600 532.200 436.200 540.000 ;
        RECT 464.400 525.600 472.200 526.200 ;
        RECT 462.600 525.000 474.000 525.600 ;
        RECT 429.600 486.000 436.200 525.000 ;
        RECT 448.800 520.800 456.000 525.000 ;
        RECT 461.400 524.400 475.200 525.000 ;
        RECT 460.200 523.800 476.400 524.400 ;
        RECT 459.600 523.200 477.000 523.800 ;
        RECT 459.000 522.600 477.600 523.200 ;
        RECT 457.800 522.000 478.200 522.600 ;
        RECT 457.200 520.800 478.800 522.000 ;
        RECT 448.800 520.200 465.000 520.800 ;
        RECT 468.600 520.200 479.400 520.800 ;
        RECT 448.800 519.600 462.600 520.200 ;
        RECT 470.400 519.600 480.000 520.200 ;
        RECT 448.800 519.000 461.400 519.600 ;
        RECT 471.600 519.000 480.000 519.600 ;
        RECT 448.800 518.400 460.200 519.000 ;
        RECT 472.200 518.400 480.600 519.000 ;
        RECT 448.800 517.800 459.600 518.400 ;
        RECT 472.800 517.800 480.600 518.400 ;
        RECT 448.800 517.200 459.000 517.800 ;
        RECT 473.400 517.200 480.600 517.800 ;
        RECT 448.800 516.600 458.400 517.200 ;
        RECT 473.400 516.600 481.200 517.200 ;
        RECT 448.800 515.400 457.800 516.600 ;
        RECT 474.000 515.400 481.200 516.600 ;
        RECT 448.800 514.200 457.200 515.400 ;
        RECT 474.600 514.200 481.200 515.400 ;
        RECT 448.800 512.400 456.600 514.200 ;
        RECT 474.600 512.400 481.800 514.200 ;
        RECT 448.800 486.000 456.000 512.400 ;
        RECT 475.200 486.000 481.800 512.400 ;
        RECT 177.000 485.400 180.600 486.000 ;
        RECT 100.800 484.800 106.800 485.400 ;
        RECT 109.200 484.800 113.400 485.400 ;
        RECT 126.600 484.800 135.600 485.400 ;
        RECT 144.000 484.800 154.800 485.400 ;
        RECT 37.200 483.600 40.200 484.800 ;
        RECT 102.000 484.200 107.400 484.800 ;
        RECT 109.200 484.200 114.600 484.800 ;
        RECT 127.800 484.200 136.200 484.800 ;
        RECT 145.800 484.200 154.800 484.800 ;
        RECT 103.200 483.600 115.200 484.200 ;
        RECT 129.000 483.600 136.800 484.200 ;
        RECT 147.000 483.600 154.800 484.200 ;
        RECT 159.000 484.200 162.000 485.400 ;
        RECT 169.800 484.800 173.400 485.400 ;
        RECT 177.600 484.800 180.600 485.400 ;
        RECT 186.600 485.400 194.400 486.000 ;
        RECT 186.600 484.800 193.800 485.400 ;
        RECT 198.600 484.800 201.600 486.000 ;
        RECT 375.000 485.400 388.200 486.000 ;
        RECT 377.400 484.800 386.400 485.400 ;
        RECT 168.600 484.200 175.200 484.800 ;
        RECT 177.600 484.200 181.200 484.800 ;
        RECT 186.600 484.200 193.200 484.800 ;
        RECT 198.600 484.200 208.200 484.800 ;
        RECT 159.000 483.600 162.600 484.200 ;
        RECT 168.000 483.600 176.400 484.200 ;
        RECT 37.200 483.000 40.800 483.600 ;
        RECT 103.800 483.000 117.000 483.600 ;
        RECT 130.200 483.000 137.400 483.600 ;
        RECT 148.800 483.000 154.800 483.600 ;
        RECT 37.800 482.400 40.800 483.000 ;
        RECT 105.000 482.400 118.200 483.000 ;
        RECT 131.400 482.400 138.000 483.000 ;
        RECT 150.000 482.400 154.800 483.000 ;
        RECT 159.600 482.400 162.600 483.600 ;
        RECT 167.400 483.000 177.000 483.600 ;
        RECT 178.200 483.000 181.800 484.200 ;
        RECT 186.600 483.600 192.600 484.200 ;
        RECT 198.000 483.600 209.400 484.200 ;
        RECT 166.800 482.400 182.400 483.000 ;
        RECT 37.800 481.800 41.400 482.400 ;
        RECT 105.600 481.800 120.000 482.400 ;
        RECT 134.400 481.800 139.200 482.400 ;
        RECT 38.400 481.200 41.400 481.800 ;
        RECT 106.800 481.200 122.400 481.800 ;
        RECT 135.000 481.200 139.800 481.800 ;
        RECT 38.400 480.600 42.000 481.200 ;
        RECT 106.800 480.600 124.800 481.200 ;
        RECT 135.600 480.600 141.000 481.200 ;
        RECT 39.000 480.000 42.000 480.600 ;
        RECT 105.000 480.000 127.800 480.600 ;
        RECT 136.800 480.000 141.600 480.600 ;
        RECT 151.800 480.000 154.200 482.400 ;
        RECT 159.600 481.800 163.200 482.400 ;
        RECT 160.200 480.600 163.200 481.800 ;
        RECT 166.800 481.800 170.400 482.400 ;
        RECT 173.400 481.800 182.400 482.400 ;
        RECT 186.600 482.400 192.000 483.600 ;
        RECT 196.200 483.000 210.000 483.600 ;
        RECT 195.000 482.400 210.000 483.000 ;
        RECT 166.800 480.600 169.800 481.800 ;
        RECT 174.600 481.200 183.000 481.800 ;
        RECT 186.600 481.200 191.400 482.400 ;
        RECT 193.800 481.800 210.000 482.400 ;
        RECT 192.600 481.200 201.000 481.800 ;
        RECT 175.800 480.600 183.600 481.200 ;
        RECT 186.600 480.600 201.000 481.200 ;
        RECT 205.200 480.600 210.000 481.800 ;
        RECT 39.000 479.400 42.600 480.000 ;
        RECT 103.800 479.400 114.600 480.000 ;
        RECT 117.600 479.400 130.200 480.000 ;
        RECT 137.400 479.400 142.800 480.000 ;
        RECT 39.600 478.800 42.600 479.400 ;
        RECT 102.600 478.800 111.000 479.400 ;
        RECT 120.000 478.800 132.600 479.400 ;
        RECT 138.000 478.800 144.000 479.400 ;
        RECT 39.600 478.200 43.200 478.800 ;
        RECT 102.000 478.200 108.600 478.800 ;
        RECT 122.400 478.200 133.800 478.800 ;
        RECT 139.200 478.200 145.200 478.800 ;
        RECT 40.200 477.600 43.200 478.200 ;
        RECT 100.800 477.600 106.800 478.200 ;
        RECT 124.800 477.600 133.200 478.200 ;
        RECT 140.400 477.600 146.400 478.200 ;
        RECT 40.200 477.000 43.800 477.600 ;
        RECT 100.200 477.000 105.600 477.600 ;
        RECT 141.000 477.000 147.600 477.600 ;
        RECT 40.800 476.400 43.800 477.000 ;
        RECT 99.000 476.400 104.400 477.000 ;
        RECT 142.200 476.400 148.800 477.000 ;
        RECT 40.800 475.800 44.400 476.400 ;
        RECT 98.400 475.800 103.200 476.400 ;
        RECT 144.000 475.800 150.000 476.400 ;
        RECT 151.800 475.800 154.800 480.000 ;
        RECT 160.800 479.400 163.800 480.600 ;
        RECT 160.800 478.800 164.400 479.400 ;
        RECT 161.400 478.200 164.400 478.800 ;
        RECT 166.200 478.200 169.200 480.600 ;
        RECT 176.400 480.000 184.200 480.600 ;
        RECT 177.600 479.400 184.200 480.000 ;
        RECT 186.600 479.400 200.400 480.600 ;
        RECT 205.200 480.000 209.400 480.600 ;
        RECT 205.800 479.400 208.800 480.000 ;
        RECT 178.200 478.800 184.800 479.400 ;
        RECT 186.600 478.800 194.400 479.400 ;
        RECT 178.800 478.200 185.400 478.800 ;
        RECT 161.400 477.600 165.000 478.200 ;
        RECT 162.000 476.400 165.000 477.600 ;
        RECT 166.800 476.400 169.800 478.200 ;
        RECT 180.000 477.600 185.400 478.200 ;
        RECT 186.600 478.200 193.200 478.800 ;
        RECT 196.200 478.200 199.800 479.400 ;
        RECT 186.600 477.600 192.600 478.200 ;
        RECT 195.600 477.600 199.200 478.200 ;
        RECT 180.600 477.000 192.000 477.600 ;
        RECT 195.000 477.000 198.600 477.600 ;
        RECT 181.200 476.400 191.400 477.000 ;
        RECT 193.800 476.400 198.000 477.000 ;
        RECT 162.000 475.800 165.600 476.400 ;
        RECT 166.800 475.800 170.400 476.400 ;
        RECT 182.400 475.800 190.800 476.400 ;
        RECT 193.200 475.800 197.400 476.400 ;
        RECT 41.400 475.200 44.400 475.800 ;
        RECT 97.800 475.200 102.600 475.800 ;
        RECT 145.200 475.200 155.400 475.800 ;
        RECT 41.400 474.600 45.000 475.200 ;
        RECT 97.200 474.600 102.000 475.200 ;
        RECT 147.600 474.600 155.400 475.200 ;
        RECT 162.600 475.200 165.600 475.800 ;
        RECT 167.400 475.200 170.400 475.800 ;
        RECT 183.000 475.200 190.800 475.800 ;
        RECT 192.000 475.200 197.400 475.800 ;
        RECT 199.200 475.200 205.800 475.800 ;
        RECT 162.600 474.600 166.200 475.200 ;
        RECT 167.400 474.600 171.000 475.200 ;
        RECT 183.600 474.600 207.000 475.200 ;
        RECT 42.000 474.000 45.000 474.600 ;
        RECT 96.600 474.000 100.800 474.600 ;
        RECT 127.800 474.000 130.200 474.600 ;
        RECT 42.000 473.400 45.600 474.000 ;
        RECT 96.000 473.400 100.200 474.000 ;
        RECT 126.600 473.400 130.200 474.000 ;
        RECT 152.400 474.000 155.400 474.600 ;
        RECT 163.200 474.000 166.200 474.600 ;
        RECT 168.000 474.000 171.600 474.600 ;
        RECT 183.600 474.000 208.200 474.600 ;
        RECT 152.400 473.400 156.000 474.000 ;
        RECT 163.200 473.400 166.800 474.000 ;
        RECT 168.000 473.400 172.800 474.000 ;
        RECT 181.200 473.400 208.800 474.000 ;
        RECT 42.600 472.800 45.600 473.400 ;
        RECT 95.400 472.800 99.600 473.400 ;
        RECT 126.000 472.800 129.600 473.400 ;
        RECT 42.600 472.200 46.200 472.800 ;
        RECT 94.800 472.200 99.000 472.800 ;
        RECT 125.400 472.200 129.000 472.800 ;
        RECT 153.000 472.200 156.000 473.400 ;
        RECT 163.800 472.800 166.800 473.400 ;
        RECT 168.600 472.800 208.800 473.400 ;
        RECT 163.800 472.200 167.400 472.800 ;
        RECT 169.200 472.200 199.200 472.800 ;
        RECT 205.800 472.200 208.800 472.800 ;
        RECT 43.200 471.600 46.800 472.200 ;
        RECT 94.200 471.600 98.400 472.200 ;
        RECT 124.800 471.600 128.400 472.200 ;
        RECT 43.800 471.000 46.800 471.600 ;
        RECT 93.600 471.000 97.800 471.600 ;
        RECT 124.200 471.000 127.800 471.600 ;
        RECT 153.600 471.000 156.600 472.200 ;
        RECT 164.400 471.600 167.400 472.200 ;
        RECT 169.800 471.600 195.000 472.200 ;
        RECT 205.800 471.600 209.400 472.200 ;
        RECT 164.400 471.000 168.000 471.600 ;
        RECT 171.000 471.000 185.400 471.600 ;
        RECT 43.800 470.400 47.400 471.000 ;
        RECT 93.600 470.400 97.200 471.000 ;
        RECT 123.600 470.400 127.200 471.000 ;
        RECT 44.400 469.800 47.400 470.400 ;
        RECT 93.000 469.800 96.600 470.400 ;
        RECT 123.000 469.800 127.200 470.400 ;
        RECT 154.200 469.800 157.200 471.000 ;
        RECT 165.000 470.400 168.000 471.000 ;
        RECT 172.800 470.400 184.800 471.000 ;
        RECT 165.000 469.800 168.600 470.400 ;
        RECT 44.400 469.200 48.000 469.800 ;
        RECT 45.000 468.600 48.000 469.200 ;
        RECT 92.400 469.200 96.000 469.800 ;
        RECT 121.800 469.200 126.600 469.800 ;
        RECT 154.800 469.200 157.800 469.800 ;
        RECT 165.600 469.200 168.600 469.800 ;
        RECT 180.600 469.800 184.800 470.400 ;
        RECT 187.800 470.400 192.600 471.600 ;
        RECT 187.800 469.800 193.200 470.400 ;
        RECT 205.800 469.800 208.800 471.600 ;
        RECT 180.600 469.200 184.200 469.800 ;
        RECT 187.800 469.200 193.800 469.800 ;
        RECT 205.200 469.200 208.800 469.800 ;
        RECT 92.400 468.600 95.400 469.200 ;
        RECT 120.600 468.600 126.000 469.200 ;
        RECT 155.400 468.600 158.400 469.200 ;
        RECT 165.600 468.600 169.200 469.200 ;
        RECT 45.000 468.000 48.600 468.600 ;
        RECT 91.800 468.000 95.400 468.600 ;
        RECT 120.000 468.000 126.000 468.600 ;
        RECT 156.000 468.000 158.400 468.600 ;
        RECT 45.600 467.400 48.600 468.000 ;
        RECT 91.200 467.400 94.800 468.000 ;
        RECT 118.800 467.400 125.400 468.000 ;
        RECT 156.000 467.400 159.000 468.000 ;
        RECT 166.200 467.400 169.800 468.600 ;
        RECT 180.000 468.000 183.600 469.200 ;
        RECT 188.400 468.600 194.400 469.200 ;
        RECT 204.600 468.600 208.200 469.200 ;
        RECT 188.400 468.000 195.600 468.600 ;
        RECT 204.000 468.000 208.200 468.600 ;
        RECT 179.400 467.400 183.000 468.000 ;
        RECT 188.400 467.400 196.800 468.000 ;
        RECT 202.800 467.400 207.600 468.000 ;
        RECT 214.200 467.400 217.200 468.000 ;
        RECT 45.600 466.800 49.200 467.400 ;
        RECT 91.200 466.800 94.200 467.400 ;
        RECT 118.200 466.800 125.400 467.400 ;
        RECT 156.600 466.800 159.600 467.400 ;
        RECT 166.800 466.800 170.400 467.400 ;
        RECT 179.400 466.800 182.400 467.400 ;
        RECT 46.200 465.600 49.800 466.800 ;
        RECT 90.600 466.200 94.200 466.800 ;
        RECT 117.600 466.200 124.800 466.800 ;
        RECT 156.600 466.200 160.200 466.800 ;
        RECT 167.400 466.200 170.400 466.800 ;
        RECT 178.800 466.200 182.400 466.800 ;
        RECT 187.800 466.800 198.600 467.400 ;
        RECT 200.400 466.800 207.000 467.400 ;
        RECT 212.400 466.800 219.000 467.400 ;
        RECT 187.800 466.200 206.400 466.800 ;
        RECT 211.200 466.200 219.600 466.800 ;
        RECT 90.600 465.600 93.600 466.200 ;
        RECT 117.000 465.600 124.800 466.200 ;
        RECT 157.200 465.600 160.800 466.200 ;
        RECT 167.400 465.600 171.000 466.200 ;
        RECT 178.800 465.600 181.800 466.200 ;
        RECT 46.800 465.000 50.400 465.600 ;
        RECT 47.400 464.400 50.400 465.000 ;
        RECT 90.000 465.000 93.600 465.600 ;
        RECT 116.400 465.000 124.200 465.600 ;
        RECT 90.000 464.400 93.000 465.000 ;
        RECT 115.800 464.400 124.200 465.000 ;
        RECT 157.800 465.000 161.400 465.600 ;
        RECT 168.000 465.000 171.600 465.600 ;
        RECT 178.200 465.000 181.800 465.600 ;
        RECT 187.800 465.000 190.800 466.200 ;
        RECT 192.600 465.600 205.200 466.200 ;
        RECT 210.600 465.600 220.800 466.200 ;
        RECT 193.800 465.000 204.600 465.600 ;
        RECT 210.000 465.000 221.400 465.600 ;
        RECT 157.800 464.400 162.000 465.000 ;
        RECT 168.600 464.400 172.200 465.000 ;
        RECT 178.200 464.400 181.200 465.000 ;
        RECT 47.400 463.800 51.000 464.400 ;
        RECT 48.000 463.200 51.000 463.800 ;
        RECT 89.400 463.800 93.000 464.400 ;
        RECT 115.200 463.800 119.400 464.400 ;
        RECT 89.400 463.200 92.400 463.800 ;
        RECT 114.600 463.200 118.800 463.800 ;
        RECT 48.000 462.600 51.600 463.200 ;
        RECT 88.800 462.600 92.400 463.200 ;
        RECT 114.000 462.600 118.200 463.200 ;
        RECT 120.600 462.600 123.600 464.400 ;
        RECT 158.400 463.800 162.600 464.400 ;
        RECT 168.600 463.800 172.800 464.400 ;
        RECT 159.000 463.200 163.200 463.800 ;
        RECT 169.200 463.200 172.800 463.800 ;
        RECT 177.600 463.800 181.200 464.400 ;
        RECT 187.200 463.800 190.800 465.000 ;
        RECT 195.600 464.400 202.800 465.000 ;
        RECT 209.400 464.400 214.200 465.000 ;
        RECT 216.600 464.400 222.000 465.000 ;
        RECT 192.600 463.800 193.200 464.400 ;
        RECT 197.400 463.800 201.600 464.400 ;
        RECT 208.800 463.800 213.000 464.400 ;
        RECT 218.400 463.800 222.600 464.400 ;
        RECT 159.000 462.600 163.800 463.200 ;
        RECT 169.800 462.600 173.400 463.200 ;
        RECT 177.600 462.600 180.600 463.800 ;
        RECT 186.600 463.200 195.000 463.800 ;
        RECT 198.000 463.200 201.600 463.800 ;
        RECT 208.200 463.200 212.400 463.800 ;
        RECT 219.000 463.200 222.600 463.800 ;
        RECT 186.600 462.600 195.600 463.200 ;
        RECT 198.000 462.600 202.200 463.200 ;
        RECT 48.600 462.000 52.200 462.600 ;
        RECT 49.200 461.400 52.200 462.000 ;
        RECT 88.800 461.400 91.800 462.600 ;
        RECT 113.400 462.000 117.600 462.600 ;
        RECT 49.200 460.800 52.800 461.400 ;
        RECT 49.800 460.200 52.800 460.800 ;
        RECT 88.200 460.800 91.800 461.400 ;
        RECT 112.800 461.400 117.000 462.000 ;
        RECT 112.800 460.800 116.400 461.400 ;
        RECT 49.800 459.600 53.400 460.200 ;
        RECT 50.400 459.000 54.000 459.600 ;
        RECT 88.200 459.000 91.200 460.800 ;
        RECT 112.200 460.200 115.800 460.800 ;
        RECT 111.600 459.000 115.200 460.200 ;
        RECT 120.000 459.600 123.000 462.600 ;
        RECT 157.800 462.000 164.400 462.600 ;
        RECT 170.400 462.000 174.600 462.600 ;
        RECT 156.000 461.400 159.600 462.000 ;
        RECT 161.400 461.400 165.000 462.000 ;
        RECT 171.000 461.400 175.200 462.000 ;
        RECT 154.800 460.800 159.000 461.400 ;
        RECT 162.600 460.800 165.000 461.400 ;
        RECT 171.600 460.800 175.800 461.400 ;
        RECT 154.200 460.200 158.400 460.800 ;
        RECT 153.000 459.600 157.800 460.200 ;
        RECT 172.200 459.600 175.800 460.800 ;
        RECT 120.000 459.000 122.400 459.600 ;
        RECT 152.400 459.000 156.600 459.600 ;
        RECT 171.600 459.000 175.800 459.600 ;
        RECT 177.000 459.000 180.000 462.600 ;
        RECT 186.000 462.000 196.200 462.600 ;
        RECT 198.600 462.000 202.200 462.600 ;
        RECT 207.600 462.600 211.800 463.200 ;
        RECT 219.600 462.600 223.200 463.200 ;
        RECT 207.600 462.000 211.200 462.600 ;
        RECT 186.000 461.400 196.800 462.000 ;
        RECT 199.200 461.400 202.800 462.000 ;
        RECT 207.000 461.400 210.600 462.000 ;
        RECT 220.200 461.400 223.800 462.600 ;
        RECT 185.400 460.800 197.400 461.400 ;
        RECT 184.800 460.200 192.600 460.800 ;
        RECT 193.800 460.200 198.000 460.800 ;
        RECT 199.800 460.200 203.400 461.400 ;
        RECT 206.400 460.200 210.000 461.400 ;
        RECT 220.800 460.800 223.800 461.400 ;
        RECT 184.200 459.600 187.800 460.200 ;
        RECT 183.000 459.000 187.800 459.600 ;
        RECT 189.000 459.000 192.000 460.200 ;
        RECT 194.400 459.600 198.600 460.200 ;
        RECT 200.400 459.600 204.000 460.200 ;
        RECT 205.800 459.600 209.400 460.200 ;
        RECT 195.000 459.000 199.200 459.600 ;
        RECT 201.000 459.000 204.600 459.600 ;
        RECT 205.800 459.000 208.800 459.600 ;
        RECT 221.400 459.000 224.400 460.800 ;
        RECT 51.000 458.400 54.000 459.000 ;
        RECT 51.000 457.800 54.600 458.400 ;
        RECT 51.600 456.600 55.200 457.800 ;
        RECT 52.200 456.000 55.800 456.600 ;
        RECT 87.600 456.000 90.600 459.000 ;
        RECT 111.000 458.400 114.600 459.000 ;
        RECT 110.400 457.800 114.000 458.400 ;
        RECT 110.400 457.200 113.400 457.800 ;
        RECT 109.800 456.600 113.400 457.200 ;
        RECT 109.800 456.000 112.800 456.600 ;
        RECT 52.800 454.800 56.400 456.000 ;
        RECT 53.400 454.200 57.000 454.800 ;
        RECT 54.000 453.000 57.600 454.200 ;
        RECT 54.600 452.400 58.200 453.000 ;
        RECT 55.200 451.200 58.800 452.400 ;
        RECT 87.000 451.200 90.000 456.000 ;
        RECT 109.200 455.400 112.800 456.000 ;
        RECT 119.400 455.400 122.400 459.000 ;
        RECT 151.800 458.400 156.000 459.000 ;
        RECT 171.000 458.400 175.200 459.000 ;
        RECT 177.000 458.400 187.200 459.000 ;
        RECT 151.200 457.800 155.400 458.400 ;
        RECT 171.000 457.800 174.600 458.400 ;
        RECT 177.600 457.800 186.600 458.400 ;
        RECT 150.000 457.200 154.800 457.800 ;
        RECT 170.400 457.200 174.000 457.800 ;
        RECT 177.600 457.200 185.400 457.800 ;
        RECT 149.400 456.600 154.200 457.200 ;
        RECT 169.800 456.600 174.000 457.200 ;
        RECT 178.200 456.600 184.800 457.200 ;
        RECT 188.400 456.600 192.000 459.000 ;
        RECT 195.600 458.400 199.800 459.000 ;
        RECT 201.600 458.400 208.800 459.000 ;
        RECT 196.200 457.800 200.400 458.400 ;
        RECT 201.600 457.800 208.200 458.400 ;
        RECT 196.800 457.200 201.000 457.800 ;
        RECT 148.800 456.000 153.000 456.600 ;
        RECT 169.800 456.000 173.400 456.600 ;
        RECT 179.400 456.000 183.600 456.600 ;
        RECT 148.800 455.400 152.400 456.000 ;
        RECT 169.800 455.400 172.800 456.000 ;
        RECT 109.200 454.800 112.200 455.400 ;
        RECT 108.600 454.200 112.200 454.800 ;
        RECT 120.000 454.800 122.400 455.400 ;
        RECT 148.200 454.800 151.800 455.400 ;
        RECT 169.200 454.800 172.800 455.400 ;
        RECT 189.000 454.800 192.000 456.600 ;
        RECT 197.400 456.600 201.000 457.200 ;
        RECT 202.200 457.200 208.200 457.800 ;
        RECT 202.200 456.600 207.600 457.200 ;
        RECT 197.400 456.000 207.600 456.600 ;
        RECT 198.000 455.400 207.600 456.000 ;
        RECT 198.600 454.800 207.000 455.400 ;
        RECT 108.600 453.600 111.600 454.200 ;
        RECT 108.000 453.000 111.600 453.600 ;
        RECT 108.000 452.400 111.000 453.000 ;
        RECT 120.000 452.400 123.000 454.800 ;
        RECT 147.600 454.200 151.200 454.800 ;
        RECT 147.000 453.600 150.600 454.200 ;
        RECT 146.400 453.000 150.000 453.600 ;
        RECT 169.200 453.000 172.200 454.800 ;
        RECT 145.800 452.400 150.000 453.000 ;
        RECT 155.400 452.400 156.000 453.000 ;
        RECT 55.800 450.600 59.400 451.200 ;
        RECT 87.600 450.600 90.000 451.200 ;
        RECT 107.400 451.800 111.000 452.400 ;
        RECT 107.400 450.600 110.400 451.800 ;
        RECT 56.400 449.400 60.000 450.600 ;
        RECT 57.000 448.800 60.600 449.400 ;
        RECT 57.600 447.600 61.200 448.800 ;
        RECT 87.600 448.200 90.600 450.600 ;
        RECT 106.800 450.000 110.400 450.600 ;
        RECT 120.600 450.600 123.000 452.400 ;
        RECT 145.200 451.800 149.400 452.400 ;
        RECT 145.200 451.200 148.800 451.800 ;
        RECT 155.400 451.200 156.600 452.400 ;
        RECT 168.600 451.200 172.200 453.000 ;
        RECT 189.000 454.200 194.400 454.800 ;
        RECT 189.000 453.600 195.000 454.200 ;
        RECT 199.200 453.600 207.000 454.800 ;
        RECT 189.000 453.000 195.600 453.600 ;
        RECT 199.800 453.000 206.400 453.600 ;
        RECT 222.000 453.000 225.000 459.000 ;
        RECT 189.000 452.400 196.800 453.000 ;
        RECT 189.000 451.800 197.400 452.400 ;
        RECT 189.600 451.200 197.400 451.800 ;
        RECT 200.400 451.800 204.000 453.000 ;
        RECT 200.400 451.200 204.600 451.800 ;
        RECT 221.400 451.200 224.400 453.000 ;
        RECT 144.600 450.600 148.200 451.200 ;
        RECT 106.800 448.800 109.800 450.000 ;
        RECT 120.600 448.800 123.600 450.600 ;
        RECT 144.000 449.400 147.600 450.600 ;
        RECT 155.400 450.000 157.200 451.200 ;
        RECT 143.400 448.800 147.000 449.400 ;
        RECT 155.400 448.800 157.800 450.000 ;
        RECT 106.200 448.200 109.800 448.800 ;
        RECT 58.200 447.000 61.800 447.600 ;
        RECT 58.800 446.400 62.400 447.000 ;
        RECT 88.200 446.400 91.200 448.200 ;
        RECT 106.200 446.400 109.200 448.200 ;
        RECT 121.200 447.600 123.600 448.800 ;
        RECT 142.800 448.200 146.400 448.800 ;
        RECT 156.000 448.200 157.800 448.800 ;
        RECT 142.800 447.600 145.800 448.200 ;
        RECT 59.400 445.200 63.000 446.400 ;
        RECT 88.800 445.200 91.800 446.400 ;
        RECT 60.000 444.600 63.600 445.200 ;
        RECT 88.800 444.600 92.400 445.200 ;
        RECT 60.600 444.000 64.200 444.600 ;
        RECT 89.400 444.000 93.000 444.600 ;
        RECT 60.600 443.400 64.800 444.000 ;
        RECT 61.200 442.800 64.800 443.400 ;
        RECT 90.000 443.400 93.000 444.000 ;
        RECT 90.000 442.800 93.600 443.400 ;
        RECT 61.800 442.200 65.400 442.800 ;
        RECT 90.600 442.200 94.200 442.800 ;
        RECT 62.400 441.600 66.000 442.200 ;
        RECT 90.600 441.600 94.800 442.200 ;
        RECT 63.000 441.000 66.600 441.600 ;
        RECT 91.200 441.000 95.400 441.600 ;
        RECT 63.000 440.400 67.200 441.000 ;
        RECT 91.800 440.400 96.000 441.000 ;
        RECT 63.600 439.800 67.200 440.400 ;
        RECT 92.400 439.800 96.600 440.400 ;
        RECT 64.200 439.200 67.800 439.800 ;
        RECT 93.000 439.200 97.200 439.800 ;
        RECT 64.800 438.600 68.400 439.200 ;
        RECT 93.000 438.600 97.800 439.200 ;
        RECT 64.800 438.000 69.000 438.600 ;
        RECT 93.000 438.000 98.400 438.600 ;
        RECT 65.400 437.400 69.600 438.000 ;
        RECT 66.000 436.800 69.600 437.400 ;
        RECT 92.400 437.400 99.600 438.000 ;
        RECT 105.600 437.400 108.600 446.400 ;
        RECT 121.200 445.800 124.200 447.600 ;
        RECT 142.200 447.000 145.800 447.600 ;
        RECT 142.200 446.400 145.200 447.000 ;
        RECT 141.600 445.800 145.200 446.400 ;
        RECT 156.000 445.800 158.400 448.200 ;
        RECT 121.800 444.000 124.800 445.800 ;
        RECT 141.000 445.200 144.600 445.800 ;
        RECT 141.000 444.600 144.000 445.200 ;
        RECT 140.400 444.000 144.000 444.600 ;
        RECT 121.800 443.400 125.400 444.000 ;
        RECT 140.400 443.400 143.400 444.000 ;
        RECT 122.400 442.200 125.400 443.400 ;
        RECT 139.800 442.800 143.400 443.400 ;
        RECT 122.400 441.600 126.000 442.200 ;
        RECT 139.800 441.600 142.800 442.800 ;
        RECT 123.000 440.400 126.000 441.600 ;
        RECT 139.200 440.400 142.200 441.600 ;
        RECT 123.600 439.200 126.600 440.400 ;
        RECT 138.600 439.800 142.200 440.400 ;
        RECT 138.600 439.200 141.600 439.800 ;
        RECT 123.600 438.600 127.200 439.200 ;
        RECT 92.400 436.800 100.800 437.400 ;
        RECT 66.600 436.200 70.200 436.800 ;
        RECT 92.400 436.200 102.000 436.800 ;
        RECT 67.200 435.600 70.800 436.200 ;
        RECT 92.400 435.600 95.400 436.200 ;
        RECT 97.200 435.600 103.200 436.200 ;
        RECT 106.200 435.600 108.600 437.400 ;
        RECT 123.000 438.000 127.200 438.600 ;
        RECT 138.000 438.600 141.600 439.200 ;
        RECT 123.000 437.400 127.800 438.000 ;
        RECT 138.000 437.400 141.000 438.600 ;
        RECT 123.000 436.800 128.400 437.400 ;
        RECT 122.400 436.200 128.400 436.800 ;
        RECT 137.400 436.200 140.400 437.400 ;
        RECT 156.000 436.800 159.000 445.800 ;
        RECT 168.600 442.200 171.600 451.200 ;
        RECT 189.600 450.600 198.000 451.200 ;
        RECT 189.600 450.000 198.600 450.600 ;
        RECT 201.000 450.000 204.600 451.200 ;
        RECT 220.800 450.600 224.400 451.200 ;
        RECT 220.800 450.000 223.800 450.600 ;
        RECT 189.600 448.200 193.200 450.000 ;
        RECT 194.400 449.400 199.200 450.000 ;
        RECT 195.000 448.800 199.800 449.400 ;
        RECT 201.600 448.800 205.200 450.000 ;
        RECT 220.200 449.400 223.800 450.000 ;
        RECT 220.200 448.800 223.200 449.400 ;
        RECT 195.600 448.200 200.400 448.800 ;
        RECT 189.600 447.600 193.800 448.200 ;
        RECT 196.200 447.600 200.400 448.200 ;
        RECT 202.200 448.200 205.800 448.800 ;
        RECT 219.600 448.200 223.200 448.800 ;
        RECT 202.200 447.600 206.400 448.200 ;
        RECT 219.000 447.600 224.400 448.200 ;
        RECT 190.200 445.800 193.800 447.600 ;
        RECT 196.800 447.000 201.000 447.600 ;
        RECT 202.800 447.000 206.400 447.600 ;
        RECT 217.200 447.000 226.200 447.600 ;
        RECT 197.400 446.400 201.600 447.000 ;
        RECT 203.400 446.400 207.000 447.000 ;
        RECT 216.000 446.400 226.800 447.000 ;
        RECT 197.400 445.800 202.200 446.400 ;
        RECT 190.800 445.200 193.800 445.800 ;
        RECT 198.000 445.200 202.200 445.800 ;
        RECT 204.000 445.800 207.600 446.400 ;
        RECT 216.000 445.800 227.400 446.400 ;
        RECT 204.000 445.200 208.200 445.800 ;
        RECT 190.800 444.000 194.400 445.200 ;
        RECT 198.600 444.600 202.800 445.200 ;
        RECT 204.600 444.600 208.200 445.200 ;
        RECT 216.000 445.200 228.000 445.800 ;
        RECT 216.000 444.600 220.200 445.200 ;
        RECT 224.400 444.600 228.000 445.200 ;
        RECT 191.400 443.400 194.400 444.000 ;
        RECT 199.200 443.400 203.400 444.600 ;
        RECT 205.200 444.000 208.800 444.600 ;
        RECT 205.800 443.400 209.400 444.000 ;
        RECT 191.400 442.800 195.000 443.400 ;
        RECT 199.800 442.800 204.000 443.400 ;
        RECT 205.800 442.800 210.000 443.400 ;
        RECT 225.000 442.800 228.000 444.600 ;
        RECT 192.000 442.200 195.000 442.800 ;
        RECT 200.400 442.200 204.000 442.800 ;
        RECT 206.400 442.200 210.000 442.800 ;
        RECT 224.400 442.200 228.000 442.800 ;
        RECT 168.600 441.000 171.000 442.200 ;
        RECT 192.000 441.600 195.600 442.200 ;
        RECT 200.400 441.600 204.600 442.200 ;
        RECT 207.000 441.600 210.600 442.200 ;
        RECT 224.400 441.600 227.400 442.200 ;
        RECT 156.000 436.200 158.400 436.800 ;
        RECT 122.400 435.600 129.000 436.200 ;
        RECT 136.800 435.600 140.400 436.200 ;
        RECT 67.800 435.000 71.400 435.600 ;
        RECT 67.800 434.400 72.000 435.000 ;
        RECT 68.400 433.800 72.600 434.400 ;
        RECT 69.000 433.200 73.200 433.800 ;
        RECT 69.600 432.600 73.800 433.200 ;
        RECT 70.200 432.000 73.800 432.600 ;
        RECT 70.800 431.400 74.400 432.000 ;
        RECT 71.400 430.800 75.000 431.400 ;
        RECT 72.000 430.200 75.600 430.800 ;
        RECT 72.000 429.600 76.200 430.200 ;
        RECT 72.600 429.000 76.800 429.600 ;
        RECT 73.200 428.400 77.400 429.000 ;
        RECT 73.800 427.800 78.000 428.400 ;
        RECT 74.400 427.200 78.600 427.800 ;
        RECT 75.000 426.600 79.200 427.200 ;
        RECT 75.600 426.000 79.800 426.600 ;
        RECT 76.200 425.400 80.400 426.000 ;
        RECT 76.800 424.800 81.000 425.400 ;
        RECT 77.400 424.200 81.600 424.800 ;
        RECT 91.800 424.200 94.800 435.600 ;
        RECT 97.800 435.000 104.400 435.600 ;
        RECT 106.200 435.000 109.200 435.600 ;
        RECT 121.800 435.000 129.600 435.600 ;
        RECT 136.800 435.000 139.800 435.600 ;
        RECT 99.000 434.400 109.200 435.000 ;
        RECT 100.200 433.800 109.200 434.400 ;
        RECT 121.200 433.800 124.800 435.000 ;
        RECT 126.000 434.400 130.200 435.000 ;
        RECT 136.200 434.400 139.800 435.000 ;
        RECT 126.600 433.800 130.800 434.400 ;
        RECT 135.600 433.800 139.200 434.400 ;
        RECT 155.400 433.800 158.400 436.200 ;
        RECT 168.000 436.200 171.000 441.000 ;
        RECT 192.600 441.000 195.600 441.600 ;
        RECT 201.000 441.000 205.200 441.600 ;
        RECT 207.600 441.000 211.200 441.600 ;
        RECT 223.800 441.000 227.400 441.600 ;
        RECT 192.600 440.400 196.200 441.000 ;
        RECT 201.600 440.400 205.200 441.000 ;
        RECT 208.200 440.400 211.200 441.000 ;
        RECT 223.200 440.400 226.800 441.000 ;
        RECT 193.200 439.800 196.200 440.400 ;
        RECT 193.200 439.200 196.800 439.800 ;
        RECT 202.200 439.200 205.800 440.400 ;
        RECT 208.800 439.800 211.800 440.400 ;
        RECT 222.600 439.800 226.800 440.400 ;
        RECT 210.000 439.200 211.800 439.800 ;
        RECT 222.000 439.200 226.200 439.800 ;
        RECT 193.800 438.600 196.800 439.200 ;
        RECT 202.800 438.600 205.800 439.200 ;
        RECT 210.600 438.600 211.800 439.200 ;
        RECT 221.400 438.600 225.600 439.200 ;
        RECT 193.800 438.000 197.400 438.600 ;
        RECT 202.800 438.000 206.400 438.600 ;
        RECT 220.200 438.000 225.600 438.600 ;
        RECT 228.600 438.000 231.600 438.600 ;
        RECT 194.400 436.800 198.000 438.000 ;
        RECT 203.400 436.800 206.400 438.000 ;
        RECT 219.600 437.400 232.200 438.000 ;
        RECT 218.400 436.800 232.800 437.400 ;
        RECT 195.000 436.200 198.600 436.800 ;
        RECT 168.000 435.600 170.400 436.200 ;
        RECT 101.400 433.200 109.200 433.800 ;
        RECT 102.600 432.600 108.600 433.200 ;
        RECT 120.600 432.600 124.200 433.800 ;
        RECT 127.200 433.200 131.400 433.800 ;
        RECT 135.000 433.200 139.200 433.800 ;
        RECT 127.800 432.600 132.600 433.200 ;
        RECT 134.400 432.600 138.600 433.200 ;
        RECT 104.400 432.000 108.000 432.600 ;
        RECT 120.000 431.400 123.600 432.600 ;
        RECT 128.400 432.000 138.000 432.600 ;
        RECT 154.800 432.000 157.800 433.800 ;
        RECT 129.000 431.400 137.400 432.000 ;
        RECT 119.400 430.200 123.000 431.400 ;
        RECT 129.600 430.800 136.800 431.400 ;
        RECT 130.800 430.200 136.200 430.800 ;
        RECT 154.200 430.200 157.800 432.000 ;
        RECT 167.400 430.200 170.400 435.600 ;
        RECT 195.600 435.000 199.200 436.200 ;
        RECT 196.200 434.400 199.800 435.000 ;
        RECT 196.800 433.800 200.400 434.400 ;
        RECT 203.400 433.800 207.000 436.800 ;
        RECT 217.200 436.200 233.400 436.800 ;
        RECT 216.600 435.600 233.400 436.200 ;
        RECT 216.600 435.000 228.600 435.600 ;
        RECT 218.400 434.400 226.200 435.000 ;
        RECT 230.400 434.400 233.400 435.600 ;
        RECT 197.400 433.200 201.000 433.800 ;
        RECT 202.800 433.200 207.000 433.800 ;
        RECT 197.400 432.600 206.400 433.200 ;
        RECT 198.000 432.000 206.400 432.600 ;
        RECT 199.200 431.400 207.600 432.000 ;
        RECT 200.400 430.800 209.400 431.400 ;
        RECT 204.000 430.200 210.600 430.800 ;
        RECT 118.800 429.000 122.400 430.200 ;
        RECT 132.600 429.600 134.400 430.200 ;
        RECT 153.600 429.600 158.400 430.200 ;
        RECT 167.400 429.600 169.800 430.200 ;
        RECT 205.800 429.600 212.400 430.200 ;
        RECT 153.600 429.000 159.000 429.600 ;
        RECT 118.200 428.400 122.400 429.000 ;
        RECT 153.000 428.400 159.600 429.000 ;
        RECT 118.200 427.800 123.000 428.400 ;
        RECT 117.600 427.200 123.000 427.800 ;
        RECT 153.000 427.800 160.200 428.400 ;
        RECT 153.000 427.200 161.400 427.800 ;
        RECT 117.000 426.000 123.600 427.200 ;
        RECT 152.400 426.000 155.400 427.200 ;
        RECT 157.200 426.600 162.000 427.200 ;
        RECT 157.800 426.000 163.200 426.600 ;
        RECT 116.400 425.400 120.000 426.000 ;
        RECT 115.800 424.800 119.400 425.400 ;
        RECT 115.200 424.200 118.800 424.800 ;
        RECT 121.200 424.200 124.200 426.000 ;
        RECT 151.800 425.400 155.400 426.000 ;
        RECT 159.000 425.400 164.400 426.000 ;
        RECT 151.800 424.800 154.800 425.400 ;
        RECT 159.600 424.800 165.600 425.400 ;
        RECT 166.800 424.800 169.800 429.600 ;
        RECT 207.600 429.000 213.600 429.600 ;
        RECT 209.400 428.400 214.800 429.000 ;
        RECT 210.600 427.800 216.600 428.400 ;
        RECT 231.000 427.800 234.000 434.400 ;
        RECT 211.800 427.200 217.800 427.800 ;
        RECT 213.600 426.600 219.000 427.200 ;
        RECT 214.800 426.000 220.200 426.600 ;
        RECT 216.000 425.400 221.400 426.000 ;
        RECT 230.400 425.400 233.400 427.800 ;
        RECT 535.800 426.000 546.600 426.600 ;
        RECT 529.800 425.400 553.800 426.000 ;
        RECT 217.200 424.800 222.600 425.400 ;
        RECT 151.200 424.200 154.800 424.800 ;
        RECT 160.200 424.200 169.800 424.800 ;
        RECT 219.000 424.200 223.800 424.800 ;
        RECT 229.800 424.200 232.800 425.400 ;
        RECT 526.800 424.800 558.600 425.400 ;
        RECT 524.400 424.200 562.200 424.800 ;
        RECT 78.000 423.600 82.200 424.200 ;
        RECT 92.400 423.600 94.800 424.200 ;
        RECT 114.600 423.600 118.800 424.200 ;
        RECT 78.600 423.000 82.800 423.600 ;
        RECT 79.200 422.400 83.400 423.000 ;
        RECT 79.800 421.800 84.000 422.400 ;
        RECT 92.400 421.800 95.400 423.600 ;
        RECT 114.600 423.000 118.200 423.600 ;
        RECT 114.000 422.400 117.600 423.000 ;
        RECT 113.400 421.800 117.000 422.400 ;
        RECT 121.800 421.800 124.800 424.200 ;
        RECT 150.600 423.600 154.800 424.200 ;
        RECT 161.400 423.600 169.800 424.200 ;
        RECT 220.200 423.600 224.400 424.200 ;
        RECT 229.200 423.600 232.800 424.200 ;
        RECT 522.000 423.600 565.200 424.200 ;
        RECT 150.600 423.000 155.400 423.600 ;
        RECT 162.600 423.000 169.800 423.600 ;
        RECT 221.400 423.000 225.600 423.600 ;
        RECT 228.600 423.000 232.200 423.600 ;
        RECT 520.200 423.000 534.600 423.600 ;
        RECT 547.800 423.000 567.600 423.600 ;
        RECT 150.000 422.400 155.400 423.000 ;
        RECT 163.200 422.400 169.800 423.000 ;
        RECT 222.000 422.400 226.800 423.000 ;
        RECT 228.000 422.400 232.200 423.000 ;
        RECT 518.400 422.400 529.800 423.000 ;
        RECT 554.400 422.400 570.600 423.000 ;
        RECT 150.000 421.800 156.000 422.400 ;
        RECT 163.200 421.800 169.200 422.400 ;
        RECT 223.200 421.800 231.600 422.400 ;
        RECT 516.600 421.800 526.800 422.400 ;
        RECT 558.600 421.800 572.400 422.400 ;
        RECT 80.400 421.200 84.600 421.800 ;
        RECT 92.400 421.200 96.000 421.800 ;
        RECT 112.800 421.200 116.400 421.800 ;
        RECT 81.000 420.600 85.200 421.200 ;
        RECT 81.600 420.000 85.800 420.600 ;
        RECT 93.000 420.000 96.000 421.200 ;
        RECT 112.200 420.600 116.400 421.200 ;
        RECT 111.600 420.000 115.800 420.600 ;
        RECT 82.200 419.400 86.400 420.000 ;
        RECT 93.000 419.400 96.600 420.000 ;
        RECT 82.800 418.800 87.000 419.400 ;
        RECT 93.600 418.800 96.600 419.400 ;
        RECT 111.000 419.400 115.200 420.000 ;
        RECT 111.000 418.800 114.600 419.400 ;
        RECT 122.400 418.800 125.400 421.800 ;
        RECT 149.400 421.200 156.000 421.800 ;
        RECT 148.800 420.600 156.000 421.200 ;
        RECT 163.800 421.200 168.600 421.800 ;
        RECT 224.400 421.200 231.000 421.800 ;
        RECT 515.400 421.200 524.400 421.800 ;
        RECT 562.200 421.200 574.200 421.800 ;
        RECT 163.800 420.600 168.000 421.200 ;
        RECT 225.000 420.600 229.800 421.200 ;
        RECT 514.200 420.600 522.000 421.200 ;
        RECT 565.200 420.600 576.000 421.200 ;
        RECT 148.800 420.000 156.600 420.600 ;
        RECT 164.400 420.000 168.000 420.600 ;
        RECT 226.200 420.000 229.800 420.600 ;
        RECT 513.000 420.000 520.200 420.600 ;
        RECT 567.600 420.000 577.800 420.600 ;
        RECT 148.200 419.400 156.600 420.000 ;
        RECT 83.400 418.200 88.200 418.800 ;
        RECT 93.600 418.200 97.200 418.800 ;
        RECT 110.400 418.200 114.000 418.800 ;
        RECT 84.000 417.600 88.800 418.200 ;
        RECT 94.200 417.600 97.200 418.200 ;
        RECT 109.800 417.600 113.400 418.200 ;
        RECT 84.600 417.000 89.400 417.600 ;
        RECT 94.200 417.000 97.800 417.600 ;
        RECT 109.200 417.000 112.800 417.600 ;
        RECT 85.800 416.400 90.000 417.000 ;
        RECT 94.800 416.400 97.800 417.000 ;
        RECT 108.600 416.400 112.200 417.000 ;
        RECT 86.400 415.800 90.600 416.400 ;
        RECT 94.800 415.800 98.400 416.400 ;
        RECT 108.000 415.800 112.200 416.400 ;
        RECT 123.000 415.800 126.000 418.800 ;
        RECT 147.600 418.200 151.200 419.400 ;
        RECT 152.400 418.800 156.600 419.400 ;
        RECT 165.000 419.400 168.000 420.000 ;
        RECT 226.800 419.400 229.800 420.000 ;
        RECT 511.200 419.400 519.000 420.000 ;
        RECT 570.000 419.400 579.000 420.000 ;
        RECT 165.000 418.800 168.600 419.400 ;
        RECT 227.400 418.800 230.400 419.400 ;
        RECT 510.600 418.800 517.200 419.400 ;
        RECT 571.800 418.800 580.200 419.400 ;
        RECT 153.000 418.200 156.600 418.800 ;
        RECT 165.600 418.200 169.200 418.800 ;
        RECT 228.000 418.200 231.000 418.800 ;
        RECT 509.400 418.200 516.000 418.800 ;
        RECT 573.600 418.200 582.000 418.800 ;
        RECT 147.000 417.600 150.600 418.200 ;
        RECT 153.000 417.600 157.200 418.200 ;
        RECT 146.400 416.400 150.000 417.600 ;
        RECT 145.800 415.800 149.400 416.400 ;
        RECT 87.000 415.200 91.800 415.800 ;
        RECT 95.400 415.200 99.000 415.800 ;
        RECT 107.400 415.200 111.600 415.800 ;
        RECT 87.600 414.600 92.400 415.200 ;
        RECT 96.000 414.600 99.000 415.200 ;
        RECT 106.800 414.600 111.000 415.200 ;
        RECT 87.600 414.000 93.000 414.600 ;
        RECT 96.000 414.000 99.600 414.600 ;
        RECT 106.200 414.000 110.400 414.600 ;
        RECT 87.600 413.400 94.200 414.000 ;
        RECT 96.600 413.400 100.200 414.000 ;
        RECT 105.600 413.400 109.800 414.000 ;
        RECT 86.400 412.800 94.800 413.400 ;
        RECT 97.200 412.800 101.400 413.400 ;
        RECT 104.400 412.800 108.600 413.400 ;
        RECT 123.600 412.800 126.600 415.800 ;
        RECT 145.200 414.600 148.800 415.800 ;
        RECT 153.600 415.200 157.200 417.600 ;
        RECT 166.200 417.600 169.200 418.200 ;
        RECT 228.600 417.600 231.000 418.200 ;
        RECT 508.200 417.600 514.200 418.200 ;
        RECT 575.400 417.600 583.200 418.200 ;
        RECT 166.200 417.000 169.800 417.600 ;
        RECT 228.600 417.000 231.600 417.600 ;
        RECT 507.000 417.000 513.000 417.600 ;
        RECT 576.600 417.000 584.400 417.600 ;
        RECT 166.800 416.400 169.800 417.000 ;
        RECT 167.400 415.800 169.800 416.400 ;
        RECT 229.200 416.400 231.600 417.000 ;
        RECT 506.400 416.400 511.800 417.000 ;
        RECT 578.400 416.400 586.200 417.000 ;
        RECT 229.200 415.800 232.200 416.400 ;
        RECT 505.200 415.800 511.200 416.400 ;
        RECT 579.600 415.800 587.400 416.400 ;
        RECT 168.000 415.200 170.400 415.800 ;
        RECT 144.600 414.000 148.200 414.600 ;
        RECT 154.200 414.000 157.200 415.200 ;
        RECT 168.600 414.600 169.800 415.200 ;
        RECT 229.800 414.600 232.200 415.800 ;
        RECT 504.000 415.200 510.000 415.800 ;
        RECT 581.400 415.200 588.600 415.800 ;
        RECT 503.400 414.600 508.800 415.200 ;
        RECT 582.600 414.600 589.800 415.200 ;
        RECT 230.400 414.000 232.200 414.600 ;
        RECT 502.200 414.000 507.600 414.600 ;
        RECT 584.400 414.000 591.000 414.600 ;
        RECT 144.000 413.400 147.600 414.000 ;
        RECT 85.800 412.200 95.400 412.800 ;
        RECT 97.800 412.200 108.000 412.800 ;
        RECT 124.200 412.200 126.600 412.800 ;
        RECT 143.400 412.200 147.000 413.400 ;
        RECT 84.600 411.600 89.400 412.200 ;
        RECT 91.200 411.600 96.600 412.200 ;
        RECT 98.400 411.600 107.400 412.200 ;
        RECT 84.000 411.000 88.800 411.600 ;
        RECT 92.400 411.000 97.200 411.600 ;
        RECT 99.000 411.000 106.800 411.600 ;
        RECT 82.800 410.400 88.200 411.000 ;
        RECT 93.000 410.400 98.400 411.000 ;
        RECT 99.600 410.400 106.200 411.000 ;
        RECT 81.600 409.800 87.000 410.400 ;
        RECT 94.200 409.800 99.000 410.400 ;
        RECT 101.400 409.800 105.000 410.400 ;
        RECT 81.000 409.200 86.400 409.800 ;
        RECT 94.800 409.200 99.600 409.800 ;
        RECT 101.400 409.200 104.400 409.800 ;
        RECT 124.200 409.200 127.200 412.200 ;
        RECT 142.800 411.600 146.400 412.200 ;
        RECT 142.200 411.000 145.800 411.600 ;
        RECT 141.600 410.400 145.200 411.000 ;
        RECT 141.000 409.800 145.200 410.400 ;
        RECT 141.000 409.200 144.600 409.800 ;
        RECT 79.800 408.600 85.200 409.200 ;
        RECT 96.000 408.600 104.400 409.200 ;
        RECT 78.600 408.000 84.600 408.600 ;
        RECT 96.600 408.000 104.400 408.600 ;
        RECT 78.000 407.400 83.400 408.000 ;
        RECT 97.800 407.400 104.400 408.000 ;
        RECT 76.800 406.800 82.200 407.400 ;
        RECT 98.400 406.800 104.400 407.400 ;
        RECT 76.200 406.200 81.600 406.800 ;
        RECT 99.600 406.200 104.400 406.800 ;
        RECT 75.000 405.600 80.400 406.200 ;
        RECT 100.800 405.600 104.400 406.200 ;
        RECT 124.800 408.600 127.200 409.200 ;
        RECT 140.400 408.600 144.000 409.200 ;
        RECT 154.200 408.600 157.800 414.000 ;
        RECT 230.400 409.800 232.800 414.000 ;
        RECT 501.600 413.400 507.000 414.000 ;
        RECT 585.600 413.400 592.200 414.000 ;
        RECT 501.000 412.800 505.800 413.400 ;
        RECT 586.800 412.800 593.400 413.400 ;
        RECT 500.400 412.200 505.200 412.800 ;
        RECT 588.000 412.200 594.600 412.800 ;
        RECT 499.800 411.600 504.000 412.200 ;
        RECT 589.200 411.600 595.800 412.200 ;
        RECT 499.200 411.000 503.400 411.600 ;
        RECT 590.400 411.000 597.000 411.600 ;
        RECT 498.000 410.400 502.800 411.000 ;
        RECT 591.600 410.400 598.200 411.000 ;
        RECT 497.400 409.800 501.600 410.400 ;
        RECT 592.800 409.800 599.400 410.400 ;
        RECT 231.000 408.600 232.800 409.800 ;
        RECT 496.800 409.200 501.000 409.800 ;
        RECT 594.000 409.200 600.600 409.800 ;
        RECT 496.200 408.600 500.400 409.200 ;
        RECT 595.200 408.600 601.200 409.200 ;
        RECT 124.800 405.600 127.800 408.600 ;
        RECT 139.800 408.000 143.400 408.600 ;
        RECT 139.200 407.400 142.800 408.000 ;
        RECT 154.200 407.400 157.200 408.600 ;
        RECT 138.600 406.800 142.800 407.400 ;
        RECT 138.000 406.200 142.200 406.800 ;
        RECT 137.400 405.600 141.600 406.200 ;
        RECT 153.600 405.600 157.200 407.400 ;
        RECT 73.800 405.000 79.800 405.600 ;
        RECT 73.200 404.400 78.600 405.000 ;
        RECT 72.000 403.800 77.400 404.400 ;
        RECT 71.400 403.200 76.800 403.800 ;
        RECT 70.200 402.600 75.600 403.200 ;
        RECT 69.600 402.000 75.000 402.600 ;
        RECT 68.400 401.400 73.800 402.000 ;
        RECT 67.800 400.800 73.200 401.400 ;
        RECT 66.600 400.200 72.000 400.800 ;
        RECT 66.000 399.600 71.400 400.200 ;
        RECT 64.800 399.000 70.200 399.600 ;
        RECT 64.200 398.400 69.600 399.000 ;
        RECT 63.600 397.800 68.400 398.400 ;
        RECT 62.400 397.200 67.800 397.800 ;
        RECT 61.800 396.600 66.600 397.200 ;
        RECT 101.400 396.600 104.400 405.600 ;
        RECT 125.400 403.800 128.400 405.600 ;
        RECT 136.800 405.000 141.600 405.600 ;
        RECT 153.000 405.000 156.600 405.600 ;
        RECT 136.200 404.400 142.200 405.000 ;
        RECT 152.400 404.400 156.600 405.000 ;
        RECT 135.600 403.800 142.800 404.400 ;
        RECT 152.400 403.800 156.000 404.400 ;
        RECT 126.000 402.600 129.000 403.800 ;
        RECT 135.000 403.200 143.400 403.800 ;
        RECT 151.200 403.200 156.000 403.800 ;
        RECT 134.400 402.600 144.600 403.200 ;
        RECT 150.600 402.600 155.400 403.200 ;
        RECT 126.000 402.000 129.600 402.600 ;
        RECT 133.200 402.000 138.000 402.600 ;
        RECT 139.200 402.000 146.400 402.600 ;
        RECT 148.200 402.000 154.800 402.600 ;
        RECT 230.400 402.000 232.800 408.600 ;
        RECT 495.600 408.000 499.200 408.600 ;
        RECT 596.400 408.000 602.400 408.600 ;
        RECT 495.000 407.400 498.600 408.000 ;
        RECT 597.600 407.400 603.600 408.000 ;
        RECT 494.400 406.800 498.000 407.400 ;
        RECT 598.800 406.800 604.800 407.400 ;
        RECT 493.800 406.200 497.400 406.800 ;
        RECT 599.400 406.200 606.000 406.800 ;
        RECT 493.200 405.600 496.800 406.200 ;
        RECT 600.600 405.600 607.200 406.200 ;
        RECT 492.600 405.000 496.200 405.600 ;
        RECT 601.800 405.000 608.400 405.600 ;
        RECT 492.000 404.400 496.200 405.000 ;
        RECT 603.000 404.400 609.600 405.000 ;
        RECT 491.400 403.800 495.600 404.400 ;
        RECT 604.200 403.800 610.800 404.400 ;
        RECT 491.400 403.200 495.000 403.800 ;
        RECT 605.400 403.200 612.000 403.800 ;
        RECT 490.800 402.600 494.400 403.200 ;
        RECT 606.600 402.600 613.200 403.200 ;
        RECT 490.200 402.000 493.800 402.600 ;
        RECT 607.800 402.000 614.400 402.600 ;
        RECT 126.600 401.400 130.800 402.000 ;
        RECT 132.000 401.400 137.400 402.000 ;
        RECT 140.400 401.400 154.200 402.000 ;
        RECT 229.800 401.400 232.800 402.000 ;
        RECT 489.600 401.400 493.800 402.000 ;
        RECT 609.000 401.400 615.000 402.000 ;
        RECT 126.600 400.800 136.800 401.400 ;
        RECT 141.000 400.800 153.600 401.400 ;
        RECT 127.200 400.200 135.600 400.800 ;
        RECT 142.200 400.200 153.000 400.800 ;
        RECT 127.800 399.600 135.000 400.200 ;
        RECT 143.400 399.600 152.400 400.200 ;
        RECT 229.800 399.600 232.200 401.400 ;
        RECT 489.600 400.800 493.200 401.400 ;
        RECT 610.200 400.800 616.200 401.400 ;
        RECT 489.000 400.200 492.600 400.800 ;
        RECT 611.400 400.200 617.400 400.800 ;
        RECT 129.000 399.000 133.800 399.600 ;
        RECT 144.600 399.000 151.200 399.600 ;
        RECT 129.600 397.800 132.600 399.000 ;
        RECT 147.600 398.400 149.400 399.000 ;
        RECT 229.200 398.400 232.200 399.600 ;
        RECT 488.400 399.000 492.000 400.200 ;
        RECT 612.600 399.600 618.600 400.200 ;
        RECT 613.200 399.000 619.200 399.600 ;
        RECT 487.800 398.400 491.400 399.000 ;
        RECT 614.400 398.400 620.400 399.000 ;
        RECT 60.600 396.000 66.000 396.600 ;
        RECT 60.000 395.400 64.800 396.000 ;
        RECT 58.800 394.800 64.200 395.400 ;
        RECT 58.200 394.200 63.000 394.800 ;
        RECT 57.000 393.600 62.400 394.200 ;
        RECT 102.000 393.600 105.000 396.600 ;
        RECT 130.200 396.000 133.200 397.800 ;
        RECT 229.200 397.200 231.600 398.400 ;
        RECT 487.800 397.800 490.800 398.400 ;
        RECT 615.600 397.800 621.000 398.400 ;
        RECT 487.200 397.200 490.800 397.800 ;
        RECT 616.800 397.200 622.200 397.800 ;
        RECT 228.600 396.600 231.600 397.200 ;
        RECT 486.600 396.600 490.200 397.200 ;
        RECT 617.400 396.600 622.800 397.200 ;
        RECT 130.800 394.200 133.800 396.000 ;
        RECT 225.000 395.400 226.800 396.000 ;
        RECT 228.600 395.400 231.000 396.600 ;
        RECT 486.600 396.000 489.600 396.600 ;
        RECT 534.000 396.000 537.000 396.600 ;
        RECT 618.600 396.000 624.000 396.600 ;
        RECT 222.000 394.800 231.000 395.400 ;
        RECT 486.000 395.400 489.600 396.000 ;
        RECT 529.200 395.400 541.200 396.000 ;
        RECT 619.800 395.400 624.600 396.000 ;
        RECT 486.000 394.800 489.000 395.400 ;
        RECT 526.800 394.800 543.600 395.400 ;
        RECT 620.400 394.800 625.800 395.400 ;
        RECT 220.200 394.200 230.400 394.800 ;
        RECT 56.400 393.000 61.800 393.600 ;
        RECT 55.800 392.400 60.600 393.000 ;
        RECT 102.600 392.400 105.600 393.600 ;
        RECT 131.400 393.000 134.400 394.200 ;
        RECT 218.400 393.600 230.400 394.200 ;
        RECT 485.400 394.200 489.000 394.800 ;
        RECT 525.000 394.200 546.000 394.800 ;
        RECT 621.600 394.200 626.400 394.800 ;
        RECT 485.400 393.600 488.400 394.200 ;
        RECT 523.800 393.600 547.200 394.200 ;
        RECT 622.800 393.600 627.600 394.200 ;
        RECT 217.200 393.000 229.800 393.600 ;
        RECT 131.400 392.400 135.000 393.000 ;
        RECT 216.000 392.400 224.400 393.000 ;
        RECT 226.800 392.400 229.800 393.000 ;
        RECT 484.800 393.000 488.400 393.600 ;
        RECT 522.600 393.000 532.800 393.600 ;
        RECT 537.600 393.000 549.000 393.600 ;
        RECT 623.400 393.000 628.800 393.600 ;
        RECT 484.800 392.400 487.800 393.000 ;
        RECT 521.400 392.400 529.200 393.000 ;
        RECT 541.200 392.400 550.200 393.000 ;
        RECT 624.600 392.400 630.000 393.000 ;
        RECT 54.600 391.800 60.000 392.400 ;
        RECT 79.200 391.800 81.000 392.400 ;
        RECT 102.600 391.800 106.200 392.400 ;
        RECT 54.000 391.200 58.800 391.800 ;
        RECT 78.000 391.200 81.600 391.800 ;
        RECT 100.800 391.200 101.400 391.800 ;
        RECT 52.800 390.600 58.200 391.200 ;
        RECT 76.200 390.600 81.600 391.200 ;
        RECT 100.200 390.600 101.400 391.200 ;
        RECT 103.200 391.200 106.800 391.800 ;
        RECT 132.000 391.200 135.000 392.400 ;
        RECT 214.800 391.800 222.000 392.400 ;
        RECT 213.600 391.200 220.200 391.800 ;
        RECT 226.800 391.200 229.200 392.400 ;
        RECT 484.200 391.200 487.200 392.400 ;
        RECT 520.200 391.800 527.400 392.400 ;
        RECT 543.600 391.800 551.400 392.400 ;
        RECT 625.200 391.800 631.200 392.400 ;
        RECT 519.600 391.200 525.600 391.800 ;
        RECT 545.400 391.200 552.000 391.800 ;
        RECT 626.400 391.200 631.800 391.800 ;
        RECT 103.200 390.600 107.400 391.200 ;
        RECT 132.600 390.600 135.600 391.200 ;
        RECT 213.000 390.600 219.000 391.200 ;
        RECT 226.200 390.600 228.600 391.200 ;
        RECT 52.200 390.000 57.600 390.600 ;
        RECT 75.000 390.000 81.600 390.600 ;
        RECT 99.000 390.000 101.400 390.600 ;
        RECT 103.800 390.000 108.600 390.600 ;
        RECT 133.200 390.000 135.600 390.600 ;
        RECT 211.800 390.000 217.800 390.600 ;
        RECT 225.600 390.000 228.600 390.600 ;
        RECT 483.600 390.000 486.600 391.200 ;
        RECT 518.400 390.600 524.400 391.200 ;
        RECT 547.200 390.600 553.200 391.200 ;
        RECT 627.600 390.600 633.000 391.200 ;
        RECT 517.800 390.000 523.200 390.600 ;
        RECT 548.400 390.000 554.400 390.600 ;
        RECT 628.200 390.000 634.200 390.600 ;
        RECT 51.600 389.400 57.600 390.000 ;
        RECT 73.800 389.400 81.600 390.000 ;
        RECT 98.400 389.400 101.400 390.000 ;
        RECT 104.400 389.400 109.800 390.000 ;
        RECT 134.400 389.400 135.000 390.000 ;
        RECT 211.200 389.400 216.600 390.000 ;
        RECT 225.600 389.400 228.000 390.000 ;
        RECT 483.000 389.400 486.600 390.000 ;
        RECT 517.200 389.400 522.000 390.000 ;
        RECT 549.600 389.400 555.000 390.000 ;
        RECT 629.400 389.400 634.800 390.000 ;
        RECT 50.400 388.800 57.600 389.400 ;
        RECT 72.600 388.800 81.000 389.400 ;
        RECT 97.800 388.800 102.600 389.400 ;
        RECT 104.400 388.800 113.400 389.400 ;
        RECT 118.800 388.800 126.000 389.400 ;
        RECT 210.600 388.800 215.400 389.400 ;
        RECT 225.000 388.800 228.000 389.400 ;
        RECT 49.800 388.200 57.600 388.800 ;
        RECT 71.400 388.200 77.400 388.800 ;
        RECT 49.200 387.600 57.600 388.200 ;
        RECT 70.200 387.600 76.800 388.200 ;
        RECT 48.000 387.000 52.800 387.600 ;
        RECT 47.400 386.400 52.200 387.000 ;
        RECT 46.200 385.800 51.600 386.400 ;
        RECT 45.600 385.200 50.400 385.800 ;
        RECT 54.600 385.200 57.600 387.600 ;
        RECT 69.000 387.000 75.600 387.600 ;
        RECT 78.600 387.000 81.000 388.800 ;
        RECT 97.200 388.200 126.000 388.800 ;
        RECT 210.000 388.200 214.800 388.800 ;
        RECT 225.000 388.200 227.400 388.800 ;
        RECT 96.600 387.600 124.800 388.200 ;
        RECT 209.400 387.600 214.200 388.200 ;
        RECT 224.400 387.600 227.400 388.200 ;
        RECT 482.400 388.200 486.000 389.400 ;
        RECT 516.600 388.800 521.400 389.400 ;
        RECT 550.800 388.800 556.200 389.400 ;
        RECT 630.000 388.800 636.000 389.400 ;
        RECT 516.000 388.200 520.200 388.800 ;
        RECT 551.400 388.200 556.800 388.800 ;
        RECT 631.200 388.200 636.600 388.800 ;
        RECT 482.400 387.600 485.400 388.200 ;
        RECT 515.400 387.600 519.600 388.200 ;
        RECT 552.600 387.600 557.400 388.200 ;
        RECT 632.400 387.600 637.800 388.200 ;
        RECT 96.000 387.000 123.600 387.600 ;
        RECT 208.800 387.000 213.600 387.600 ;
        RECT 223.800 387.000 226.800 387.600 ;
        RECT 67.800 386.400 74.400 387.000 ;
        RECT 66.600 385.800 73.200 386.400 ;
        RECT 64.800 385.200 72.000 385.800 ;
        RECT 45.000 384.600 49.800 385.200 ;
        RECT 54.600 384.600 58.200 385.200 ;
        RECT 63.000 384.600 70.800 385.200 ;
        RECT 78.600 384.600 81.600 387.000 ;
        RECT 94.800 386.400 99.600 387.000 ;
        RECT 100.800 386.400 121.800 387.000 ;
        RECT 208.200 386.400 213.000 387.000 ;
        RECT 223.200 386.400 226.800 387.000 ;
        RECT 481.800 387.000 485.400 387.600 ;
        RECT 514.800 387.000 519.000 387.600 ;
        RECT 553.200 387.000 558.000 387.600 ;
        RECT 633.000 387.000 639.000 387.600 ;
        RECT 481.800 386.400 484.800 387.000 ;
        RECT 514.200 386.400 518.400 387.000 ;
        RECT 554.400 386.400 558.600 387.000 ;
        RECT 634.200 386.400 639.600 387.000 ;
        RECT 94.200 385.800 99.000 386.400 ;
        RECT 102.000 385.800 109.200 386.400 ;
        RECT 114.000 385.800 121.200 386.400 ;
        RECT 207.600 385.800 212.400 386.400 ;
        RECT 223.200 385.800 226.200 386.400 ;
        RECT 93.600 385.200 98.400 385.800 ;
        RECT 105.000 385.200 106.800 385.800 ;
        RECT 92.400 384.600 97.200 385.200 ;
        RECT 43.800 384.000 49.200 384.600 ;
        RECT 54.600 384.000 69.600 384.600 ;
        RECT 79.200 384.000 82.200 384.600 ;
        RECT 91.200 384.000 96.600 384.600 ;
        RECT 105.000 384.000 106.200 385.200 ;
        RECT 117.600 384.600 121.200 385.800 ;
        RECT 207.000 385.200 211.800 385.800 ;
        RECT 222.600 385.200 225.600 385.800 ;
        RECT 481.200 385.200 484.800 386.400 ;
        RECT 513.600 385.800 517.800 386.400 ;
        RECT 555.000 385.800 559.200 386.400 ;
        RECT 635.400 385.800 640.800 386.400 ;
        RECT 513.000 385.200 517.200 385.800 ;
        RECT 555.600 385.200 559.800 385.800 ;
        RECT 636.000 385.200 641.400 385.800 ;
        RECT 206.400 384.600 211.200 385.200 ;
        RECT 222.000 384.600 225.000 385.200 ;
        RECT 481.200 384.600 484.200 385.200 ;
        RECT 513.000 384.600 516.600 385.200 ;
        RECT 556.200 384.600 560.400 385.200 ;
        RECT 637.200 384.600 642.600 385.200 ;
        RECT 117.000 384.000 120.600 384.600 ;
        RECT 205.800 384.000 210.600 384.600 ;
        RECT 221.400 384.000 225.000 384.600 ;
        RECT 43.200 383.400 48.000 384.000 ;
        RECT 55.200 383.400 68.400 384.000 ;
        RECT 79.200 383.400 82.800 384.000 ;
        RECT 90.000 383.400 96.000 384.000 ;
        RECT 105.000 383.400 106.800 384.000 ;
        RECT 116.400 383.400 120.000 384.000 ;
        RECT 205.200 383.400 210.000 384.000 ;
        RECT 220.800 383.400 224.400 384.000 ;
        RECT 42.000 382.800 47.400 383.400 ;
        RECT 55.800 382.800 66.600 383.400 ;
        RECT 79.800 382.800 83.400 383.400 ;
        RECT 88.800 382.800 94.800 383.400 ;
        RECT 41.400 382.200 46.200 382.800 ;
        RECT 56.400 382.200 64.800 382.800 ;
        RECT 79.800 382.200 94.200 382.800 ;
        RECT 105.000 382.200 107.400 383.400 ;
        RECT 115.800 382.800 120.000 383.400 ;
        RECT 204.600 382.800 208.800 383.400 ;
        RECT 219.600 382.800 223.800 383.400 ;
        RECT 480.600 382.800 484.200 384.600 ;
        RECT 512.400 384.000 516.000 384.600 ;
        RECT 556.800 384.000 561.000 384.600 ;
        RECT 637.800 384.000 643.200 384.600 ;
        RECT 511.800 383.400 515.400 384.000 ;
        RECT 558.000 383.400 561.600 384.000 ;
        RECT 639.000 383.400 644.400 384.000 ;
        RECT 511.800 382.800 514.800 383.400 ;
        RECT 558.000 382.800 562.200 383.400 ;
        RECT 639.600 382.800 645.000 383.400 ;
        RECT 115.200 382.200 119.400 382.800 ;
        RECT 163.800 382.200 166.200 382.800 ;
        RECT 203.400 382.200 208.200 382.800 ;
        RECT 219.000 382.200 223.200 382.800 ;
        RECT 40.800 381.600 45.600 382.200 ;
        RECT 57.000 381.600 63.000 382.200 ;
        RECT 67.800 381.600 71.400 382.200 ;
        RECT 80.400 381.600 93.000 382.200 ;
        RECT 39.600 381.000 45.000 381.600 ;
        RECT 66.000 381.000 71.400 381.600 ;
        RECT 81.000 381.000 91.800 381.600 ;
        RECT 39.000 380.400 43.800 381.000 ;
        RECT 64.200 380.400 71.400 381.000 ;
        RECT 81.600 380.400 90.600 381.000 ;
        RECT 105.000 380.400 108.000 382.200 ;
        RECT 114.600 381.600 118.800 382.200 ;
        RECT 163.200 381.600 167.400 382.200 ;
        RECT 202.800 381.600 207.600 382.200 ;
        RECT 218.400 381.600 222.600 382.200 ;
        RECT 114.000 381.000 118.200 381.600 ;
        RECT 163.200 381.000 169.200 381.600 ;
        RECT 202.200 381.000 207.000 381.600 ;
        RECT 217.800 381.000 222.000 381.600 ;
        RECT 480.000 381.000 483.600 382.800 ;
        RECT 511.200 382.200 514.800 382.800 ;
        RECT 558.600 382.200 562.800 382.800 ;
        RECT 640.800 382.200 646.200 382.800 ;
        RECT 510.600 381.600 514.200 382.200 ;
        RECT 559.200 381.600 563.400 382.200 ;
        RECT 641.400 381.600 646.800 382.200 ;
        RECT 510.600 381.000 513.600 381.600 ;
        RECT 559.800 381.000 563.400 381.600 ;
        RECT 642.600 381.000 648.000 381.600 ;
        RECT 112.800 380.400 117.600 381.000 ;
        RECT 163.800 380.400 171.000 381.000 ;
        RECT 201.000 380.400 206.400 381.000 ;
        RECT 217.200 380.400 221.400 381.000 ;
        RECT 480.000 380.400 483.000 381.000 ;
        RECT 38.400 379.800 43.200 380.400 ;
        RECT 63.600 379.800 71.400 380.400 ;
        RECT 82.800 379.800 88.800 380.400 ;
        RECT 37.200 379.200 42.000 379.800 ;
        RECT 63.000 379.200 70.200 379.800 ;
        RECT 104.400 379.200 107.400 380.400 ;
        RECT 112.200 379.800 117.000 380.400 ;
        RECT 164.400 379.800 172.800 380.400 ;
        RECT 199.800 379.800 205.800 380.400 ;
        RECT 216.000 379.800 220.800 380.400 ;
        RECT 111.000 379.200 116.400 379.800 ;
        RECT 165.600 379.200 174.600 379.800 ;
        RECT 198.600 379.200 204.600 379.800 ;
        RECT 215.400 379.200 220.200 379.800 ;
        RECT 36.600 378.600 41.400 379.200 ;
        RECT 63.000 378.600 67.800 379.200 ;
        RECT 91.800 378.600 93.000 379.200 ;
        RECT 103.800 378.600 107.400 379.200 ;
        RECT 110.400 378.600 115.200 379.200 ;
        RECT 133.200 378.600 133.800 379.200 ;
        RECT 167.400 378.600 177.000 379.200 ;
        RECT 196.800 378.600 204.000 379.200 ;
        RECT 214.800 378.600 219.000 379.200 ;
        RECT 479.400 378.600 483.000 380.400 ;
        RECT 510.000 380.400 513.600 381.000 ;
        RECT 560.400 380.400 564.000 381.000 ;
        RECT 643.200 380.400 648.600 381.000 ;
        RECT 510.000 379.200 513.000 380.400 ;
        RECT 561.000 379.200 564.600 380.400 ;
        RECT 644.400 379.800 649.200 380.400 ;
        RECT 645.000 379.200 650.400 379.800 ;
        RECT 35.400 378.000 40.800 378.600 ;
        RECT 34.800 377.400 39.600 378.000 ;
        RECT 34.200 376.800 39.000 377.400 ;
        RECT 33.000 376.200 38.400 376.800 ;
        RECT 63.000 376.200 66.000 378.600 ;
        RECT 91.200 378.000 93.600 378.600 ;
        RECT 103.200 378.000 106.800 378.600 ;
        RECT 91.200 376.800 94.200 378.000 ;
        RECT 102.600 377.400 106.800 378.000 ;
        RECT 109.800 377.400 114.600 378.600 ;
        RECT 130.800 378.000 134.400 378.600 ;
        RECT 168.600 378.000 179.400 378.600 ;
        RECT 194.400 378.000 202.800 378.600 ;
        RECT 213.600 378.000 218.400 378.600 ;
        RECT 479.400 378.000 482.400 378.600 ;
        RECT 129.000 377.400 133.800 378.000 ;
        RECT 170.400 377.400 181.800 378.000 ;
        RECT 191.400 377.400 201.600 378.000 ;
        RECT 213.000 377.400 217.200 378.000 ;
        RECT 102.000 376.800 106.200 377.400 ;
        RECT 109.800 376.800 116.400 377.400 ;
        RECT 126.600 376.800 133.200 377.400 ;
        RECT 172.200 376.800 200.400 377.400 ;
        RECT 211.800 376.800 216.600 377.400 ;
        RECT 79.800 376.200 81.600 376.800 ;
        RECT 90.000 376.200 94.800 376.800 ;
        RECT 101.400 376.200 105.600 376.800 ;
        RECT 110.400 376.200 121.200 376.800 ;
        RECT 122.400 376.200 132.600 376.800 ;
        RECT 174.000 376.200 198.600 376.800 ;
        RECT 211.200 376.200 216.000 376.800 ;
        RECT 478.800 376.200 482.400 378.000 ;
        RECT 509.400 377.400 512.400 379.200 ;
        RECT 561.600 378.600 565.200 379.200 ;
        RECT 646.200 378.600 651.000 379.200 ;
        RECT 562.200 378.000 565.800 378.600 ;
        RECT 646.800 378.000 651.600 378.600 ;
        RECT 562.800 377.400 565.800 378.000 ;
        RECT 647.400 377.400 652.800 378.000 ;
        RECT 32.400 375.600 37.200 376.200 ;
        RECT 63.000 375.600 66.600 376.200 ;
        RECT 78.600 375.600 82.800 376.200 ;
        RECT 88.200 375.600 94.800 376.200 ;
        RECT 100.200 375.600 105.000 376.200 ;
        RECT 111.000 375.600 131.400 376.200 ;
        RECT 176.400 375.600 196.800 376.200 ;
        RECT 210.000 375.600 214.800 376.200 ;
        RECT 31.200 375.000 36.600 375.600 ;
        RECT 63.600 375.000 66.600 375.600 ;
        RECT 76.800 375.000 84.600 375.600 ;
        RECT 86.400 375.000 95.400 375.600 ;
        RECT 99.000 375.000 104.400 375.600 ;
        RECT 112.200 375.000 130.200 375.600 ;
        RECT 178.800 375.000 195.000 375.600 ;
        RECT 208.800 375.000 214.200 375.600 ;
        RECT 478.800 375.000 481.800 376.200 ;
        RECT 508.800 375.000 511.800 377.400 ;
        RECT 562.800 376.800 566.400 377.400 ;
        RECT 648.600 376.800 653.400 377.400 ;
        RECT 563.400 376.200 566.400 376.800 ;
        RECT 649.200 376.200 654.000 376.800 ;
        RECT 563.400 375.600 567.000 376.200 ;
        RECT 649.800 375.600 654.600 376.200 ;
        RECT 564.000 375.000 567.000 375.600 ;
        RECT 651.000 375.000 655.800 375.600 ;
        RECT 30.600 374.400 35.400 375.000 ;
        RECT 63.600 374.400 67.200 375.000 ;
        RECT 75.600 374.400 91.200 375.000 ;
        RECT 92.400 374.400 96.000 375.000 ;
        RECT 97.800 374.400 103.800 375.000 ;
        RECT 114.000 374.400 129.000 375.000 ;
        RECT 182.400 374.400 191.400 375.000 ;
        RECT 207.000 374.400 213.000 375.000 ;
        RECT 29.400 373.800 34.800 374.400 ;
        RECT 64.200 373.800 67.800 374.400 ;
        RECT 73.800 373.800 90.600 374.400 ;
        RECT 92.400 373.800 102.600 374.400 ;
        RECT 116.400 373.800 129.000 374.400 ;
        RECT 205.200 373.800 211.800 374.400 ;
        RECT 28.800 373.200 34.200 373.800 ;
        RECT 64.200 373.200 90.000 373.800 ;
        RECT 93.000 373.200 102.000 373.800 ;
        RECT 28.200 372.600 33.000 373.200 ;
        RECT 64.800 372.600 78.600 373.200 ;
        RECT 82.200 372.600 88.800 373.200 ;
        RECT 93.600 372.600 100.800 373.200 ;
        RECT 27.000 372.000 32.400 372.600 ;
        RECT 65.400 372.000 77.400 372.600 ;
        RECT 84.600 372.000 86.400 372.600 ;
        RECT 94.200 372.000 99.600 372.600 ;
        RECT 124.800 372.000 128.400 373.800 ;
        RECT 202.800 373.200 210.600 373.800 ;
        RECT 478.200 373.200 481.800 375.000 ;
        RECT 147.000 372.600 148.800 373.200 ;
        RECT 159.000 372.600 169.800 373.200 ;
        RECT 199.200 372.600 208.800 373.200 ;
        RECT 142.800 372.000 150.000 372.600 ;
        RECT 159.000 372.000 176.400 372.600 ;
        RECT 193.200 372.000 207.000 372.600 ;
        RECT 478.200 372.000 481.200 373.200 ;
        RECT 26.400 371.400 31.200 372.000 ;
        RECT 66.600 371.400 76.200 372.000 ;
        RECT 95.400 371.400 97.800 372.000 ;
        RECT 123.600 371.400 127.800 372.000 ;
        RECT 140.400 371.400 149.400 372.000 ;
        RECT 159.600 371.400 205.200 372.000 ;
        RECT 25.200 370.800 30.600 371.400 ;
        RECT 67.800 370.800 73.800 371.400 ;
        RECT 123.000 370.800 127.800 371.400 ;
        RECT 138.600 370.800 147.600 371.400 ;
        RECT 161.400 370.800 202.800 371.400 ;
        RECT 24.600 370.200 29.400 370.800 ;
        RECT 121.800 370.200 127.200 370.800 ;
        RECT 136.200 370.200 146.400 370.800 ;
        RECT 164.400 370.200 200.400 370.800 ;
        RECT 23.400 369.600 28.800 370.200 ;
        RECT 120.600 369.600 126.600 370.200 ;
        RECT 134.400 369.600 144.600 370.200 ;
        RECT 169.800 369.600 195.600 370.200 ;
        RECT 222.600 369.600 227.400 370.200 ;
        RECT 22.800 369.000 27.600 369.600 ;
        RECT 118.800 369.000 126.600 369.600 ;
        RECT 132.000 369.000 143.400 369.600 ;
        RECT 177.000 369.000 179.400 369.600 ;
        RECT 184.800 369.000 188.400 369.600 ;
        RECT 218.400 369.000 231.600 369.600 ;
        RECT 477.600 369.000 481.200 372.000 ;
        RECT 21.600 368.400 27.000 369.000 ;
        RECT 117.600 368.400 126.600 369.000 ;
        RECT 129.000 368.400 143.400 369.000 ;
        RECT 21.000 367.800 27.000 368.400 ;
        RECT 116.400 367.800 138.600 368.400 ;
        RECT 19.800 367.200 42.600 367.800 ;
        RECT 115.200 367.200 122.400 367.800 ;
        RECT 123.600 367.200 136.200 367.800 ;
        RECT 141.000 367.200 144.000 368.400 ;
        RECT 185.400 367.800 188.400 369.000 ;
        RECT 216.000 368.400 234.000 369.000 ;
        RECT 214.200 367.800 235.800 368.400 ;
        RECT 261.000 367.800 264.000 368.400 ;
        RECT 185.400 367.200 189.000 367.800 ;
        RECT 212.400 367.200 237.000 367.800 ;
        RECT 260.400 367.200 264.600 367.800 ;
        RECT 477.600 367.200 480.600 369.000 ;
        RECT 18.600 366.600 51.000 367.200 ;
        RECT 114.000 366.600 121.200 367.200 ;
        RECT 123.600 366.600 134.400 367.200 ;
        RECT 141.600 366.600 144.600 367.200 ;
        RECT 186.000 366.600 189.000 367.200 ;
        RECT 211.200 366.600 222.000 367.200 ;
        RECT 228.000 366.600 238.200 367.200 ;
        RECT 259.800 366.600 265.200 367.200 ;
        RECT 18.000 366.000 56.400 366.600 ;
        RECT 112.200 366.000 120.000 366.600 ;
        RECT 124.200 366.000 132.000 366.600 ;
        RECT 141.600 366.000 145.200 366.600 ;
        RECT 186.000 366.000 189.600 366.600 ;
        RECT 210.000 366.000 218.400 366.600 ;
        RECT 231.600 366.000 239.400 366.600 ;
        RECT 259.800 366.000 265.800 366.600 ;
        RECT 17.400 365.400 60.000 366.000 ;
        RECT 111.000 365.400 118.800 366.000 ;
        RECT 125.400 365.400 129.000 366.000 ;
        RECT 142.200 365.400 145.200 366.000 ;
        RECT 186.600 365.400 189.600 366.000 ;
        RECT 208.800 365.400 216.000 366.000 ;
        RECT 233.400 365.400 240.600 366.000 ;
        RECT 259.800 365.400 266.400 366.000 ;
        RECT 17.400 364.800 63.600 365.400 ;
        RECT 109.200 364.800 117.600 365.400 ;
        RECT 142.200 364.800 145.800 365.400 ;
        RECT 186.600 364.800 190.200 365.400 ;
        RECT 207.600 364.800 214.200 365.400 ;
        RECT 235.200 364.800 241.200 365.400 ;
        RECT 259.200 364.800 266.400 365.400 ;
        RECT 43.800 364.200 66.600 364.800 ;
        RECT 108.000 364.200 115.800 364.800 ;
        RECT 51.600 363.600 69.600 364.200 ;
        RECT 106.200 363.600 114.600 364.200 ;
        RECT 142.800 363.600 145.800 364.800 ;
        RECT 187.200 364.200 190.800 364.800 ;
        RECT 206.400 364.200 213.000 364.800 ;
        RECT 236.400 364.200 242.400 364.800 ;
        RECT 187.200 363.600 192.000 364.200 ;
        RECT 205.200 363.600 211.800 364.200 ;
        RECT 237.600 363.600 243.000 364.200 ;
        RECT 56.400 363.000 73.200 363.600 ;
        RECT 103.800 363.000 113.400 363.600 ;
        RECT 60.600 362.400 76.200 363.000 ;
        RECT 102.000 362.400 112.200 363.000 ;
        RECT 143.400 362.400 146.400 363.600 ;
        RECT 187.800 363.000 192.600 363.600 ;
        RECT 204.000 363.000 210.600 363.600 ;
        RECT 238.800 363.000 243.600 363.600 ;
        RECT 188.400 362.400 193.800 363.000 ;
        RECT 202.800 362.400 209.400 363.000 ;
        RECT 239.400 362.400 244.200 363.000 ;
        RECT 259.200 362.400 262.200 364.800 ;
        RECT 263.400 364.200 267.000 364.800 ;
        RECT 264.000 363.600 267.600 364.200 ;
        RECT 264.600 363.000 267.600 363.600 ;
        RECT 477.000 363.600 480.600 367.200 ;
        RECT 508.200 367.200 511.200 375.000 ;
        RECT 564.000 374.400 567.600 375.000 ;
        RECT 651.600 374.400 656.400 375.000 ;
        RECT 564.600 373.800 567.600 374.400 ;
        RECT 652.200 373.800 657.000 374.400 ;
        RECT 564.600 373.200 568.200 373.800 ;
        RECT 652.800 373.200 657.600 373.800 ;
        RECT 565.200 372.600 568.200 373.200 ;
        RECT 654.000 372.600 658.200 373.200 ;
        RECT 565.200 372.000 568.800 372.600 ;
        RECT 654.600 372.000 658.800 372.600 ;
        RECT 565.800 371.400 568.800 372.000 ;
        RECT 655.200 371.400 660.000 372.000 ;
        RECT 565.800 370.800 569.400 371.400 ;
        RECT 655.800 370.800 660.600 371.400 ;
        RECT 566.400 369.600 569.400 370.800 ;
        RECT 656.400 370.200 661.200 370.800 ;
        RECT 657.600 369.600 661.800 370.200 ;
        RECT 566.400 369.000 570.000 369.600 ;
        RECT 658.200 369.000 662.400 369.600 ;
        RECT 567.000 367.800 570.000 369.000 ;
        RECT 658.800 368.400 663.000 369.000 ;
        RECT 659.400 367.800 663.600 368.400 ;
        RECT 508.200 366.000 510.600 367.200 ;
        RECT 567.600 366.000 570.600 367.800 ;
        RECT 660.000 367.200 664.200 367.800 ;
        RECT 660.600 366.600 664.800 367.200 ;
        RECT 661.200 366.000 665.400 366.600 ;
        RECT 264.600 362.400 268.200 363.000 ;
        RECT 63.600 361.800 79.200 362.400 ;
        RECT 99.600 361.800 110.400 362.400 ;
        RECT 143.400 361.800 147.000 362.400 ;
        RECT 189.000 361.800 195.600 362.400 ;
        RECT 201.600 361.800 208.200 362.400 ;
        RECT 240.600 361.800 244.800 362.400 ;
        RECT 259.200 361.800 261.600 362.400 ;
        RECT 67.200 361.200 84.000 361.800 ;
        RECT 95.400 361.200 108.600 361.800 ;
        RECT 70.200 360.600 107.400 361.200 ;
        RECT 73.200 360.000 105.000 360.600 ;
        RECT 144.000 360.000 147.000 361.800 ;
        RECT 190.200 361.200 207.000 361.800 ;
        RECT 241.200 361.200 245.400 361.800 ;
        RECT 190.800 360.600 206.400 361.200 ;
        RECT 241.800 360.600 246.000 361.200 ;
        RECT 191.400 360.000 205.200 360.600 ;
        RECT 242.400 360.000 246.600 360.600 ;
        RECT 76.200 359.400 103.200 360.000 ;
        RECT 79.800 358.800 99.600 359.400 ;
        RECT 84.000 358.200 94.800 358.800 ;
        RECT 144.600 357.600 147.600 360.000 ;
        RECT 192.600 359.400 204.000 360.000 ;
        RECT 243.000 359.400 246.600 360.000 ;
        RECT 145.200 357.000 147.600 357.600 ;
        RECT 195.600 358.800 202.800 359.400 ;
        RECT 243.600 358.800 247.200 359.400 ;
        RECT 195.600 358.200 201.600 358.800 ;
        RECT 244.200 358.200 247.800 358.800 ;
        RECT 195.600 357.600 200.400 358.200 ;
        RECT 211.200 357.600 212.400 358.200 ;
        RECT 195.600 357.000 199.200 357.600 ;
        RECT 210.000 357.000 213.600 357.600 ;
        RECT 244.800 357.000 248.400 358.200 ;
        RECT 145.200 354.600 148.200 357.000 ;
        RECT 196.200 356.400 198.000 357.000 ;
        RECT 209.400 356.400 214.800 357.000 ;
        RECT 245.400 356.400 249.000 357.000 ;
        RECT 208.800 355.800 215.400 356.400 ;
        RECT 246.000 355.800 249.000 356.400 ;
        RECT 258.600 356.400 261.600 361.800 ;
        RECT 265.200 361.800 268.200 362.400 ;
        RECT 265.200 361.200 268.800 361.800 ;
        RECT 265.800 360.600 268.800 361.200 ;
        RECT 265.800 360.000 269.400 360.600 ;
        RECT 477.000 360.000 480.000 363.600 ;
        RECT 508.200 361.800 511.200 366.000 ;
        RECT 568.200 364.200 571.200 366.000 ;
        RECT 661.800 365.400 666.000 366.000 ;
        RECT 662.400 364.800 666.600 365.400 ;
        RECT 663.000 364.200 667.200 364.800 ;
        RECT 568.800 362.400 571.800 364.200 ;
        RECT 663.600 363.600 667.800 364.200 ;
        RECT 664.200 363.000 668.400 363.600 ;
        RECT 664.800 362.400 669.000 363.000 ;
        RECT 266.400 358.800 269.400 360.000 ;
        RECT 267.000 357.600 270.000 358.800 ;
        RECT 267.000 357.000 270.600 357.600 ;
        RECT 258.600 355.800 261.000 356.400 ;
        RECT 208.200 355.200 216.000 355.800 ;
        RECT 246.000 355.200 249.600 355.800 ;
        RECT 207.600 354.600 216.600 355.200 ;
        RECT 246.600 354.600 249.600 355.200 ;
        RECT 145.200 353.400 147.600 354.600 ;
        RECT 207.000 354.000 210.600 354.600 ;
        RECT 213.000 354.000 217.200 354.600 ;
        RECT 246.600 354.000 250.200 354.600 ;
        RECT 206.400 353.400 210.600 354.000 ;
        RECT 213.600 353.400 217.800 354.000 ;
        RECT 144.600 350.400 147.600 353.400 ;
        RECT 205.800 352.800 210.000 353.400 ;
        RECT 214.200 352.800 217.800 353.400 ;
        RECT 247.200 353.400 250.200 354.000 ;
        RECT 247.200 352.800 250.800 353.400 ;
        RECT 205.800 352.200 209.400 352.800 ;
        RECT 214.800 352.200 218.400 352.800 ;
        RECT 205.200 351.600 208.800 352.200 ;
        RECT 215.400 351.600 218.400 352.200 ;
        RECT 247.800 352.200 250.800 352.800 ;
        RECT 247.800 351.600 251.400 352.200 ;
        RECT 204.600 351.000 208.200 351.600 ;
        RECT 215.400 351.000 219.000 351.600 ;
        RECT 144.000 348.600 147.000 350.400 ;
        RECT 204.000 349.800 207.600 351.000 ;
        RECT 216.000 350.400 219.000 351.000 ;
        RECT 248.400 351.000 251.400 351.600 ;
        RECT 248.400 350.400 252.000 351.000 ;
        RECT 216.000 349.800 219.600 350.400 ;
        RECT 203.400 349.200 207.000 349.800 ;
        RECT 143.400 348.000 149.400 348.600 ;
        RECT 193.800 348.000 195.000 348.600 ;
        RECT 202.800 348.000 206.400 349.200 ;
        RECT 216.600 348.600 219.600 349.800 ;
        RECT 249.000 349.200 252.000 350.400 ;
        RECT 249.000 348.600 252.600 349.200 ;
        RECT 143.400 347.400 150.600 348.000 ;
        RECT 192.600 347.400 196.800 348.000 ;
        RECT 202.200 347.400 205.800 348.000 ;
        RECT 142.200 346.800 150.000 347.400 ;
        RECT 192.000 346.800 198.000 347.400 ;
        RECT 202.200 346.800 205.200 347.400 ;
        RECT 141.000 346.200 149.400 346.800 ;
        RECT 192.000 346.200 199.200 346.800 ;
        RECT 201.600 346.200 205.200 346.800 ;
        RECT 217.200 346.800 220.200 348.600 ;
        RECT 249.600 347.400 252.600 348.600 ;
        RECT 258.000 348.000 261.000 355.800 ;
        RECT 267.600 355.800 270.600 357.000 ;
        RECT 476.400 357.000 480.000 360.000 ;
        RECT 508.800 360.600 511.200 361.800 ;
        RECT 267.600 355.200 271.200 355.800 ;
        RECT 268.200 354.000 271.200 355.200 ;
        RECT 268.800 352.200 271.800 354.000 ;
        RECT 268.800 351.600 272.400 352.200 ;
        RECT 269.400 349.800 272.400 351.600 ;
        RECT 222.000 346.800 229.200 347.400 ;
        RECT 217.200 346.200 235.200 346.800 ;
        RECT 140.400 345.600 148.200 346.200 ;
        RECT 191.400 345.600 199.800 346.200 ;
        RECT 201.000 345.600 204.600 346.200 ;
        RECT 217.200 345.600 238.800 346.200 ;
        RECT 139.200 345.000 146.400 345.600 ;
        RECT 191.400 345.000 204.000 345.600 ;
        RECT 138.000 344.400 145.200 345.000 ;
        RECT 191.400 344.400 194.400 345.000 ;
        RECT 196.200 344.400 204.000 345.000 ;
        RECT 217.200 345.000 241.200 345.600 ;
        RECT 250.200 345.000 253.200 347.400 ;
        RECT 258.000 346.800 260.400 348.000 ;
        RECT 270.000 347.400 273.000 349.800 ;
        RECT 217.200 344.400 243.600 345.000 ;
        RECT 137.400 343.800 143.400 344.400 ;
        RECT 136.200 343.200 142.200 343.800 ;
        RECT 135.000 342.600 141.000 343.200 ;
        RECT 190.800 342.600 193.800 344.400 ;
        RECT 197.400 343.800 203.400 344.400 ;
        RECT 198.600 343.200 203.400 343.800 ;
        RECT 217.200 343.200 220.200 344.400 ;
        RECT 230.400 343.800 245.400 344.400 ;
        RECT 235.800 343.200 247.200 343.800 ;
        RECT 133.800 342.000 140.400 342.600 ;
        RECT 132.600 341.400 139.200 342.000 ;
        RECT 131.400 340.800 138.000 341.400 ;
        RECT 190.200 340.800 193.200 342.600 ;
        RECT 199.200 342.000 203.400 343.200 ;
        RECT 199.800 341.400 203.400 342.000 ;
        RECT 216.600 341.400 219.600 343.200 ;
        RECT 238.800 342.600 248.400 343.200 ;
        RECT 250.800 342.600 253.800 345.000 ;
        RECT 241.200 342.000 249.600 342.600 ;
        RECT 250.800 342.000 254.400 342.600 ;
        RECT 222.600 341.400 224.400 342.000 ;
        RECT 243.600 341.400 254.400 342.000 ;
        RECT 200.400 340.800 203.400 341.400 ;
        RECT 216.000 340.800 219.600 341.400 ;
        RECT 220.800 340.800 225.600 341.400 ;
        RECT 244.800 340.800 254.400 341.400 ;
        RECT 130.200 340.200 136.800 340.800 ;
        RECT 129.600 339.600 135.600 340.200 ;
        RECT 128.400 339.000 134.400 339.600 ;
        RECT 163.200 339.000 171.000 339.600 ;
        RECT 189.600 339.000 192.600 340.800 ;
        RECT 127.200 338.400 133.200 339.000 ;
        RECT 159.000 338.400 170.400 339.000 ;
        RECT 189.000 338.400 192.600 339.000 ;
        RECT 126.600 337.800 132.000 338.400 ;
        RECT 154.800 337.800 169.200 338.400 ;
        RECT 125.400 337.200 131.400 337.800 ;
        RECT 150.600 337.200 167.400 337.800 ;
        RECT 189.000 337.200 192.000 338.400 ;
        RECT 201.000 337.200 204.000 340.800 ;
        RECT 216.000 340.200 226.200 340.800 ;
        RECT 246.600 340.200 254.400 340.800 ;
        RECT 215.400 339.600 226.800 340.200 ;
        RECT 247.800 339.600 255.000 340.200 ;
        RECT 257.400 339.600 260.400 346.800 ;
        RECT 270.600 345.000 273.600 347.400 ;
        RECT 281.400 345.000 284.400 345.600 ;
        RECT 271.200 342.600 274.200 345.000 ;
        RECT 281.400 344.400 285.000 345.000 ;
        RECT 280.800 343.800 285.600 344.400 ;
        RECT 476.400 343.800 479.400 357.000 ;
        RECT 508.800 356.400 511.800 360.600 ;
        RECT 569.400 360.000 572.400 362.400 ;
        RECT 665.400 361.800 669.600 362.400 ;
        RECT 666.000 361.200 670.200 361.800 ;
        RECT 666.600 360.600 670.800 361.200 ;
        RECT 667.200 360.000 671.400 360.600 ;
        RECT 570.000 357.600 573.000 360.000 ;
        RECT 667.800 359.400 672.000 360.000 ;
        RECT 668.400 358.800 672.000 359.400 ;
        RECT 669.000 358.200 672.600 358.800 ;
        RECT 669.600 357.600 673.200 358.200 ;
        RECT 509.400 352.800 512.400 356.400 ;
        RECT 570.600 355.800 573.600 357.600 ;
        RECT 670.200 357.000 673.800 357.600 ;
        RECT 670.200 356.400 674.400 357.000 ;
        RECT 670.800 355.800 675.000 356.400 ;
        RECT 571.200 353.400 574.200 355.800 ;
        RECT 671.400 355.200 675.600 355.800 ;
        RECT 672.000 354.600 675.600 355.200 ;
        RECT 672.600 354.000 676.200 354.600 ;
        RECT 673.200 353.400 676.800 354.000 ;
        RECT 510.000 349.800 513.000 352.800 ;
        RECT 571.800 351.600 574.800 353.400 ;
        RECT 673.800 352.800 677.400 353.400 ;
        RECT 673.800 352.200 678.000 352.800 ;
        RECT 674.400 351.600 678.000 352.200 ;
        RECT 571.800 351.000 575.400 351.600 ;
        RECT 675.000 351.000 678.600 351.600 ;
        RECT 510.600 347.400 513.600 349.800 ;
        RECT 572.400 349.200 575.400 351.000 ;
        RECT 675.600 350.400 679.200 351.000 ;
        RECT 676.200 349.800 679.800 350.400 ;
        RECT 676.200 349.200 680.400 349.800 ;
        RECT 511.200 345.600 514.200 347.400 ;
        RECT 573.000 346.800 576.000 349.200 ;
        RECT 676.800 348.600 680.400 349.200 ;
        RECT 677.400 348.000 681.000 348.600 ;
        RECT 678.000 347.400 681.600 348.000 ;
        RECT 678.000 346.800 682.200 347.400 ;
        RECT 511.800 344.400 514.800 345.600 ;
        RECT 573.600 345.000 576.600 346.800 ;
        RECT 678.600 346.200 682.200 346.800 ;
        RECT 679.200 345.600 682.800 346.200 ;
        RECT 573.600 344.400 577.200 345.000 ;
        RECT 679.800 344.400 683.400 345.600 ;
        RECT 280.200 342.600 286.200 343.800 ;
        RECT 477.000 343.200 479.400 343.800 ;
        RECT 512.400 343.800 514.800 344.400 ;
        RECT 271.800 339.600 274.800 342.600 ;
        RECT 279.600 342.000 286.800 342.600 ;
        RECT 279.600 341.400 282.600 342.000 ;
        RECT 279.000 340.800 282.600 341.400 ;
        RECT 283.800 341.400 286.800 342.000 ;
        RECT 283.800 340.800 287.400 341.400 ;
        RECT 279.000 340.200 282.000 340.800 ;
        RECT 278.400 339.600 282.000 340.200 ;
        RECT 284.400 339.600 287.400 340.800 ;
        RECT 214.800 339.000 226.800 339.600 ;
        RECT 249.600 339.000 255.000 339.600 ;
        RECT 256.800 339.000 260.400 339.600 ;
        RECT 214.800 338.400 222.600 339.000 ;
        RECT 213.600 337.800 220.800 338.400 ;
        RECT 213.000 337.200 219.600 337.800 ;
        RECT 124.800 336.600 130.200 337.200 ;
        RECT 148.200 336.600 165.000 337.200 ;
        RECT 189.000 336.600 191.400 337.200 ;
        RECT 201.000 336.600 203.400 337.200 ;
        RECT 212.400 336.600 218.400 337.200 ;
        RECT 123.600 336.000 129.000 336.600 ;
        RECT 146.400 336.000 162.000 336.600 ;
        RECT 189.600 336.000 190.800 336.600 ;
        RECT 212.400 336.000 217.200 336.600 ;
        RECT 223.800 336.000 226.800 339.000 ;
        RECT 250.200 338.400 259.800 339.000 ;
        RECT 251.400 337.800 259.800 338.400 ;
        RECT 252.600 337.200 259.800 337.800 ;
        RECT 272.400 337.200 275.400 339.600 ;
        RECT 278.400 339.000 281.400 339.600 ;
        RECT 277.800 338.400 281.400 339.000 ;
        RECT 277.800 337.200 280.800 338.400 ;
        RECT 285.000 337.800 288.000 339.600 ;
        RECT 477.000 339.000 480.000 343.200 ;
        RECT 512.400 342.600 515.400 343.800 ;
        RECT 574.200 342.600 577.200 344.400 ;
        RECT 680.400 343.800 684.000 344.400 ;
        RECT 680.400 343.200 684.600 343.800 ;
        RECT 681.000 342.600 684.600 343.200 ;
        RECT 513.000 342.000 515.400 342.600 ;
        RECT 513.000 340.800 516.000 342.000 ;
        RECT 574.800 340.800 577.800 342.600 ;
        RECT 681.600 342.000 685.200 342.600 ;
        RECT 681.600 341.400 685.800 342.000 ;
        RECT 682.200 340.800 685.800 341.400 ;
        RECT 513.600 339.000 516.600 340.800 ;
        RECT 574.800 340.200 578.400 340.800 ;
        RECT 477.600 338.400 480.000 339.000 ;
        RECT 253.200 336.600 259.800 337.200 ;
        RECT 254.400 336.000 259.800 336.600 ;
        RECT 123.000 335.400 128.400 336.000 ;
        RECT 147.000 335.400 158.400 336.000 ;
        RECT 212.400 335.400 216.000 336.000 ;
        RECT 223.200 335.400 226.800 336.000 ;
        RECT 255.000 335.400 259.800 336.000 ;
        RECT 273.000 336.000 276.000 337.200 ;
        RECT 277.200 336.600 280.800 337.200 ;
        RECT 277.200 336.000 280.200 336.600 ;
        RECT 273.000 335.400 280.200 336.000 ;
        RECT 285.600 336.000 288.600 337.800 ;
        RECT 285.600 335.400 289.200 336.000 ;
        RECT 477.600 335.400 480.600 338.400 ;
        RECT 514.200 337.200 517.200 339.000 ;
        RECT 575.400 338.400 578.400 340.200 ;
        RECT 682.800 339.600 686.400 340.800 ;
        RECT 683.400 339.000 687.000 339.600 ;
        RECT 514.800 336.000 517.800 337.200 ;
        RECT 576.000 336.600 579.000 338.400 ;
        RECT 684.000 337.800 687.600 339.000 ;
        RECT 684.600 336.600 688.200 337.800 ;
        RECT 514.800 335.400 518.400 336.000 ;
        RECT 122.400 334.800 127.200 335.400 ;
        RECT 223.200 334.800 226.200 335.400 ;
        RECT 256.200 334.800 260.400 335.400 ;
        RECT 121.800 334.200 126.600 334.800 ;
        RECT 222.600 334.200 226.200 334.800 ;
        RECT 256.800 334.200 261.000 334.800 ;
        RECT 273.000 334.200 279.600 335.400 ;
        RECT 120.600 333.600 125.400 334.200 ;
        RECT 222.000 333.600 225.600 334.200 ;
        RECT 257.400 333.600 261.600 334.200 ;
        RECT 120.000 333.000 124.800 333.600 ;
        RECT 220.800 333.000 225.600 333.600 ;
        RECT 258.000 333.000 262.200 333.600 ;
        RECT 119.400 332.400 124.200 333.000 ;
        RECT 219.000 332.400 225.600 333.000 ;
        RECT 259.200 332.400 262.800 333.000 ;
        RECT 273.600 332.400 279.000 334.200 ;
        RECT 286.200 333.000 289.200 335.400 ;
        RECT 118.800 331.800 123.000 332.400 ;
        RECT 193.800 331.800 208.800 332.400 ;
        RECT 218.400 331.800 227.400 332.400 ;
        RECT 259.800 331.800 263.400 332.400 ;
        RECT 273.600 331.800 278.400 332.400 ;
        RECT 118.200 331.200 122.400 331.800 ;
        RECT 189.600 331.200 212.400 331.800 ;
        RECT 218.400 331.200 228.600 331.800 ;
        RECT 260.400 331.200 264.000 331.800 ;
        RECT 117.600 330.600 121.800 331.200 ;
        RECT 186.600 330.600 214.800 331.200 ;
        RECT 218.400 330.600 229.800 331.200 ;
        RECT 261.000 330.600 264.600 331.200 ;
        RECT 274.200 330.600 278.400 331.800 ;
        RECT 286.800 330.600 289.800 333.000 ;
        RECT 478.200 332.400 481.200 335.400 ;
        RECT 515.400 334.200 518.400 335.400 ;
        RECT 576.600 334.800 579.600 336.600 ;
        RECT 685.200 336.000 688.800 336.600 ;
        RECT 685.800 335.400 688.800 336.000 ;
        RECT 685.800 334.800 689.400 335.400 ;
        RECT 576.600 334.200 580.200 334.800 ;
        RECT 516.000 333.000 519.000 334.200 ;
        RECT 577.200 333.000 580.200 334.200 ;
        RECT 686.400 334.200 689.400 334.800 ;
        RECT 686.400 333.600 690.000 334.200 ;
        RECT 687.000 333.000 690.000 333.600 ;
        RECT 516.000 332.400 519.600 333.000 ;
        RECT 577.200 332.400 580.800 333.000 ;
        RECT 687.000 332.400 690.600 333.000 ;
        RECT 478.200 331.800 481.800 332.400 ;
        RECT 117.000 330.000 121.200 330.600 ;
        RECT 184.200 330.000 216.600 330.600 ;
        RECT 218.400 330.000 230.400 330.600 ;
        RECT 261.000 330.000 265.200 330.600 ;
        RECT 116.400 329.400 120.600 330.000 ;
        RECT 181.800 329.400 199.800 330.000 ;
        RECT 202.800 329.400 220.200 330.000 ;
        RECT 225.600 329.400 231.000 330.000 ;
        RECT 261.600 329.400 265.800 330.000 ;
        RECT 115.800 328.800 120.000 329.400 ;
        RECT 180.000 328.800 193.200 329.400 ;
        RECT 208.800 328.800 220.200 329.400 ;
        RECT 226.800 328.800 231.600 329.400 ;
        RECT 262.200 328.800 265.800 329.400 ;
        RECT 274.200 328.800 277.800 330.600 ;
        RECT 287.400 330.000 289.800 330.600 ;
        RECT 478.800 330.000 481.800 331.800 ;
        RECT 516.600 331.200 519.600 332.400 ;
        RECT 577.800 331.200 580.800 332.400 ;
        RECT 687.600 331.800 691.200 332.400 ;
        RECT 688.200 331.200 691.200 331.800 ;
        RECT 517.200 330.000 520.200 331.200 ;
        RECT 577.800 330.600 581.400 331.200 ;
        RECT 115.800 328.200 119.400 328.800 ;
        RECT 178.200 328.200 189.600 328.800 ;
        RECT 212.400 328.200 221.400 328.800 ;
        RECT 115.200 327.600 118.800 328.200 ;
        RECT 177.600 327.600 186.600 328.200 ;
        RECT 214.200 327.600 223.200 328.200 ;
        RECT 114.600 327.000 118.200 327.600 ;
        RECT 177.000 327.000 183.600 327.600 ;
        RECT 216.600 327.000 224.400 327.600 ;
        RECT 228.000 327.000 231.600 328.800 ;
        RECT 262.800 328.200 266.400 328.800 ;
        RECT 263.400 327.600 267.000 328.200 ;
        RECT 114.000 326.400 117.600 327.000 ;
        RECT 178.200 326.400 180.600 327.000 ;
        RECT 218.400 326.400 225.600 327.000 ;
        RECT 226.800 326.400 231.600 327.000 ;
        RECT 264.000 326.400 267.600 327.600 ;
        RECT 274.200 327.000 277.200 328.800 ;
        RECT 273.600 326.400 277.200 327.000 ;
        RECT 287.400 326.400 290.400 330.000 ;
        RECT 478.800 329.400 482.400 330.000 ;
        RECT 517.200 329.400 520.800 330.000 ;
        RECT 479.400 327.600 482.400 329.400 ;
        RECT 517.800 328.800 520.800 329.400 ;
        RECT 578.400 329.400 581.400 330.600 ;
        RECT 688.200 330.000 691.800 331.200 ;
        RECT 675.000 329.400 687.000 330.000 ;
        RECT 688.200 329.400 692.400 330.000 ;
        RECT 578.400 328.800 582.000 329.400 ;
        RECT 670.800 328.800 692.400 329.400 ;
        RECT 517.800 328.200 521.400 328.800 ;
        RECT 518.400 327.600 521.400 328.200 ;
        RECT 579.000 327.600 582.000 328.800 ;
        RECT 669.600 328.200 692.400 328.800 ;
        RECT 669.000 327.600 693.000 328.200 ;
        RECT 479.400 327.000 483.000 327.600 ;
        RECT 518.400 327.000 522.000 327.600 ;
        RECT 579.000 327.000 582.600 327.600 ;
        RECT 113.400 325.800 117.600 326.400 ;
        RECT 219.600 325.800 231.000 326.400 ;
        RECT 264.600 325.800 268.200 326.400 ;
        RECT 113.400 325.200 117.000 325.800 ;
        RECT 221.400 325.200 230.400 325.800 ;
        RECT 265.200 325.200 268.200 325.800 ;
        RECT 112.800 324.600 116.400 325.200 ;
        RECT 222.600 324.600 229.800 325.200 ;
        RECT 265.200 324.600 268.800 325.200 ;
        RECT 273.600 324.600 276.600 326.400 ;
        RECT 112.200 323.400 115.800 324.600 ;
        RECT 223.800 324.000 229.800 324.600 ;
        RECT 265.800 324.000 269.400 324.600 ;
        RECT 225.000 323.400 229.800 324.000 ;
        RECT 266.400 323.400 269.400 324.000 ;
        RECT 111.600 322.800 115.200 323.400 ;
        RECT 225.600 322.800 230.400 323.400 ;
        RECT 266.400 322.800 270.000 323.400 ;
        RECT 111.600 322.200 114.600 322.800 ;
        RECT 226.800 322.200 231.600 322.800 ;
        RECT 267.000 322.200 270.000 322.800 ;
        RECT 273.000 322.200 276.000 324.600 ;
        RECT 111.000 321.600 114.600 322.200 ;
        RECT 227.400 321.600 232.200 322.200 ;
        RECT 267.000 321.600 270.600 322.200 ;
        RECT 111.000 321.000 114.000 321.600 ;
        RECT 228.000 321.000 232.800 321.600 ;
        RECT 267.600 321.000 270.600 321.600 ;
        RECT 110.400 319.800 113.400 321.000 ;
        RECT 153.600 320.400 156.600 321.000 ;
        RECT 229.200 320.400 233.400 321.000 ;
        RECT 267.600 320.400 271.200 321.000 ;
        RECT 152.400 319.800 159.000 320.400 ;
        RECT 229.800 319.800 234.000 320.400 ;
        RECT 109.800 318.600 112.800 319.800 ;
        RECT 151.800 319.200 161.400 319.800 ;
        RECT 230.400 319.200 234.600 319.800 ;
        RECT 268.200 319.200 271.200 320.400 ;
        RECT 272.400 319.200 275.400 322.200 ;
        RECT 288.000 321.600 291.000 326.400 ;
        RECT 303.600 325.800 306.000 326.400 ;
        RECT 302.400 325.200 307.200 325.800 ;
        RECT 480.000 325.200 483.000 327.000 ;
        RECT 519.000 325.800 522.000 327.000 ;
        RECT 579.600 325.800 582.600 327.000 ;
        RECT 668.400 327.000 693.000 327.600 ;
        RECT 668.400 325.800 678.600 327.000 ;
        RECT 684.000 326.400 693.000 327.000 ;
        RECT 687.000 325.800 693.000 326.400 ;
        RECT 301.800 324.600 307.800 325.200 ;
        RECT 480.000 324.600 483.600 325.200 ;
        RECT 301.200 323.400 308.400 324.600 ;
        RECT 480.600 323.400 483.600 324.600 ;
        RECT 519.600 324.600 522.600 325.800 ;
        RECT 579.600 325.200 583.200 325.800 ;
        RECT 669.600 325.200 681.000 325.800 ;
        RECT 688.800 325.200 693.000 325.800 ;
        RECT 519.600 324.000 523.200 324.600 ;
        RECT 580.200 324.000 583.200 325.200 ;
        RECT 671.400 324.600 682.800 325.200 ;
        RECT 690.600 324.600 692.400 325.200 ;
        RECT 673.800 324.000 684.600 324.600 ;
        RECT 520.200 323.400 523.200 324.000 ;
        RECT 300.600 322.800 304.200 323.400 ;
        RECT 305.400 322.800 309.000 323.400 ;
        RECT 300.000 322.200 303.600 322.800 ;
        RECT 306.000 322.200 309.600 322.800 ;
        RECT 480.600 322.200 484.200 323.400 ;
        RECT 520.200 322.800 523.800 323.400 ;
        RECT 154.800 318.600 162.600 319.200 ;
        RECT 231.000 318.600 235.200 319.200 ;
        RECT 109.200 318.000 112.800 318.600 ;
        RECT 156.600 318.000 164.400 318.600 ;
        RECT 231.600 318.000 235.200 318.600 ;
        RECT 268.800 318.600 275.400 319.200 ;
        RECT 109.200 316.800 112.200 318.000 ;
        RECT 158.400 317.400 166.200 318.000 ;
        RECT 232.200 317.400 235.800 318.000 ;
        RECT 268.800 317.400 274.800 318.600 ;
        RECT 160.200 316.800 167.400 317.400 ;
        RECT 232.800 316.800 236.400 317.400 ;
        RECT 108.600 315.000 111.600 316.800 ;
        RECT 161.400 316.200 168.600 316.800 ;
        RECT 163.200 315.600 170.400 316.200 ;
        RECT 233.400 315.600 237.000 316.800 ;
        RECT 269.400 315.600 274.800 317.400 ;
        RECT 164.400 315.000 171.600 315.600 ;
        RECT 234.000 315.000 237.600 315.600 ;
        RECT 108.600 313.800 111.000 315.000 ;
        RECT 165.600 314.400 172.800 315.000 ;
        RECT 234.600 314.400 237.600 315.000 ;
        RECT 270.000 314.400 274.200 315.600 ;
        RECT 288.600 315.000 291.600 321.600 ;
        RECT 299.400 321.000 303.000 322.200 ;
        RECT 306.600 321.000 309.600 322.200 ;
        RECT 481.200 321.600 484.200 322.200 ;
        RECT 520.800 322.200 523.800 322.800 ;
        RECT 580.800 322.800 583.800 324.000 ;
        RECT 676.200 323.400 685.800 324.000 ;
        RECT 678.600 322.800 687.000 323.400 ;
        RECT 580.800 322.200 584.400 322.800 ;
        RECT 681.000 322.200 688.200 322.800 ;
        RECT 520.800 321.600 524.400 322.200 ;
        RECT 298.800 320.400 302.400 321.000 ;
        RECT 306.600 320.400 310.200 321.000 ;
        RECT 481.200 320.400 484.800 321.600 ;
        RECT 521.400 321.000 524.400 321.600 ;
        RECT 581.400 321.600 584.400 322.200 ;
        RECT 682.800 321.600 688.800 322.200 ;
        RECT 521.400 320.400 525.000 321.000 ;
        RECT 581.400 320.400 585.000 321.600 ;
        RECT 684.000 321.000 690.000 321.600 ;
        RECT 685.200 320.400 690.600 321.000 ;
        RECT 298.800 319.800 301.800 320.400 ;
        RECT 298.200 319.200 301.800 319.800 ;
        RECT 307.200 319.200 310.200 320.400 ;
        RECT 481.800 319.200 484.800 320.400 ;
        RECT 522.000 319.800 525.000 320.400 ;
        RECT 582.000 319.800 585.000 320.400 ;
        RECT 686.400 319.800 691.200 320.400 ;
        RECT 522.000 319.200 525.600 319.800 ;
        RECT 582.000 319.200 585.600 319.800 ;
        RECT 687.600 319.200 691.800 319.800 ;
        RECT 297.600 318.000 301.200 319.200 ;
        RECT 297.000 317.400 300.600 318.000 ;
        RECT 297.000 316.800 300.000 317.400 ;
        RECT 307.800 316.800 310.800 319.200 ;
        RECT 481.800 318.600 485.400 319.200 ;
        RECT 522.600 318.600 525.600 319.200 ;
        RECT 582.600 318.600 585.600 319.200 ;
        RECT 688.200 318.600 691.800 319.200 ;
        RECT 482.400 317.400 485.400 318.600 ;
        RECT 523.200 318.000 526.200 318.600 ;
        RECT 523.200 317.400 526.800 318.000 ;
        RECT 582.600 317.400 586.200 318.600 ;
        RECT 622.200 317.400 623.400 318.000 ;
        RECT 688.800 317.400 691.800 318.600 ;
        RECT 482.400 316.800 486.000 317.400 ;
        RECT 296.400 316.200 300.000 316.800 ;
        RECT 296.400 315.600 299.400 316.200 ;
        RECT 166.800 313.800 174.000 314.400 ;
        RECT 234.600 313.800 238.200 314.400 ;
        RECT 270.000 313.800 273.600 314.400 ;
        RECT 108.000 312.000 111.000 313.800 ;
        RECT 168.600 313.200 175.200 313.800 ;
        RECT 235.200 313.200 238.200 313.800 ;
        RECT 169.800 312.600 176.400 313.200 ;
        RECT 171.000 312.000 177.600 312.600 ;
        RECT 235.800 312.000 238.800 313.200 ;
        RECT 108.600 310.800 111.000 312.000 ;
        RECT 172.200 311.400 178.800 312.000 ;
        RECT 235.800 311.400 239.400 312.000 ;
        RECT 173.400 310.800 180.000 311.400 ;
        RECT 236.400 310.800 239.400 311.400 ;
        RECT 108.600 307.200 111.600 310.800 ;
        RECT 174.600 310.200 181.200 310.800 ;
        RECT 236.400 310.200 240.000 310.800 ;
        RECT 270.600 310.200 273.600 313.800 ;
        RECT 175.800 309.600 182.400 310.200 ;
        RECT 177.000 309.000 183.600 309.600 ;
        RECT 237.000 309.000 240.000 310.200 ;
        RECT 271.200 309.600 273.600 310.200 ;
        RECT 289.200 313.800 291.600 315.000 ;
        RECT 295.800 315.000 299.400 315.600 ;
        RECT 295.800 314.400 298.800 315.000 ;
        RECT 295.200 313.800 298.800 314.400 ;
        RECT 308.400 313.800 311.400 316.800 ;
        RECT 483.000 315.000 486.000 316.800 ;
        RECT 523.800 316.800 526.800 317.400 ;
        RECT 583.200 316.800 586.200 317.400 ;
        RECT 613.800 316.800 624.600 317.400 ;
        RECT 523.800 316.200 527.400 316.800 ;
        RECT 583.200 316.200 586.800 316.800 ;
        RECT 610.200 316.200 624.600 316.800 ;
        RECT 524.400 315.600 527.400 316.200 ;
        RECT 524.400 315.000 528.000 315.600 ;
        RECT 583.800 315.000 586.800 316.200 ;
        RECT 606.600 315.600 624.600 316.200 ;
        RECT 603.600 315.000 624.600 315.600 ;
        RECT 289.200 309.600 292.200 313.800 ;
        RECT 295.200 313.200 298.200 313.800 ;
        RECT 294.600 312.600 298.200 313.200 ;
        RECT 309.000 313.200 311.400 313.800 ;
        RECT 483.600 313.200 486.600 315.000 ;
        RECT 525.000 313.800 528.600 315.000 ;
        RECT 584.400 313.800 587.400 315.000 ;
        RECT 601.200 314.400 623.400 315.000 ;
        RECT 689.400 314.400 692.400 317.400 ;
        RECT 598.800 313.800 621.600 314.400 ;
        RECT 525.600 313.200 529.200 313.800 ;
        RECT 584.400 313.200 588.000 313.800 ;
        RECT 597.000 313.200 609.600 313.800 ;
        RECT 613.200 313.200 620.400 313.800 ;
        RECT 294.600 312.000 297.600 312.600 ;
        RECT 294.000 311.400 297.600 312.000 ;
        RECT 294.000 310.800 297.000 311.400 ;
        RECT 293.400 310.200 297.000 310.800 ;
        RECT 293.400 309.600 296.400 310.200 ;
        RECT 178.200 308.400 184.800 309.000 ;
        RECT 237.000 308.400 240.600 309.000 ;
        RECT 179.400 307.800 185.400 308.400 ;
        RECT 180.600 307.200 186.600 307.800 ;
        RECT 109.200 304.800 112.200 307.200 ;
        RECT 181.800 306.600 187.800 307.200 ;
        RECT 237.600 306.600 240.600 308.400 ;
        RECT 183.000 306.000 189.000 306.600 ;
        RECT 184.200 305.400 189.600 306.000 ;
        RECT 184.800 304.800 190.800 305.400 ;
        RECT 109.800 303.000 112.800 304.800 ;
        RECT 186.000 304.200 191.400 304.800 ;
        RECT 238.200 304.200 241.200 306.600 ;
        RECT 271.200 304.800 274.200 309.600 ;
        RECT 289.200 309.000 296.400 309.600 ;
        RECT 289.200 307.800 295.800 309.000 ;
        RECT 289.200 306.600 295.200 307.800 ;
        RECT 289.200 305.400 294.600 306.600 ;
        RECT 271.200 304.200 273.600 304.800 ;
        RECT 187.200 303.600 192.600 304.200 ;
        RECT 187.800 303.000 193.800 303.600 ;
        RECT 110.400 301.800 113.400 303.000 ;
        RECT 189.000 302.400 194.400 303.000 ;
        RECT 190.200 301.800 195.600 302.400 ;
        RECT 110.400 301.200 114.000 301.800 ;
        RECT 190.800 301.200 196.200 301.800 ;
        RECT 111.000 300.600 114.000 301.200 ;
        RECT 192.000 300.600 196.800 301.200 ;
        RECT 238.800 300.600 241.800 304.200 ;
        RECT 270.600 301.200 273.600 304.200 ;
        RECT 289.200 304.200 294.000 305.400 ;
        RECT 289.200 303.000 293.400 304.200 ;
        RECT 289.200 301.800 292.800 303.000 ;
        RECT 111.000 299.400 114.600 300.600 ;
        RECT 192.600 300.000 198.000 300.600 ;
        RECT 239.400 300.000 241.800 300.600 ;
        RECT 193.800 299.400 198.600 300.000 ;
        RECT 111.600 298.200 115.200 299.400 ;
        RECT 194.400 298.800 199.200 299.400 ;
        RECT 195.600 298.200 200.400 298.800 ;
        RECT 112.200 297.600 115.800 298.200 ;
        RECT 196.200 297.600 201.000 298.200 ;
        RECT 112.800 297.000 116.400 297.600 ;
        RECT 196.800 297.000 201.600 297.600 ;
        RECT 112.800 296.400 117.000 297.000 ;
        RECT 198.000 296.400 202.800 297.000 ;
        RECT 113.400 295.200 117.600 296.400 ;
        RECT 198.600 295.800 203.400 296.400 ;
        RECT 199.200 295.200 205.200 295.800 ;
        RECT 105.000 294.600 118.800 295.200 ;
        RECT 200.400 294.600 206.400 295.200 ;
        RECT 100.800 294.000 123.000 294.600 ;
        RECT 201.000 294.000 207.600 294.600 ;
        RECT 99.000 293.400 126.000 294.000 ;
        RECT 201.600 293.400 208.800 294.000 ;
        RECT 97.200 292.800 129.000 293.400 ;
        RECT 202.200 292.800 210.000 293.400 ;
        RECT 96.600 292.200 131.400 292.800 ;
        RECT 202.800 292.200 210.600 292.800 ;
        RECT 96.000 291.600 104.400 292.200 ;
        RECT 119.400 291.600 133.200 292.200 ;
        RECT 203.400 291.600 211.800 292.200 ;
        RECT 95.400 291.000 100.800 291.600 ;
        RECT 123.600 291.000 134.400 291.600 ;
        RECT 204.000 291.000 213.000 291.600 ;
        RECT 95.400 290.400 99.000 291.000 ;
        RECT 126.600 290.400 135.600 291.000 ;
        RECT 204.600 290.400 214.200 291.000 ;
        RECT 95.400 289.200 98.400 290.400 ;
        RECT 129.000 289.800 136.200 290.400 ;
        RECT 205.200 289.800 214.800 290.400 ;
        RECT 239.400 289.800 242.400 300.000 ;
        RECT 270.000 299.400 273.000 301.200 ;
        RECT 289.200 300.600 292.200 301.800 ;
        RECT 288.600 299.400 291.600 300.600 ;
        RECT 269.400 298.200 272.400 299.400 ;
        RECT 288.000 298.200 291.000 299.400 ;
        RECT 268.800 297.600 272.400 298.200 ;
        RECT 287.400 297.600 291.000 298.200 ;
        RECT 268.800 297.000 273.000 297.600 ;
        RECT 287.400 297.000 290.400 297.600 ;
        RECT 309.000 297.000 312.000 313.200 ;
        RECT 484.200 312.000 487.200 313.200 ;
        RECT 526.200 312.600 529.200 313.200 ;
        RECT 526.200 312.000 529.800 312.600 ;
        RECT 484.200 311.400 487.800 312.000 ;
        RECT 484.800 310.200 487.800 311.400 ;
        RECT 526.800 311.400 529.800 312.000 ;
        RECT 585.000 312.000 588.000 313.200 ;
        RECT 595.200 312.600 606.600 313.200 ;
        RECT 613.200 312.600 619.200 313.200 ;
        RECT 593.400 312.000 603.600 312.600 ;
        RECT 612.000 312.000 618.000 312.600 ;
        RECT 585.000 311.400 588.600 312.000 ;
        RECT 591.600 311.400 601.200 312.000 ;
        RECT 611.400 311.400 616.800 312.000 ;
        RECT 690.000 311.400 693.000 314.400 ;
        RECT 526.800 310.800 530.400 311.400 ;
        RECT 527.400 310.200 530.400 310.800 ;
        RECT 585.600 310.800 588.600 311.400 ;
        RECT 590.400 310.800 598.800 311.400 ;
        RECT 610.200 310.800 616.200 311.400 ;
        RECT 585.600 310.200 597.000 310.800 ;
        RECT 609.000 310.200 615.000 310.800 ;
        RECT 484.800 309.600 488.400 310.200 ;
        RECT 527.400 309.600 531.000 310.200 ;
        RECT 586.200 309.600 595.200 310.200 ;
        RECT 608.400 309.600 613.800 310.200 ;
        RECT 485.400 309.000 488.400 309.600 ;
        RECT 528.000 309.000 531.600 309.600 ;
        RECT 586.200 309.000 593.400 309.600 ;
        RECT 607.200 309.000 612.600 309.600 ;
        RECT 485.400 308.400 489.000 309.000 ;
        RECT 486.000 307.200 489.000 308.400 ;
        RECT 528.600 308.400 531.600 309.000 ;
        RECT 586.800 308.400 592.200 309.000 ;
        RECT 606.600 308.400 612.000 309.000 ;
        RECT 690.600 308.400 693.600 311.400 ;
        RECT 528.600 307.800 532.200 308.400 ;
        RECT 587.400 307.800 590.400 308.400 ;
        RECT 605.400 307.800 610.800 308.400 ;
        RECT 691.200 307.800 693.600 308.400 ;
        RECT 486.600 306.000 489.600 307.200 ;
        RECT 529.200 306.600 532.800 307.800 ;
        RECT 604.200 307.200 610.200 307.800 ;
        RECT 603.600 306.600 609.000 307.200 ;
        RECT 529.800 306.000 533.400 306.600 ;
        RECT 602.400 306.000 607.800 306.600 ;
        RECT 486.600 305.400 490.200 306.000 ;
        RECT 487.200 304.800 490.200 305.400 ;
        RECT 530.400 305.400 533.400 306.000 ;
        RECT 601.800 305.400 607.200 306.000 ;
        RECT 530.400 304.800 534.000 305.400 ;
        RECT 600.600 304.800 606.000 305.400 ;
        RECT 487.200 304.200 490.800 304.800 ;
        RECT 487.800 303.600 490.800 304.200 ;
        RECT 531.000 303.600 534.600 304.800 ;
        RECT 600.000 304.200 605.400 304.800 ;
        RECT 691.200 304.200 694.200 307.800 ;
        RECT 598.800 303.600 604.200 304.200 ;
        RECT 691.800 303.600 694.200 304.200 ;
        RECT 487.800 303.000 491.400 303.600 ;
        RECT 531.600 303.000 535.200 303.600 ;
        RECT 597.600 303.000 603.000 303.600 ;
        RECT 488.400 301.800 491.400 303.000 ;
        RECT 532.200 301.800 535.800 303.000 ;
        RECT 597.000 302.400 602.400 303.000 ;
        RECT 595.800 301.800 601.200 302.400 ;
        RECT 489.000 300.600 492.000 301.800 ;
        RECT 532.800 301.200 536.400 301.800 ;
        RECT 595.200 301.200 600.600 301.800 ;
        RECT 533.400 300.600 536.400 301.200 ;
        RECT 594.000 300.600 599.400 301.200 ;
        RECT 489.000 300.000 492.600 300.600 ;
        RECT 533.400 300.000 537.000 300.600 ;
        RECT 592.800 300.000 598.800 300.600 ;
        RECT 489.600 299.400 492.600 300.000 ;
        RECT 534.000 299.400 537.600 300.000 ;
        RECT 592.200 299.400 597.600 300.000 ;
        RECT 489.600 298.800 493.200 299.400 ;
        RECT 490.200 298.200 493.200 298.800 ;
        RECT 534.600 298.800 537.600 299.400 ;
        RECT 591.000 298.800 596.400 299.400 ;
        RECT 534.600 298.200 538.200 298.800 ;
        RECT 590.400 298.200 595.800 298.800 ;
        RECT 691.800 298.200 694.800 303.600 ;
        RECT 490.200 297.600 493.800 298.200 ;
        RECT 490.800 297.000 493.800 297.600 ;
        RECT 535.200 297.000 538.800 298.200 ;
        RECT 589.200 297.600 594.600 298.200 ;
        RECT 692.400 297.600 694.800 298.200 ;
        RECT 588.600 297.000 594.000 297.600 ;
        RECT 268.200 296.400 273.000 297.000 ;
        RECT 286.800 296.400 290.400 297.000 ;
        RECT 268.200 295.800 273.600 296.400 ;
        RECT 267.600 294.600 274.200 295.800 ;
        RECT 286.800 295.200 289.800 296.400 ;
        RECT 267.000 294.000 274.800 294.600 ;
        RECT 286.200 294.000 289.200 295.200 ;
        RECT 266.400 293.400 270.000 294.000 ;
        RECT 265.800 292.800 270.000 293.400 ;
        RECT 271.800 292.800 274.800 294.000 ;
        RECT 285.600 293.400 289.200 294.000 ;
        RECT 265.200 292.200 269.400 292.800 ;
        RECT 264.600 291.600 268.800 292.200 ;
        RECT 272.400 291.600 275.400 292.800 ;
        RECT 285.600 292.200 288.600 293.400 ;
        RECT 308.400 292.200 311.400 297.000 ;
        RECT 490.800 296.400 494.400 297.000 ;
        RECT 535.800 296.400 539.400 297.000 ;
        RECT 587.400 296.400 592.800 297.000 ;
        RECT 491.400 295.800 494.400 296.400 ;
        RECT 491.400 295.200 495.000 295.800 ;
        RECT 536.400 295.200 540.000 296.400 ;
        RECT 586.800 295.800 591.600 296.400 ;
        RECT 585.600 295.200 591.000 295.800 ;
        RECT 492.000 294.600 495.000 295.200 ;
        RECT 537.000 294.600 540.600 295.200 ;
        RECT 585.000 294.600 589.800 295.200 ;
        RECT 492.000 294.000 495.600 294.600 ;
        RECT 492.600 293.400 496.200 294.000 ;
        RECT 537.600 293.400 541.200 294.600 ;
        RECT 585.000 293.400 589.200 294.600 ;
        RECT 493.200 292.800 496.200 293.400 ;
        RECT 538.200 292.800 541.800 293.400 ;
        RECT 585.000 292.800 589.800 293.400 ;
        RECT 493.200 292.200 496.800 292.800 ;
        RECT 264.000 291.000 268.200 291.600 ;
        RECT 272.400 291.000 276.000 291.600 ;
        RECT 285.000 291.000 288.000 292.200 ;
        RECT 263.400 290.400 267.600 291.000 ;
        RECT 262.800 289.800 267.600 290.400 ;
        RECT 273.000 289.800 276.000 291.000 ;
        RECT 284.400 290.400 288.000 291.000 ;
        RECT 130.800 289.200 136.800 289.800 ;
        RECT 205.800 289.200 216.000 289.800 ;
        RECT 239.400 289.200 241.800 289.800 ;
        RECT 261.600 289.200 267.000 289.800 ;
        RECT 95.400 288.600 99.000 289.200 ;
        RECT 133.200 288.600 136.800 289.200 ;
        RECT 206.400 288.600 217.200 289.200 ;
        RECT 96.000 287.400 99.600 288.600 ;
        RECT 135.000 288.000 136.200 288.600 ;
        RECT 207.000 288.000 211.200 288.600 ;
        RECT 212.400 288.000 218.400 288.600 ;
        RECT 207.600 287.400 211.200 288.000 ;
        RECT 213.600 287.400 219.000 288.000 ;
        RECT 96.600 286.800 100.800 287.400 ;
        RECT 208.200 286.800 211.800 287.400 ;
        RECT 214.200 286.800 220.200 287.400 ;
        RECT 97.200 286.200 101.400 286.800 ;
        RECT 208.800 286.200 212.400 286.800 ;
        RECT 215.400 286.200 221.400 286.800 ;
        RECT 238.800 286.200 241.800 289.200 ;
        RECT 261.000 288.600 266.400 289.200 ;
        RECT 273.600 288.600 276.600 289.800 ;
        RECT 284.400 289.200 287.400 290.400 ;
        RECT 260.400 288.000 265.800 288.600 ;
        RECT 273.600 288.000 277.200 288.600 ;
        RECT 283.800 288.000 286.800 289.200 ;
        RECT 307.800 288.600 310.800 292.200 ;
        RECT 493.800 291.600 496.800 292.200 ;
        RECT 538.800 291.600 542.400 292.800 ;
        RECT 585.600 292.200 590.400 292.800 ;
        RECT 586.200 291.600 591.000 292.200 ;
        RECT 493.800 291.000 497.400 291.600 ;
        RECT 539.400 291.000 543.000 291.600 ;
        RECT 587.400 291.000 591.600 291.600 ;
        RECT 494.400 290.400 497.400 291.000 ;
        RECT 494.400 289.800 498.000 290.400 ;
        RECT 540.000 289.800 543.600 291.000 ;
        RECT 588.000 290.400 592.200 291.000 ;
        RECT 588.600 289.800 592.800 290.400 ;
        RECT 495.000 289.200 498.000 289.800 ;
        RECT 540.600 289.200 544.200 289.800 ;
        RECT 589.200 289.200 593.400 289.800 ;
        RECT 495.000 288.600 498.600 289.200 ;
        RECT 259.800 287.400 265.200 288.000 ;
        RECT 259.200 286.800 264.000 287.400 ;
        RECT 274.200 286.800 277.200 288.000 ;
        RECT 283.200 287.400 286.800 288.000 ;
        RECT 258.000 286.200 263.400 286.800 ;
        RECT 274.200 286.200 277.800 286.800 ;
        RECT 283.200 286.200 286.200 287.400 ;
        RECT 97.800 285.600 102.000 286.200 ;
        RECT 209.400 285.600 212.400 286.200 ;
        RECT 216.600 285.600 222.600 286.200 ;
        RECT 98.400 285.000 102.600 285.600 ;
        RECT 99.000 284.400 103.800 285.000 ;
        RECT 210.000 284.400 213.000 285.600 ;
        RECT 217.800 285.000 223.200 285.600 ;
        RECT 238.200 285.000 241.200 286.200 ;
        RECT 257.400 285.600 262.800 286.200 ;
        RECT 256.200 285.000 262.200 285.600 ;
        RECT 274.800 285.000 277.800 286.200 ;
        RECT 218.400 284.400 224.400 285.000 ;
        RECT 99.600 283.800 104.400 284.400 ;
        RECT 210.600 283.800 213.600 284.400 ;
        RECT 219.600 283.800 225.600 284.400 ;
        RECT 237.600 283.800 241.200 285.000 ;
        RECT 255.000 284.400 261.000 285.000 ;
        RECT 274.800 284.400 278.400 285.000 ;
        RECT 282.600 284.400 285.600 286.200 ;
        RECT 307.200 285.600 310.200 288.600 ;
        RECT 495.600 288.000 499.200 288.600 ;
        RECT 541.200 288.000 544.800 289.200 ;
        RECT 589.800 288.600 594.000 289.200 ;
        RECT 590.400 288.000 594.600 288.600 ;
        RECT 496.200 287.400 499.200 288.000 ;
        RECT 541.800 287.400 545.400 288.000 ;
        RECT 591.000 287.400 595.200 288.000 ;
        RECT 496.200 286.800 499.800 287.400 ;
        RECT 496.800 286.200 499.800 286.800 ;
        RECT 542.400 286.200 546.000 287.400 ;
        RECT 591.600 286.800 595.800 287.400 ;
        RECT 592.200 286.200 596.400 286.800 ;
        RECT 496.800 285.600 500.400 286.200 ;
        RECT 543.000 285.600 546.600 286.200 ;
        RECT 592.800 285.600 597.600 286.200 ;
        RECT 253.800 283.800 260.400 284.400 ;
        RECT 100.200 283.200 105.600 283.800 ;
        RECT 211.200 283.200 213.600 283.800 ;
        RECT 220.800 283.200 226.200 283.800 ;
        RECT 237.600 283.200 240.600 283.800 ;
        RECT 252.600 283.200 259.200 283.800 ;
        RECT 100.800 282.600 106.200 283.200 ;
        RECT 211.800 282.600 214.200 283.200 ;
        RECT 221.400 282.600 227.400 283.200 ;
        RECT 237.000 282.600 240.600 283.200 ;
        RECT 251.400 282.600 258.000 283.200 ;
        RECT 275.400 282.600 278.400 284.400 ;
        RECT 282.000 283.200 285.000 284.400 ;
        RECT 306.600 283.200 309.600 285.600 ;
        RECT 497.400 285.000 501.000 285.600 ;
        RECT 543.600 285.000 547.200 285.600 ;
        RECT 593.400 285.000 598.200 285.600 ;
        RECT 498.000 284.400 501.000 285.000 ;
        RECT 544.200 284.400 547.200 285.000 ;
        RECT 594.600 284.400 598.800 285.000 ;
        RECT 498.000 283.800 501.600 284.400 ;
        RECT 544.200 283.800 547.800 284.400 ;
        RECT 595.200 283.800 599.400 284.400 ;
        RECT 498.600 283.200 501.600 283.800 ;
        RECT 544.800 283.200 548.400 283.800 ;
        RECT 595.800 283.200 600.000 283.800 ;
        RECT 281.400 282.600 285.000 283.200 ;
        RECT 102.000 282.000 107.400 282.600 ;
        RECT 212.400 282.000 214.200 282.600 ;
        RECT 222.600 282.000 228.000 282.600 ;
        RECT 237.000 282.000 240.000 282.600 ;
        RECT 250.200 282.000 256.800 282.600 ;
        RECT 102.600 281.400 108.600 282.000 ;
        RECT 103.800 280.800 109.200 281.400 ;
        RECT 213.000 280.800 214.800 282.000 ;
        RECT 223.800 281.400 229.200 282.000 ;
        RECT 224.400 280.800 230.400 281.400 ;
        RECT 236.400 280.800 240.000 282.000 ;
        RECT 248.400 281.400 255.600 282.000 ;
        RECT 247.200 280.800 255.000 281.400 ;
        RECT 104.400 280.200 110.400 280.800 ;
        RECT 213.600 280.200 214.800 280.800 ;
        RECT 225.600 280.200 231.000 280.800 ;
        RECT 236.400 280.200 239.400 280.800 ;
        RECT 105.600 279.600 112.200 280.200 ;
        RECT 214.200 279.600 215.400 280.200 ;
        RECT 226.800 279.600 232.200 280.200 ;
        RECT 235.800 279.600 239.400 280.200 ;
        RECT 246.000 280.200 253.800 280.800 ;
        RECT 276.000 280.200 279.000 282.600 ;
        RECT 281.400 281.400 284.400 282.600 ;
        RECT 246.000 279.600 252.600 280.200 ;
        RECT 276.600 279.600 279.600 280.200 ;
        RECT 280.800 279.600 283.800 281.400 ;
        RECT 306.000 280.800 309.000 283.200 ;
        RECT 498.600 282.600 502.200 283.200 ;
        RECT 499.200 282.000 502.800 282.600 ;
        RECT 545.400 282.000 549.000 283.200 ;
        RECT 596.400 282.600 600.600 283.200 ;
        RECT 597.000 282.000 601.200 282.600 ;
        RECT 692.400 282.000 695.400 297.600 ;
        RECT 499.800 281.400 502.800 282.000 ;
        RECT 546.000 281.400 549.600 282.000 ;
        RECT 597.600 281.400 601.800 282.000 ;
        RECT 499.800 280.800 503.400 281.400 ;
        RECT 106.800 279.000 113.400 279.600 ;
        RECT 214.800 279.000 215.400 279.600 ;
        RECT 227.400 279.000 232.800 279.600 ;
        RECT 235.800 279.000 238.800 279.600 ;
        RECT 246.000 279.000 250.800 279.600 ;
        RECT 108.000 278.400 114.600 279.000 ;
        RECT 228.600 278.400 234.000 279.000 ;
        RECT 235.200 278.400 238.800 279.000 ;
        RECT 246.600 278.400 249.600 279.000 ;
        RECT 109.200 277.800 116.400 278.400 ;
        RECT 229.200 277.800 238.200 278.400 ;
        RECT 110.400 277.200 118.200 277.800 ;
        RECT 230.400 277.200 238.200 277.800 ;
        RECT 247.200 277.800 249.600 278.400 ;
        RECT 276.600 277.800 283.200 279.600 ;
        RECT 305.400 278.400 308.400 280.800 ;
        RECT 500.400 280.200 503.400 280.800 ;
        RECT 546.600 280.200 550.200 281.400 ;
        RECT 598.200 280.800 602.400 281.400 ;
        RECT 692.400 280.800 694.800 282.000 ;
        RECT 598.800 280.200 603.000 280.800 ;
        RECT 500.400 279.600 504.000 280.200 ;
        RECT 547.200 279.600 550.800 280.200 ;
        RECT 599.400 279.600 603.600 280.200 ;
        RECT 501.000 279.000 504.600 279.600 ;
        RECT 547.800 279.000 551.400 279.600 ;
        RECT 600.000 279.000 604.200 279.600 ;
        RECT 501.600 278.400 504.600 279.000 ;
        RECT 247.200 277.200 250.200 277.800 ;
        RECT 111.600 276.600 119.400 277.200 ;
        RECT 231.000 276.600 238.200 277.200 ;
        RECT 112.800 276.000 121.800 276.600 ;
        RECT 232.200 276.000 238.200 276.600 ;
        RECT 114.600 275.400 123.600 276.000 ;
        RECT 232.800 275.400 238.200 276.000 ;
        RECT 247.800 276.600 250.200 277.200 ;
        RECT 247.800 275.400 250.800 276.600 ;
        RECT 277.200 276.000 282.600 277.800 ;
        RECT 304.800 276.000 307.800 278.400 ;
        RECT 501.600 277.800 505.200 278.400 ;
        RECT 548.400 277.800 552.000 279.000 ;
        RECT 600.600 278.400 605.400 279.000 ;
        RECT 601.200 277.800 606.000 278.400 ;
        RECT 502.200 277.200 505.800 277.800 ;
        RECT 549.000 277.200 552.600 277.800 ;
        RECT 601.800 277.200 606.600 277.800 ;
        RECT 502.200 276.600 506.400 277.200 ;
        RECT 502.800 276.000 506.400 276.600 ;
        RECT 549.600 276.000 553.200 277.200 ;
        RECT 603.000 276.600 607.200 277.200 ;
        RECT 603.600 276.000 607.800 276.600 ;
        RECT 277.200 275.400 282.000 276.000 ;
        RECT 115.800 274.800 126.000 275.400 ;
        RECT 234.000 274.800 239.400 275.400 ;
        RECT 117.600 274.200 128.400 274.800 ;
        RECT 234.600 274.200 240.000 274.800 ;
        RECT 248.400 274.200 251.400 275.400 ;
        RECT 277.800 274.800 282.000 275.400 ;
        RECT 119.400 273.600 130.800 274.200 ;
        RECT 235.800 273.600 240.600 274.200 ;
        RECT 248.400 273.600 252.000 274.200 ;
        RECT 121.200 273.000 133.200 273.600 ;
        RECT 236.400 273.000 241.800 273.600 ;
        RECT 122.400 272.400 135.600 273.000 ;
        RECT 237.600 272.400 242.400 273.000 ;
        RECT 249.000 272.400 252.000 273.600 ;
        RECT 277.800 273.000 281.400 274.800 ;
        RECT 304.200 274.200 307.200 276.000 ;
        RECT 503.400 274.800 507.000 276.000 ;
        RECT 550.200 275.400 553.800 276.000 ;
        RECT 604.200 275.400 608.400 276.000 ;
        RECT 550.800 274.800 554.400 275.400 ;
        RECT 604.800 274.800 609.000 275.400 ;
        RECT 691.800 274.800 694.800 280.800 ;
        RECT 504.000 274.200 507.600 274.800 ;
        RECT 124.800 271.800 138.600 272.400 ;
        RECT 238.200 271.800 243.000 272.400 ;
        RECT 126.600 271.200 141.000 271.800 ;
        RECT 239.400 271.200 244.200 271.800 ;
        RECT 249.600 271.200 252.600 272.400 ;
        RECT 126.600 270.600 154.200 271.200 ;
        RECT 240.000 270.600 244.800 271.200 ;
        RECT 114.000 270.000 159.600 270.600 ;
        RECT 240.600 270.000 246.000 270.600 ;
        RECT 250.200 270.000 253.200 271.200 ;
        RECT 278.400 270.000 281.400 273.000 ;
        RECT 303.600 273.600 307.200 274.200 ;
        RECT 303.600 271.800 306.600 273.600 ;
        RECT 504.600 273.000 508.200 274.200 ;
        RECT 551.400 273.600 555.000 274.800 ;
        RECT 605.400 274.200 609.600 274.800 ;
        RECT 606.000 273.600 610.200 274.200 ;
        RECT 552.000 273.000 555.600 273.600 ;
        RECT 606.600 273.000 610.800 273.600 ;
        RECT 505.200 272.400 508.800 273.000 ;
        RECT 303.000 270.000 306.000 271.800 ;
        RECT 505.800 271.200 509.400 272.400 ;
        RECT 552.600 271.800 556.200 273.000 ;
        RECT 607.200 272.400 611.400 273.000 ;
        RECT 607.800 271.800 612.600 272.400 ;
        RECT 553.200 271.200 556.800 271.800 ;
        RECT 608.400 271.200 613.200 271.800 ;
        RECT 506.400 270.600 510.000 271.200 ;
        RECT 553.800 270.600 557.400 271.200 ;
        RECT 609.600 270.600 613.800 271.200 ;
        RECT 691.200 270.600 694.200 274.800 ;
        RECT 507.000 270.000 510.000 270.600 ;
        RECT 106.200 269.400 160.200 270.000 ;
        RECT 241.800 269.400 246.600 270.000 ;
        RECT 250.800 269.400 253.800 270.000 ;
        RECT 100.200 268.800 160.800 269.400 ;
        RECT 242.400 268.800 247.200 269.400 ;
        RECT 250.800 268.800 254.400 269.400 ;
        RECT 95.400 268.200 160.800 268.800 ;
        RECT 243.000 268.200 247.800 268.800 ;
        RECT 251.400 268.200 254.400 268.800 ;
        RECT 91.200 267.600 126.000 268.200 ;
        RECT 156.000 267.600 160.200 268.200 ;
        RECT 244.200 267.600 249.000 268.200 ;
        RECT 251.400 267.600 255.000 268.200 ;
        RECT 87.600 267.000 112.800 267.600 ;
        RECT 244.800 267.000 249.600 267.600 ;
        RECT 252.000 267.000 255.000 267.600 ;
        RECT 84.000 266.400 105.600 267.000 ;
        RECT 245.400 266.400 250.200 267.000 ;
        RECT 81.000 265.800 99.600 266.400 ;
        RECT 246.600 265.800 250.800 266.400 ;
        RECT 252.000 265.800 255.600 267.000 ;
        RECT 279.000 266.400 282.000 270.000 ;
        RECT 302.400 268.200 305.400 270.000 ;
        RECT 507.000 269.400 510.600 270.000 ;
        RECT 554.400 269.400 558.000 270.600 ;
        RECT 610.200 270.000 614.400 270.600 ;
        RECT 691.200 270.000 693.600 270.600 ;
        RECT 610.800 269.400 615.000 270.000 ;
        RECT 507.600 268.800 511.200 269.400 ;
        RECT 555.000 268.800 558.600 269.400 ;
        RECT 611.400 268.800 615.600 269.400 ;
        RECT 301.800 267.600 305.400 268.200 ;
        RECT 508.200 268.200 511.200 268.800 ;
        RECT 555.600 268.200 559.200 268.800 ;
        RECT 612.000 268.200 616.200 268.800 ;
        RECT 508.200 267.600 511.800 268.200 ;
        RECT 301.800 266.400 304.800 267.600 ;
        RECT 508.800 267.000 511.800 267.600 ;
        RECT 556.200 267.000 559.800 268.200 ;
        RECT 612.600 267.600 616.800 268.200 ;
        RECT 613.200 267.000 617.400 267.600 ;
        RECT 314.400 266.400 327.000 267.000 ;
        RECT 508.800 266.400 512.400 267.000 ;
        RECT 556.800 266.400 560.400 267.000 ;
        RECT 613.800 266.400 618.000 267.000 ;
        RECT 690.600 266.400 693.600 270.000 ;
        RECT 279.600 265.800 282.000 266.400 ;
        RECT 301.200 265.800 304.800 266.400 ;
        RECT 309.000 265.800 331.800 266.400 ;
        RECT 509.400 265.800 513.000 266.400 ;
        RECT 78.600 265.200 94.800 265.800 ;
        RECT 247.200 265.200 256.200 265.800 ;
        RECT 76.200 264.600 91.200 265.200 ;
        RECT 247.800 264.600 256.800 265.200 ;
        RECT 74.400 264.000 87.000 264.600 ;
        RECT 248.400 264.000 256.800 264.600 ;
        RECT 72.600 263.400 84.000 264.000 ;
        RECT 249.600 263.400 257.400 264.000 ;
        RECT 70.800 262.800 81.000 263.400 ;
        RECT 250.200 262.800 258.000 263.400 ;
        RECT 69.600 262.200 78.600 262.800 ;
        RECT 250.800 262.200 258.000 262.800 ;
        RECT 68.400 261.600 76.200 262.200 ;
        RECT 251.400 261.600 258.600 262.200 ;
        RECT 67.800 261.000 74.400 261.600 ;
        RECT 252.600 261.000 259.200 261.600 ;
        RECT 67.200 260.400 72.600 261.000 ;
        RECT 253.200 260.400 259.800 261.000 ;
        RECT 66.600 259.800 71.400 260.400 ;
        RECT 253.800 259.800 259.800 260.400 ;
        RECT 279.600 259.800 282.600 265.800 ;
        RECT 301.200 265.200 334.200 265.800 ;
        RECT 510.000 265.200 513.000 265.800 ;
        RECT 557.400 265.800 561.000 266.400 ;
        RECT 614.400 265.800 618.600 266.400 ;
        RECT 557.400 265.200 561.600 265.800 ;
        RECT 615.000 265.200 619.200 265.800 ;
        RECT 301.200 264.600 336.600 265.200 ;
        RECT 510.000 264.600 513.600 265.200 ;
        RECT 558.000 264.600 561.600 265.200 ;
        RECT 615.600 264.600 619.800 265.200 ;
        RECT 300.000 264.000 339.000 264.600 ;
        RECT 510.600 264.000 513.600 264.600 ;
        RECT 558.600 264.000 562.200 264.600 ;
        RECT 616.200 264.000 620.400 264.600 ;
        RECT 297.600 263.400 313.800 264.000 ;
        RECT 327.600 263.400 340.800 264.000 ;
        RECT 510.600 263.400 514.200 264.000 ;
        RECT 559.200 263.400 562.800 264.000 ;
        RECT 616.800 263.400 621.000 264.000 ;
        RECT 690.000 263.400 693.000 266.400 ;
        RECT 295.200 262.800 308.400 263.400 ;
        RECT 331.800 262.800 342.600 263.400 ;
        RECT 511.200 262.800 514.800 263.400 ;
        RECT 559.200 262.800 563.400 263.400 ;
        RECT 617.400 262.800 621.600 263.400 ;
        RECT 690.000 262.800 692.400 263.400 ;
        RECT 292.800 262.200 305.400 262.800 ;
        RECT 334.800 262.200 344.400 262.800 ;
        RECT 511.800 262.200 514.800 262.800 ;
        RECT 559.800 262.200 563.400 262.800 ;
        RECT 618.000 262.200 622.200 262.800 ;
        RECT 291.000 261.600 301.800 262.200 ;
        RECT 336.600 261.600 346.200 262.200 ;
        RECT 511.800 261.600 515.400 262.200 ;
        RECT 288.600 261.000 299.400 261.600 ;
        RECT 339.000 261.000 347.400 261.600 ;
        RECT 512.400 261.000 515.400 261.600 ;
        RECT 560.400 261.600 564.000 262.200 ;
        RECT 618.600 261.600 622.800 262.200 ;
        RECT 560.400 261.000 564.600 261.600 ;
        RECT 619.200 261.000 623.400 261.600 ;
        RECT 286.800 260.400 297.600 261.000 ;
        RECT 340.800 260.400 348.600 261.000 ;
        RECT 512.400 260.400 516.000 261.000 ;
        RECT 561.000 260.400 564.600 261.000 ;
        RECT 619.800 260.400 624.000 261.000 ;
        RECT 285.000 259.800 295.200 260.400 ;
        RECT 342.600 259.800 349.800 260.400 ;
        RECT 513.000 259.800 516.000 260.400 ;
        RECT 561.600 259.800 565.200 260.400 ;
        RECT 620.400 259.800 624.600 260.400 ;
        RECT 689.400 259.800 692.400 262.800 ;
        RECT 66.600 259.200 70.200 259.800 ;
        RECT 254.400 259.200 260.400 259.800 ;
        RECT 280.200 259.200 292.800 259.800 ;
        RECT 343.800 259.200 351.000 259.800 ;
        RECT 513.000 259.200 516.600 259.800 ;
        RECT 562.200 259.200 565.800 259.800 ;
        RECT 621.000 259.200 625.200 259.800 ;
        RECT 66.000 258.600 70.200 259.200 ;
        RECT 255.000 258.600 261.000 259.200 ;
        RECT 280.200 258.600 291.000 259.200 ;
        RECT 345.600 258.600 352.200 259.200 ;
        RECT 513.600 258.600 517.200 259.200 ;
        RECT 66.600 258.000 70.200 258.600 ;
        RECT 255.600 258.000 261.000 258.600 ;
        RECT 279.600 258.000 289.200 258.600 ;
        RECT 346.800 258.000 353.400 258.600 ;
        RECT 514.200 258.000 517.200 258.600 ;
        RECT 562.800 258.600 565.800 259.200 ;
        RECT 621.600 258.600 625.800 259.200 ;
        RECT 562.800 258.000 566.400 258.600 ;
        RECT 622.200 258.000 626.400 258.600 ;
        RECT 66.600 257.400 71.400 258.000 ;
        RECT 256.800 257.400 261.600 258.000 ;
        RECT 278.400 257.400 287.400 258.000 ;
        RECT 348.000 257.400 354.600 258.000 ;
        RECT 514.200 257.400 517.800 258.000 ;
        RECT 563.400 257.400 567.000 258.000 ;
        RECT 622.800 257.400 627.000 258.000 ;
        RECT 688.800 257.400 691.800 259.800 ;
        RECT 67.200 256.800 72.600 257.400 ;
        RECT 257.400 256.800 261.600 257.400 ;
        RECT 276.600 256.800 285.600 257.400 ;
        RECT 349.200 256.800 355.200 257.400 ;
        RECT 514.800 256.800 517.800 257.400 ;
        RECT 564.000 256.800 567.000 257.400 ;
        RECT 623.400 256.800 627.600 257.400 ;
        RECT 688.800 256.800 691.200 257.400 ;
        RECT 67.200 256.200 74.400 256.800 ;
        RECT 183.600 256.200 194.400 256.800 ;
        RECT 258.000 256.200 262.200 256.800 ;
        RECT 275.400 256.200 283.800 256.800 ;
        RECT 350.400 256.200 356.400 256.800 ;
        RECT 514.800 256.200 518.400 256.800 ;
        RECT 564.000 256.200 567.600 256.800 ;
        RECT 624.000 256.200 628.200 256.800 ;
        RECT 68.400 255.600 76.800 256.200 ;
        RECT 177.600 255.600 195.600 256.200 ;
        RECT 258.600 255.600 262.800 256.200 ;
        RECT 274.200 255.600 282.000 256.200 ;
        RECT 351.600 255.600 357.000 256.200 ;
        RECT 515.400 255.600 518.400 256.200 ;
        RECT 564.600 255.600 568.200 256.200 ;
        RECT 624.600 255.600 628.800 256.200 ;
        RECT 69.600 255.000 78.600 255.600 ;
        RECT 172.800 255.000 195.600 255.600 ;
        RECT 259.200 255.000 263.400 255.600 ;
        RECT 272.400 255.000 280.200 255.600 ;
        RECT 352.800 255.000 358.200 255.600 ;
        RECT 515.400 255.000 519.000 255.600 ;
        RECT 70.800 254.400 81.600 255.000 ;
        RECT 168.000 254.400 195.600 255.000 ;
        RECT 259.800 254.400 264.000 255.000 ;
        RECT 271.800 254.400 278.400 255.000 ;
        RECT 353.400 254.400 358.800 255.000 ;
        RECT 516.000 254.400 519.000 255.000 ;
        RECT 565.200 255.000 568.200 255.600 ;
        RECT 625.200 255.000 629.400 255.600 ;
        RECT 565.200 254.400 568.800 255.000 ;
        RECT 625.800 254.400 630.000 255.000 ;
        RECT 688.200 254.400 691.200 256.800 ;
        RECT 72.600 253.800 84.000 254.400 ;
        RECT 163.800 253.800 190.800 254.400 ;
        RECT 260.400 253.800 264.600 254.400 ;
        RECT 270.600 253.800 277.200 254.400 ;
        RECT 354.600 253.800 359.400 254.400 ;
        RECT 516.000 253.800 519.600 254.400 ;
        RECT 74.400 253.200 87.000 253.800 ;
        RECT 160.200 253.200 183.000 253.800 ;
        RECT 261.000 253.200 265.200 253.800 ;
        RECT 269.400 253.200 276.000 253.800 ;
        RECT 355.200 253.200 360.000 253.800 ;
        RECT 516.600 253.200 519.600 253.800 ;
        RECT 565.800 253.800 569.400 254.400 ;
        RECT 626.400 253.800 630.600 254.400 ;
        RECT 565.800 253.200 570.000 253.800 ;
        RECT 627.000 253.200 631.200 253.800 ;
        RECT 76.800 252.600 90.000 253.200 ;
        RECT 156.000 252.600 177.000 253.200 ;
        RECT 261.600 252.600 265.800 253.200 ;
        RECT 268.200 252.600 274.800 253.200 ;
        RECT 356.400 252.600 360.600 253.200 ;
        RECT 516.600 252.600 520.200 253.200 ;
        RECT 566.400 252.600 570.000 253.200 ;
        RECT 627.600 252.600 631.800 253.200 ;
        RECT 78.600 252.000 93.000 252.600 ;
        RECT 152.400 252.000 172.200 252.600 ;
        RECT 262.800 252.000 265.800 252.600 ;
        RECT 267.000 252.000 273.600 252.600 ;
        RECT 357.000 252.000 361.200 252.600 ;
        RECT 517.200 252.000 520.200 252.600 ;
        RECT 81.000 251.400 96.600 252.000 ;
        RECT 148.800 251.400 168.000 252.000 ;
        RECT 263.400 251.400 272.400 252.000 ;
        RECT 357.600 251.400 361.200 252.000 ;
        RECT 517.800 251.400 520.800 252.000 ;
        RECT 567.000 251.400 570.600 252.600 ;
        RECT 628.200 252.000 632.400 252.600 ;
        RECT 687.600 252.000 690.600 254.400 ;
        RECT 628.800 251.400 633.000 252.000 ;
        RECT 84.000 250.800 100.800 251.400 ;
        RECT 145.200 250.800 163.800 251.400 ;
        RECT 264.000 250.800 271.200 251.400 ;
        RECT 358.200 250.800 361.800 251.400 ;
        RECT 517.800 250.800 521.400 251.400 ;
        RECT 567.600 250.800 571.200 251.400 ;
        RECT 629.400 250.800 633.600 251.400 ;
        RECT 87.000 250.200 105.600 250.800 ;
        RECT 141.600 250.200 159.600 250.800 ;
        RECT 264.000 250.200 270.000 250.800 ;
        RECT 358.200 250.200 362.400 250.800 ;
        RECT 90.000 249.600 112.800 250.200 ;
        RECT 137.400 249.600 156.000 250.200 ;
        RECT 218.400 249.600 225.000 250.200 ;
        RECT 263.400 249.600 268.800 250.200 ;
        RECT 358.800 249.600 362.400 250.200 ;
        RECT 518.400 250.200 521.400 250.800 ;
        RECT 568.200 250.200 571.200 250.800 ;
        RECT 630.000 250.200 634.200 250.800 ;
        RECT 518.400 249.600 522.000 250.200 ;
        RECT 568.200 249.600 571.800 250.200 ;
        RECT 630.600 249.600 634.800 250.200 ;
        RECT 687.000 249.600 690.000 252.000 ;
        RECT 93.000 249.000 152.400 249.600 ;
        RECT 215.400 249.000 225.000 249.600 ;
        RECT 262.200 249.000 267.600 249.600 ;
        RECT 96.600 248.400 148.800 249.000 ;
        RECT 213.000 248.400 225.000 249.000 ;
        RECT 261.600 248.400 267.000 249.000 ;
        RECT 359.400 248.400 363.000 249.600 ;
        RECT 519.000 249.000 522.000 249.600 ;
        RECT 568.800 249.000 571.800 249.600 ;
        RECT 631.200 249.000 635.400 249.600 ;
        RECT 519.000 248.400 522.600 249.000 ;
        RECT 568.800 248.400 572.400 249.000 ;
        RECT 631.800 248.400 636.000 249.000 ;
        RECT 100.800 247.800 145.200 248.400 ;
        RECT 210.600 247.800 223.800 248.400 ;
        RECT 260.400 247.800 265.800 248.400 ;
        RECT 360.000 247.800 363.000 248.400 ;
        RECT 106.200 247.200 141.600 247.800 ;
        RECT 208.800 247.200 221.400 247.800 ;
        RECT 259.800 247.200 264.600 247.800 ;
        RECT 360.000 247.200 363.600 247.800 ;
        RECT 519.600 247.200 522.600 248.400 ;
        RECT 569.400 247.800 573.000 248.400 ;
        RECT 632.400 247.800 636.000 248.400 ;
        RECT 570.000 247.200 573.000 247.800 ;
        RECT 633.000 247.200 636.600 247.800 ;
        RECT 686.400 247.200 689.400 249.600 ;
        RECT 114.000 246.600 138.000 247.200 ;
        RECT 206.400 246.600 218.400 247.200 ;
        RECT 258.600 246.600 264.000 247.200 ;
        RECT 360.600 246.600 363.600 247.200 ;
        RECT 114.000 246.000 134.400 246.600 ;
        RECT 204.600 246.000 215.400 246.600 ;
        RECT 258.000 246.000 262.800 246.600 ;
        RECT 360.600 246.000 364.200 246.600 ;
        RECT 114.000 245.400 130.800 246.000 ;
        RECT 202.200 245.400 213.000 246.000 ;
        RECT 257.400 245.400 262.200 246.000 ;
        RECT 361.200 245.400 364.200 246.000 ;
        RECT 520.200 246.000 523.200 247.200 ;
        RECT 570.000 246.600 573.600 247.200 ;
        RECT 633.600 246.600 637.200 247.200 ;
        RECT 570.600 246.000 573.600 246.600 ;
        RECT 634.200 246.000 637.800 246.600 ;
        RECT 520.200 245.400 523.800 246.000 ;
        RECT 570.600 245.400 574.200 246.000 ;
        RECT 111.000 244.800 127.800 245.400 ;
        RECT 200.400 244.800 210.600 245.400 ;
        RECT 256.200 244.800 261.000 245.400 ;
        RECT 361.200 244.800 364.800 245.400 ;
        RECT 108.000 244.200 124.200 244.800 ;
        RECT 198.600 244.200 208.800 244.800 ;
        RECT 255.600 244.200 260.400 244.800 ;
        RECT 361.800 244.200 364.800 244.800 ;
        RECT 520.800 244.800 523.800 245.400 ;
        RECT 571.200 244.800 574.200 245.400 ;
        RECT 634.800 245.400 638.400 246.000 ;
        RECT 634.800 244.800 639.000 245.400 ;
        RECT 685.800 244.800 688.800 247.200 ;
        RECT 520.800 244.200 524.400 244.800 ;
        RECT 571.200 244.200 574.800 244.800 ;
        RECT 635.400 244.200 639.600 244.800 ;
        RECT 104.400 243.600 120.600 244.200 ;
        RECT 196.800 243.600 206.400 244.200 ;
        RECT 255.000 243.600 259.800 244.200 ;
        RECT 361.800 243.600 365.400 244.200 ;
        RECT 101.400 243.000 117.600 243.600 ;
        RECT 195.000 243.000 204.600 243.600 ;
        RECT 254.400 243.000 258.600 243.600 ;
        RECT 98.400 242.400 114.000 243.000 ;
        RECT 193.200 242.400 202.800 243.000 ;
        RECT 253.200 242.400 258.000 243.000 ;
        RECT 362.400 242.400 365.400 243.600 ;
        RECT 521.400 243.600 524.400 244.200 ;
        RECT 571.800 243.600 574.800 244.200 ;
        RECT 636.000 243.600 640.200 244.200 ;
        RECT 521.400 243.000 525.000 243.600 ;
        RECT 571.800 243.000 575.400 243.600 ;
        RECT 636.600 243.000 640.800 243.600 ;
        RECT 685.200 243.000 688.200 244.800 ;
        RECT 522.000 242.400 525.000 243.000 ;
        RECT 572.400 242.400 575.400 243.000 ;
        RECT 637.200 242.400 640.800 243.000 ;
        RECT 684.600 242.400 688.200 243.000 ;
        RECT 95.400 241.800 111.000 242.400 ;
        RECT 191.400 241.800 200.400 242.400 ;
        RECT 252.600 241.800 257.400 242.400 ;
        RECT 93.000 241.200 107.400 241.800 ;
        RECT 189.600 241.200 198.600 241.800 ;
        RECT 252.000 241.200 256.800 241.800 ;
        RECT 363.000 241.200 366.000 242.400 ;
        RECT 522.000 241.800 525.600 242.400 ;
        RECT 572.400 241.800 576.000 242.400 ;
        RECT 637.800 241.800 641.400 242.400 ;
        RECT 90.000 240.600 104.400 241.200 ;
        RECT 187.800 240.600 196.800 241.200 ;
        RECT 251.400 240.600 255.600 241.200 ;
        RECT 363.000 240.600 366.600 241.200 ;
        RECT 522.600 240.600 525.600 241.800 ;
        RECT 573.000 241.200 576.000 241.800 ;
        RECT 638.400 241.200 642.000 241.800 ;
        RECT 573.000 240.600 576.600 241.200 ;
        RECT 87.000 240.000 101.400 240.600 ;
        RECT 186.000 240.000 195.000 240.600 ;
        RECT 250.800 240.000 255.000 240.600 ;
        RECT 84.600 239.400 98.400 240.000 ;
        RECT 184.800 239.400 193.200 240.000 ;
        RECT 250.200 239.400 254.400 240.000 ;
        RECT 363.600 239.400 366.600 240.600 ;
        RECT 523.200 239.400 526.200 240.600 ;
        RECT 573.600 240.000 576.600 240.600 ;
        RECT 639.000 240.600 642.600 241.200 ;
        RECT 684.600 240.600 687.600 242.400 ;
        RECT 639.000 240.000 643.200 240.600 ;
        RECT 573.600 239.400 577.200 240.000 ;
        RECT 639.600 239.400 643.800 240.000 ;
        RECT 82.200 238.800 95.400 239.400 ;
        RECT 183.000 238.800 191.400 239.400 ;
        RECT 249.600 238.800 253.800 239.400 ;
        RECT 363.600 238.800 367.200 239.400 ;
        RECT 523.200 238.800 526.800 239.400 ;
        RECT 79.800 238.200 93.000 238.800 ;
        RECT 181.200 238.200 190.200 238.800 ;
        RECT 249.000 238.200 253.200 238.800 ;
        RECT 77.400 237.600 90.000 238.200 ;
        RECT 180.000 237.600 188.400 238.200 ;
        RECT 248.400 237.600 252.600 238.200 ;
        RECT 75.000 237.000 87.600 237.600 ;
        RECT 178.200 237.000 186.600 237.600 ;
        RECT 247.800 237.000 252.000 237.600 ;
        RECT 364.200 237.000 367.200 238.800 ;
        RECT 523.800 238.200 526.800 238.800 ;
        RECT 574.200 238.800 577.200 239.400 ;
        RECT 640.200 238.800 644.400 239.400 ;
        RECT 684.000 238.800 687.000 240.600 ;
        RECT 574.200 238.200 577.800 238.800 ;
        RECT 640.800 238.200 644.400 238.800 ;
        RECT 683.400 238.200 687.000 238.800 ;
        RECT 523.800 237.600 527.400 238.200 ;
        RECT 73.200 236.400 84.600 237.000 ;
        RECT 176.400 236.400 184.800 237.000 ;
        RECT 247.200 236.400 251.400 237.000 ;
        RECT 70.800 235.800 82.200 236.400 ;
        RECT 175.200 235.800 183.600 236.400 ;
        RECT 246.600 235.800 250.800 236.400 ;
        RECT 69.000 235.200 79.800 235.800 ;
        RECT 173.400 235.200 181.800 235.800 ;
        RECT 246.000 235.200 250.200 235.800 ;
        RECT 364.800 235.200 367.800 237.000 ;
        RECT 524.400 236.400 527.400 237.600 ;
        RECT 574.800 237.600 577.800 238.200 ;
        RECT 641.400 237.600 645.000 238.200 ;
        RECT 574.800 237.000 578.400 237.600 ;
        RECT 642.000 237.000 645.600 237.600 ;
        RECT 683.400 237.000 686.400 238.200 ;
        RECT 575.400 236.400 578.400 237.000 ;
        RECT 642.600 236.400 646.200 237.000 ;
        RECT 682.800 236.400 686.400 237.000 ;
        RECT 525.000 235.200 528.000 236.400 ;
        RECT 575.400 235.800 579.000 236.400 ;
        RECT 642.600 235.800 646.800 236.400 ;
        RECT 66.600 234.600 77.400 235.200 ;
        RECT 172.200 234.600 180.000 235.200 ;
        RECT 245.400 234.600 249.600 235.200 ;
        RECT 64.800 234.000 75.000 234.600 ;
        RECT 170.400 234.000 178.800 234.600 ;
        RECT 244.800 234.000 249.000 234.600 ;
        RECT 63.000 233.400 73.200 234.000 ;
        RECT 169.200 233.400 177.000 234.000 ;
        RECT 244.200 233.400 248.400 234.000 ;
        RECT 61.200 232.800 70.800 233.400 ;
        RECT 167.400 232.800 175.800 233.400 ;
        RECT 243.600 232.800 247.800 233.400 ;
        RECT 365.400 232.800 368.400 235.200 ;
        RECT 525.000 234.600 528.600 235.200 ;
        RECT 576.000 234.600 579.000 235.800 ;
        RECT 643.200 235.200 647.400 235.800 ;
        RECT 643.800 234.600 647.400 235.200 ;
        RECT 682.800 234.600 685.800 236.400 ;
        RECT 525.600 233.400 528.600 234.600 ;
        RECT 576.600 233.400 579.600 234.600 ;
        RECT 644.400 234.000 648.000 234.600 ;
        RECT 645.000 233.400 648.600 234.000 ;
        RECT 525.600 232.800 529.200 233.400 ;
        RECT 576.600 232.800 580.200 233.400 ;
        RECT 645.000 232.800 649.200 233.400 ;
        RECT 682.200 232.800 685.200 234.600 ;
        RECT 59.400 232.200 69.000 232.800 ;
        RECT 166.200 232.200 174.000 232.800 ;
        RECT 243.600 232.200 247.200 232.800 ;
        RECT 58.200 231.600 67.200 232.200 ;
        RECT 165.000 231.600 172.800 232.200 ;
        RECT 243.000 231.600 246.600 232.200 ;
        RECT 57.000 231.000 65.400 231.600 ;
        RECT 163.200 231.000 171.000 231.600 ;
        RECT 242.400 231.000 246.000 231.600 ;
        RECT 55.800 230.400 63.600 231.000 ;
        RECT 162.000 230.400 169.800 231.000 ;
        RECT 241.800 230.400 245.400 231.000 ;
        RECT 366.000 230.400 369.000 232.800 ;
        RECT 526.200 231.600 529.200 232.800 ;
        RECT 577.200 232.200 580.200 232.800 ;
        RECT 645.600 232.200 649.800 232.800 ;
        RECT 577.200 231.600 580.800 232.200 ;
        RECT 646.200 231.600 649.800 232.200 ;
        RECT 54.600 229.800 61.800 230.400 ;
        RECT 160.200 229.800 168.000 230.400 ;
        RECT 241.200 229.800 245.400 230.400 ;
        RECT 54.000 229.200 60.000 229.800 ;
        RECT 159.000 229.200 166.800 229.800 ;
        RECT 240.600 229.200 244.800 229.800 ;
        RECT 53.400 228.600 58.800 229.200 ;
        RECT 157.800 228.600 165.000 229.200 ;
        RECT 240.600 228.600 244.200 229.200 ;
        RECT 52.800 228.000 57.600 228.600 ;
        RECT 156.000 228.000 163.800 228.600 ;
        RECT 240.000 228.000 243.600 228.600 ;
        RECT 366.600 228.000 369.600 230.400 ;
        RECT 526.800 229.800 529.800 231.600 ;
        RECT 577.800 230.400 580.800 231.600 ;
        RECT 646.800 231.000 650.400 231.600 ;
        RECT 681.600 231.000 684.600 232.800 ;
        RECT 647.400 230.400 651.000 231.000 ;
        RECT 527.400 228.000 530.400 229.800 ;
        RECT 578.400 229.200 581.400 230.400 ;
        RECT 648.000 229.800 651.600 230.400 ;
        RECT 681.000 229.800 684.000 231.000 ;
        RECT 648.000 229.200 652.200 229.800 ;
        RECT 578.400 228.600 582.000 229.200 ;
        RECT 648.600 228.600 652.200 229.200 ;
        RECT 680.400 229.200 684.000 229.800 ;
        RECT 52.200 227.400 56.400 228.000 ;
        RECT 154.800 227.400 162.000 228.000 ;
        RECT 239.400 227.400 243.000 228.000 ;
        RECT 51.600 226.800 55.800 227.400 ;
        RECT 153.600 226.800 160.800 227.400 ;
        RECT 51.600 225.600 55.200 226.800 ;
        RECT 151.800 226.200 159.600 226.800 ;
        RECT 238.800 226.200 242.400 227.400 ;
        RECT 150.600 225.600 157.800 226.200 ;
        RECT 238.200 225.600 241.800 226.200 ;
        RECT 51.600 225.000 55.800 225.600 ;
        RECT 149.400 225.000 156.600 225.600 ;
        RECT 237.600 225.000 241.200 225.600 ;
        RECT 367.200 225.000 370.200 228.000 ;
        RECT 528.000 226.200 531.000 228.000 ;
        RECT 579.000 227.400 582.000 228.600 ;
        RECT 649.200 228.000 652.800 228.600 ;
        RECT 680.400 228.000 683.400 229.200 ;
        RECT 649.800 227.400 653.400 228.000 ;
        RECT 679.800 227.400 683.400 228.000 ;
        RECT 579.000 226.800 582.600 227.400 ;
        RECT 52.200 224.400 57.600 225.000 ;
        RECT 148.200 224.400 154.800 225.000 ;
        RECT 52.200 223.800 59.400 224.400 ;
        RECT 146.400 223.800 153.000 224.400 ;
        RECT 237.000 223.800 240.600 225.000 ;
        RECT 53.400 223.200 61.200 223.800 ;
        RECT 145.200 223.200 151.800 223.800 ;
        RECT 236.400 223.200 240.000 223.800 ;
        RECT 54.000 222.600 63.600 223.200 ;
        RECT 144.000 222.600 150.600 223.200 ;
        RECT 55.200 222.000 66.600 222.600 ;
        RECT 142.800 222.000 149.400 222.600 ;
        RECT 235.800 222.000 239.400 223.200 ;
        RECT 57.000 221.400 70.200 222.000 ;
        RECT 141.600 221.400 148.200 222.000 ;
        RECT 234.600 221.400 238.800 222.000 ;
        RECT 58.800 220.800 73.800 221.400 ;
        RECT 139.800 220.800 147.600 221.400 ;
        RECT 233.400 220.800 238.200 221.400 ;
        RECT 61.200 220.200 78.600 220.800 ;
        RECT 135.600 220.200 146.400 220.800 ;
        RECT 231.600 220.200 238.200 220.800 ;
        RECT 334.200 220.200 334.800 222.000 ;
        RECT 367.800 221.400 370.800 225.000 ;
        RECT 528.600 223.800 531.600 226.200 ;
        RECT 579.600 225.600 582.600 226.800 ;
        RECT 650.400 226.800 654.000 227.400 ;
        RECT 650.400 226.200 654.600 226.800 ;
        RECT 679.800 226.200 682.800 227.400 ;
        RECT 651.000 225.600 654.600 226.200 ;
        RECT 679.200 225.600 682.800 226.200 ;
        RECT 580.200 223.800 583.200 225.600 ;
        RECT 651.600 225.000 655.200 225.600 ;
        RECT 652.200 224.400 655.800 225.000 ;
        RECT 679.200 224.400 682.200 225.600 ;
        RECT 652.800 223.800 656.400 224.400 ;
        RECT 529.200 222.000 532.200 223.800 ;
        RECT 580.800 222.000 583.800 223.800 ;
        RECT 652.800 223.200 657.000 223.800 ;
        RECT 678.600 223.200 681.600 224.400 ;
        RECT 653.400 222.600 657.000 223.200 ;
        RECT 678.000 222.600 681.600 223.200 ;
        RECT 654.000 222.000 657.600 222.600 ;
        RECT 529.200 221.400 532.800 222.000 ;
        RECT 63.600 219.600 84.000 220.200 ;
        RECT 128.400 219.600 144.600 220.200 ;
        RECT 230.400 219.600 237.600 220.200 ;
        RECT 334.200 219.600 335.400 220.200 ;
        RECT 66.600 219.000 91.200 219.600 ;
        RECT 120.000 219.000 143.400 219.600 ;
        RECT 228.600 219.000 237.000 219.600 ;
        RECT 70.200 218.400 141.600 219.000 ;
        RECT 227.400 218.400 237.000 219.000 ;
        RECT 74.400 217.800 140.400 218.400 ;
        RECT 225.600 217.800 236.400 218.400 ;
        RECT 78.600 217.200 129.600 217.800 ;
        RECT 130.800 217.200 139.200 217.800 ;
        RECT 224.400 217.200 235.800 217.800 ;
        RECT 84.600 216.600 124.800 217.200 ;
        RECT 130.800 216.600 138.000 217.200 ;
        RECT 222.600 216.600 229.800 217.200 ;
        RECT 232.200 216.600 235.800 217.200 ;
        RECT 333.600 216.600 335.400 219.600 ;
        RECT 368.400 217.800 371.400 221.400 ;
        RECT 529.800 219.000 532.800 221.400 ;
        RECT 581.400 220.200 584.400 222.000 ;
        RECT 654.600 221.400 658.200 222.000 ;
        RECT 678.000 221.400 681.000 222.600 ;
        RECT 655.200 220.800 658.800 221.400 ;
        RECT 677.400 220.800 681.000 221.400 ;
        RECT 655.200 220.200 659.400 220.800 ;
        RECT 581.400 219.600 585.000 220.200 ;
        RECT 655.800 219.600 659.400 220.200 ;
        RECT 677.400 219.600 680.400 220.800 ;
        RECT 91.800 216.000 118.200 216.600 ;
        RECT 129.600 216.000 136.800 216.600 ;
        RECT 220.800 216.000 228.600 216.600 ;
        RECT 232.200 216.000 235.200 216.600 ;
        RECT 128.400 215.400 135.600 216.000 ;
        RECT 219.600 215.400 226.800 216.000 ;
        RECT 231.600 215.400 235.200 216.000 ;
        RECT 127.200 214.800 134.400 215.400 ;
        RECT 217.800 214.800 225.600 215.400 ;
        RECT 231.600 214.800 234.600 215.400 ;
        RECT 126.000 214.200 132.600 214.800 ;
        RECT 216.000 214.200 223.800 214.800 ;
        RECT 231.000 214.200 234.600 214.800 ;
        RECT 124.800 213.600 131.400 214.200 ;
        RECT 214.800 213.600 222.600 214.200 ;
        RECT 231.000 213.600 234.000 214.200 ;
        RECT 123.600 213.000 130.200 213.600 ;
        RECT 213.000 213.000 220.800 213.600 ;
        RECT 230.400 213.000 234.000 213.600 ;
        RECT 333.000 213.000 335.400 216.600 ;
        RECT 369.000 214.200 372.000 217.800 ;
        RECT 530.400 216.600 533.400 219.000 ;
        RECT 582.000 217.800 585.000 219.600 ;
        RECT 656.400 219.000 660.000 219.600 ;
        RECT 657.000 218.400 660.600 219.000 ;
        RECT 676.800 218.400 679.800 219.600 ;
        RECT 657.600 217.800 661.200 218.400 ;
        RECT 676.200 217.800 679.800 218.400 ;
        RECT 122.400 212.400 129.000 213.000 ;
        RECT 211.200 212.400 219.600 213.000 ;
        RECT 230.400 212.400 233.400 213.000 ;
        RECT 121.200 211.800 127.800 212.400 ;
        RECT 209.400 211.800 217.800 212.400 ;
        RECT 229.800 211.800 233.400 212.400 ;
        RECT 332.400 212.400 335.400 213.000 ;
        RECT 369.600 213.600 372.000 214.200 ;
        RECT 120.000 211.200 126.600 211.800 ;
        RECT 207.600 211.200 216.600 211.800 ;
        RECT 229.800 211.200 232.800 211.800 ;
        RECT 118.800 210.600 125.400 211.200 ;
        RECT 205.800 210.600 214.800 211.200 ;
        RECT 229.200 210.600 232.800 211.200 ;
        RECT 117.600 210.000 124.200 210.600 ;
        RECT 204.600 210.000 213.000 210.600 ;
        RECT 229.200 210.000 232.200 210.600 ;
        RECT 116.400 209.400 123.000 210.000 ;
        RECT 202.800 209.400 211.200 210.000 ;
        RECT 228.600 209.400 232.200 210.000 ;
        RECT 332.400 209.400 334.800 212.400 ;
        RECT 369.600 209.400 372.600 213.600 ;
        RECT 531.000 213.000 534.000 216.600 ;
        RECT 582.600 215.400 585.600 217.800 ;
        RECT 657.600 217.200 661.800 217.800 ;
        RECT 676.200 217.200 679.200 217.800 ;
        RECT 658.200 216.600 661.800 217.200 ;
        RECT 675.600 216.600 679.200 217.200 ;
        RECT 658.800 216.000 662.400 216.600 ;
        RECT 659.400 215.400 663.000 216.000 ;
        RECT 675.600 215.400 678.600 216.600 ;
        RECT 583.200 213.000 586.200 215.400 ;
        RECT 660.000 214.800 663.600 215.400 ;
        RECT 675.000 214.800 678.600 215.400 ;
        RECT 660.000 214.200 664.200 214.800 ;
        RECT 675.000 214.200 678.000 214.800 ;
        RECT 660.600 213.600 664.200 214.200 ;
        RECT 674.400 213.600 678.000 214.200 ;
        RECT 661.200 213.000 664.800 213.600 ;
        RECT 674.400 213.000 677.400 213.600 ;
        RECT 115.200 208.800 121.800 209.400 ;
        RECT 200.400 208.800 210.000 209.400 ;
        RECT 228.600 208.800 231.600 209.400 ;
        RECT 114.000 208.200 120.600 208.800 ;
        RECT 198.600 208.200 208.200 208.800 ;
        RECT 228.000 208.200 231.600 208.800 ;
        RECT 113.400 207.600 119.400 208.200 ;
        RECT 196.800 207.600 206.400 208.200 ;
        RECT 228.000 207.600 231.000 208.200 ;
        RECT 112.200 207.000 118.200 207.600 ;
        RECT 195.000 207.000 204.600 207.600 ;
        RECT 227.400 207.000 231.000 207.600 ;
        RECT 111.000 206.400 117.000 207.000 ;
        RECT 193.200 206.400 202.800 207.000 ;
        RECT 109.800 205.800 115.800 206.400 ;
        RECT 190.800 205.800 201.000 206.400 ;
        RECT 227.400 205.800 230.400 207.000 ;
        RECT 331.800 206.400 334.800 209.400 ;
        RECT 370.200 208.800 372.600 209.400 ;
        RECT 531.600 208.800 534.600 213.000 ;
        RECT 583.800 210.000 586.800 213.000 ;
        RECT 661.800 212.400 665.400 213.000 ;
        RECT 673.800 212.400 677.400 213.000 ;
        RECT 662.400 211.800 666.000 212.400 ;
        RECT 662.400 211.200 666.600 211.800 ;
        RECT 673.800 211.200 676.800 212.400 ;
        RECT 663.000 210.600 666.600 211.200 ;
        RECT 663.600 210.000 667.200 210.600 ;
        RECT 673.200 210.000 676.200 211.200 ;
        RECT 331.800 205.800 334.200 206.400 ;
        RECT 108.600 205.200 114.600 205.800 ;
        RECT 189.000 205.200 199.200 205.800 ;
        RECT 107.400 204.600 114.000 205.200 ;
        RECT 186.600 204.600 196.800 205.200 ;
        RECT 226.800 204.600 229.800 205.800 ;
        RECT 106.800 204.000 112.800 204.600 ;
        RECT 184.800 204.000 195.000 204.600 ;
        RECT 226.200 204.000 229.800 204.600 ;
        RECT 105.600 203.400 111.600 204.000 ;
        RECT 182.400 203.400 193.200 204.000 ;
        RECT 104.400 202.800 110.400 203.400 ;
        RECT 180.000 202.800 191.400 203.400 ;
        RECT 226.200 202.800 229.200 204.000 ;
        RECT 331.200 202.800 334.200 205.800 ;
        RECT 370.200 203.400 373.200 208.800 ;
        RECT 531.600 208.200 535.200 208.800 ;
        RECT 532.200 205.800 535.200 208.200 ;
        RECT 584.400 207.000 587.400 210.000 ;
        RECT 664.200 209.400 667.800 210.000 ;
        RECT 672.600 209.400 676.200 210.000 ;
        RECT 664.200 208.800 668.400 209.400 ;
        RECT 672.600 208.800 675.600 209.400 ;
        RECT 664.800 208.200 668.400 208.800 ;
        RECT 672.000 208.200 675.600 208.800 ;
        RECT 665.400 207.600 669.000 208.200 ;
        RECT 672.000 207.600 675.000 208.200 ;
        RECT 666.000 207.000 669.600 207.600 ;
        RECT 671.400 207.000 675.000 207.600 ;
        RECT 532.200 204.000 534.600 205.800 ;
        RECT 103.200 202.200 109.200 202.800 ;
        RECT 177.600 202.200 189.000 202.800 ;
        RECT 225.600 202.200 229.200 202.800 ;
        RECT 102.600 201.600 108.000 202.200 ;
        RECT 175.800 201.600 187.200 202.200 ;
        RECT 101.400 201.000 107.400 201.600 ;
        RECT 172.800 201.000 184.800 201.600 ;
        RECT 225.600 201.000 228.600 202.200 ;
        RECT 100.200 200.400 106.200 201.000 ;
        RECT 170.400 200.400 184.800 201.000 ;
        RECT 99.600 199.800 105.000 200.400 ;
        RECT 168.000 199.800 180.000 200.400 ;
        RECT 98.400 199.200 103.800 199.800 ;
        RECT 165.000 199.200 178.200 199.800 ;
        RECT 97.800 198.600 103.200 199.200 ;
        RECT 162.600 198.600 175.800 199.200 ;
        RECT 96.600 198.000 102.000 198.600 ;
        RECT 159.600 198.000 173.400 198.600 ;
        RECT 96.000 197.400 100.800 198.000 ;
        RECT 156.600 197.400 170.400 198.000 ;
        RECT 94.800 196.800 100.200 197.400 ;
        RECT 153.600 196.800 168.000 197.400 ;
        RECT 94.200 196.200 99.000 196.800 ;
        RECT 150.000 196.200 165.000 196.800 ;
        RECT 93.600 195.600 98.400 196.200 ;
        RECT 147.000 195.600 162.600 196.200 ;
        RECT 93.000 195.000 97.200 195.600 ;
        RECT 142.800 195.000 159.600 195.600 ;
        RECT 92.400 194.400 96.600 195.000 ;
        RECT 139.200 194.400 156.600 195.000 ;
        RECT 92.400 193.800 96.000 194.400 ;
        RECT 135.000 193.800 153.600 194.400 ;
        RECT 91.800 192.600 95.400 193.800 ;
        RECT 129.600 193.200 150.000 193.800 ;
        RECT 124.200 192.600 146.400 193.200 ;
        RECT 91.800 192.000 97.200 192.600 ;
        RECT 117.600 192.000 142.800 192.600 ;
        RECT 92.400 191.400 138.600 192.000 ;
        RECT 92.400 190.800 134.400 191.400 ;
        RECT 93.600 190.200 129.600 190.800 ;
        RECT 94.800 189.600 123.600 190.200 ;
        RECT 97.800 189.000 116.400 189.600 ;
        RECT 181.800 180.600 184.800 200.400 ;
        RECT 225.000 199.200 228.000 201.000 ;
        RECT 330.600 199.800 333.600 202.800 ;
        RECT 370.200 201.000 373.800 203.400 ;
        RECT 224.400 196.800 227.400 199.200 ;
        RECT 330.000 197.400 333.000 199.800 ;
        RECT 370.800 199.200 373.800 201.000 ;
        RECT 401.400 199.800 415.200 200.400 ;
        RECT 392.400 199.200 416.400 199.800 ;
        RECT 370.800 198.600 378.600 199.200 ;
        RECT 385.200 198.600 417.000 199.200 ;
        RECT 370.800 198.000 417.600 198.600 ;
        RECT 370.800 197.400 418.200 198.000 ;
        RECT 329.400 196.800 333.000 197.400 ;
        RECT 371.400 196.800 400.200 197.400 ;
        RECT 414.600 196.800 419.400 197.400 ;
        RECT 531.600 196.800 534.600 204.000 ;
        RECT 585.000 202.800 588.000 207.000 ;
        RECT 666.600 206.400 670.200 207.000 ;
        RECT 671.400 206.400 674.400 207.000 ;
        RECT 667.200 205.800 674.400 206.400 ;
        RECT 667.200 205.200 673.800 205.800 ;
        RECT 667.800 204.600 673.800 205.200 ;
        RECT 668.400 204.000 673.200 204.600 ;
        RECT 669.600 203.400 673.200 204.000 ;
        RECT 670.200 202.800 672.600 203.400 ;
        RECT 585.600 196.800 588.600 202.800 ;
        RECT 670.800 202.200 672.000 202.800 ;
        RECT 223.800 194.400 226.800 196.800 ;
        RECT 329.400 195.600 333.600 196.800 ;
        RECT 371.400 196.200 373.800 196.800 ;
        RECT 375.000 196.200 391.800 196.800 ;
        RECT 415.200 196.200 421.200 196.800 ;
        RECT 531.600 196.200 534.000 196.800 ;
        RECT 372.000 195.600 373.200 196.200 ;
        RECT 378.600 195.600 384.000 196.200 ;
        RECT 415.800 195.600 421.800 196.200 ;
        RECT 329.400 195.000 334.200 195.600 ;
        RECT 416.400 195.000 423.000 195.600 ;
        RECT 328.800 194.400 334.800 195.000 ;
        RECT 416.400 194.400 423.600 195.000 ;
        RECT 223.800 193.800 226.200 194.400 ;
        RECT 223.200 192.000 226.200 193.800 ;
        RECT 328.800 193.800 335.400 194.400 ;
        RECT 405.000 193.800 411.600 194.400 ;
        RECT 415.800 193.800 424.800 194.400 ;
        RECT 328.800 193.200 336.000 193.800 ;
        RECT 328.800 192.600 336.600 193.200 ;
        RECT 403.800 192.600 418.800 193.800 ;
        RECT 420.600 193.200 425.400 193.800 ;
        RECT 420.600 192.600 426.000 193.200 ;
        RECT 223.800 190.800 225.600 192.000 ;
        RECT 328.200 190.800 331.200 192.600 ;
        RECT 333.000 192.000 337.200 192.600 ;
        RECT 404.400 192.000 426.600 192.600 ;
        RECT 531.000 192.000 534.000 196.200 ;
        RECT 586.200 195.600 588.600 196.800 ;
        RECT 333.600 191.400 337.800 192.000 ;
        RECT 405.600 191.400 426.600 192.000 ;
        RECT 334.200 190.800 338.400 191.400 ;
        RECT 411.000 190.800 427.200 191.400 ;
        RECT 327.600 190.200 331.200 190.800 ;
        RECT 334.800 190.200 339.600 190.800 ;
        RECT 414.000 190.200 430.200 190.800 ;
        RECT 327.600 189.000 330.600 190.200 ;
        RECT 335.400 189.600 340.200 190.200 ;
        RECT 418.200 189.600 432.600 190.200 ;
        RECT 336.000 189.000 340.800 189.600 ;
        RECT 421.200 189.000 435.000 189.600 ;
        RECT 530.400 189.000 533.400 192.000 ;
        RECT 327.000 188.400 330.600 189.000 ;
        RECT 337.200 188.400 342.000 189.000 ;
        RECT 423.600 188.400 437.400 189.000 ;
        RECT 327.000 186.600 330.000 188.400 ;
        RECT 337.800 187.800 342.600 188.400 ;
        RECT 426.600 187.800 439.800 188.400 ;
        RECT 338.400 187.200 343.800 187.800 ;
        RECT 429.000 187.200 442.200 187.800 ;
        RECT 339.000 186.600 344.400 187.200 ;
        RECT 432.000 186.600 444.000 187.200 ;
        RECT 326.400 185.400 329.400 186.600 ;
        RECT 340.200 186.000 345.600 186.600 ;
        RECT 434.400 186.000 445.800 186.600 ;
        RECT 529.800 186.000 532.800 189.000 ;
        RECT 586.200 187.200 589.200 195.600 ;
        RECT 658.200 187.800 661.200 188.400 ;
        RECT 340.800 185.400 346.800 186.000 ;
        RECT 437.400 185.400 448.200 186.000 ;
        RECT 325.800 184.800 329.400 185.400 ;
        RECT 342.000 184.800 347.400 185.400 ;
        RECT 439.800 184.800 449.400 185.400 ;
        RECT 325.800 183.600 328.800 184.800 ;
        RECT 342.600 184.200 348.600 184.800 ;
        RECT 442.200 184.200 451.200 184.800 ;
        RECT 343.800 183.600 349.800 184.200 ;
        RECT 444.000 183.600 453.000 184.200 ;
        RECT 529.200 183.600 532.200 186.000 ;
        RECT 586.200 185.400 588.600 187.200 ;
        RECT 657.600 186.600 661.800 187.800 ;
        RECT 325.200 183.000 328.800 183.600 ;
        RECT 345.000 183.000 351.000 183.600 ;
        RECT 445.800 183.000 454.800 183.600 ;
        RECT 325.200 181.800 328.200 183.000 ;
        RECT 346.200 182.400 352.200 183.000 ;
        RECT 447.600 182.400 456.600 183.000 ;
        RECT 347.400 181.800 353.400 182.400 ;
        RECT 449.400 181.800 457.800 182.400 ;
        RECT 528.600 181.800 531.600 183.600 ;
        RECT 324.600 180.600 327.600 181.800 ;
        RECT 348.600 181.200 356.400 181.800 ;
        RECT 450.600 181.200 459.000 181.800 ;
        RECT 349.800 180.600 357.000 181.200 ;
        RECT 452.400 180.600 460.200 181.200 ;
        RECT 182.400 178.800 184.800 180.600 ;
        RECT 324.000 180.000 327.600 180.600 ;
        RECT 352.200 180.000 357.000 180.600 ;
        RECT 454.200 180.000 461.400 180.600 ;
        RECT 528.000 180.000 531.000 181.800 ;
        RECT 324.000 178.800 327.000 180.000 ;
        RECT 182.400 171.000 185.400 178.800 ;
        RECT 323.400 177.600 326.400 178.800 ;
        RECT 354.600 177.600 357.600 180.000 ;
        RECT 455.400 179.400 462.000 180.000 ;
        RECT 527.400 179.400 531.000 180.000 ;
        RECT 585.600 180.000 588.600 185.400 ;
        RECT 657.000 186.000 661.800 186.600 ;
        RECT 657.000 184.800 661.200 186.000 ;
        RECT 657.000 183.600 660.600 184.800 ;
        RECT 657.000 182.400 661.200 183.600 ;
        RECT 657.000 181.800 661.800 182.400 ;
        RECT 657.000 181.200 662.400 181.800 ;
        RECT 657.600 180.600 663.600 181.200 ;
        RECT 658.200 180.000 664.800 180.600 ;
        RECT 585.600 179.400 588.000 180.000 ;
        RECT 653.400 179.400 656.400 180.000 ;
        RECT 658.200 179.400 666.000 180.000 ;
        RECT 457.200 178.800 463.200 179.400 ;
        RECT 458.400 178.200 463.800 178.800 ;
        RECT 527.400 178.200 530.400 179.400 ;
        RECT 459.600 177.600 464.400 178.200 ;
        RECT 526.800 177.600 530.400 178.200 ;
        RECT 322.800 177.000 326.400 177.600 ;
        RECT 322.800 176.400 325.800 177.000 ;
        RECT 322.200 175.800 325.800 176.400 ;
        RECT 322.200 174.600 325.200 175.800 ;
        RECT 355.200 174.600 358.200 177.600 ;
        RECT 460.800 177.000 465.000 177.600 ;
        RECT 461.400 176.400 465.600 177.000 ;
        RECT 526.800 176.400 529.800 177.600 ;
        RECT 462.000 175.800 466.200 176.400 ;
        RECT 462.600 175.200 466.800 175.800 ;
        RECT 526.200 175.200 529.200 176.400 ;
        RECT 585.000 175.800 588.000 179.400 ;
        RECT 652.800 178.200 657.000 179.400 ;
        RECT 658.800 178.800 666.000 179.400 ;
        RECT 659.400 178.200 666.600 178.800 ;
        RECT 463.200 174.600 467.400 175.200 ;
        RECT 525.600 174.600 529.200 175.200 ;
        RECT 584.400 175.200 588.000 175.800 ;
        RECT 652.200 177.000 657.000 178.200 ;
        RECT 660.600 177.600 666.600 178.200 ;
        RECT 661.200 177.000 666.000 177.600 ;
        RECT 652.200 175.800 656.400 177.000 ;
        RECT 663.000 176.400 665.400 177.000 ;
        RECT 652.200 175.200 657.000 175.800 ;
        RECT 321.600 173.400 324.600 174.600 ;
        RECT 321.000 172.800 324.600 173.400 ;
        RECT 321.000 172.200 324.000 172.800 ;
        RECT 355.800 172.200 358.800 174.600 ;
        RECT 463.800 174.000 468.000 174.600 ;
        RECT 464.400 173.400 468.600 174.000 ;
        RECT 525.600 173.400 528.600 174.600 ;
        RECT 465.000 172.800 468.600 173.400 ;
        RECT 465.600 172.200 469.200 172.800 ;
        RECT 525.000 172.200 528.000 173.400 ;
        RECT 584.400 172.800 587.400 175.200 ;
        RECT 652.800 174.600 657.600 175.200 ;
        RECT 652.800 174.000 658.200 174.600 ;
        RECT 652.800 173.400 659.400 174.000 ;
        RECT 653.400 172.800 660.000 173.400 ;
        RECT 320.400 171.600 324.000 172.200 ;
        RECT 320.400 171.000 323.400 171.600 ;
        RECT 183.000 169.800 185.400 171.000 ;
        RECT 319.800 170.400 323.400 171.000 ;
        RECT 356.400 170.400 359.400 172.200 ;
        RECT 466.200 171.000 469.800 172.200 ;
        RECT 524.400 171.600 528.000 172.200 ;
        RECT 583.800 172.200 587.400 172.800 ;
        RECT 654.000 172.200 660.600 172.800 ;
        RECT 524.400 171.000 527.400 171.600 ;
        RECT 466.800 170.400 470.400 171.000 ;
        RECT 319.800 169.800 322.800 170.400 ;
        RECT 183.000 164.400 186.000 169.800 ;
        RECT 319.200 169.200 322.800 169.800 ;
        RECT 357.000 169.200 360.000 170.400 ;
        RECT 467.400 169.800 470.400 170.400 ;
        RECT 523.800 170.400 527.400 171.000 ;
        RECT 583.800 170.400 586.800 172.200 ;
        RECT 654.600 171.600 661.200 172.200 ;
        RECT 655.200 171.000 661.800 171.600 ;
        RECT 656.400 170.400 661.800 171.000 ;
        RECT 523.800 169.800 526.800 170.400 ;
        RECT 467.400 169.200 471.000 169.800 ;
        RECT 318.600 168.600 322.200 169.200 ;
        RECT 357.000 168.600 360.600 169.200 ;
        RECT 318.600 168.000 321.600 168.600 ;
        RECT 318.000 167.400 321.600 168.000 ;
        RECT 357.600 168.000 360.600 168.600 ;
        RECT 468.000 168.000 471.000 169.200 ;
        RECT 523.200 169.200 526.800 169.800 ;
        RECT 583.200 169.800 586.800 170.400 ;
        RECT 657.000 169.800 661.800 170.400 ;
        RECT 523.200 168.600 526.200 169.200 ;
        RECT 583.200 168.600 586.200 169.800 ;
        RECT 657.600 169.200 661.200 169.800 ;
        RECT 649.800 168.600 652.800 169.200 ;
        RECT 657.600 168.600 659.400 169.200 ;
        RECT 522.600 168.000 526.200 168.600 ;
        RECT 582.600 168.000 586.200 168.600 ;
        RECT 649.200 168.000 653.400 168.600 ;
        RECT 657.000 168.000 659.400 168.600 ;
        RECT 357.600 167.400 361.200 168.000 ;
        RECT 465.600 167.400 471.600 168.000 ;
        RECT 522.600 167.400 525.600 168.000 ;
        RECT 318.000 166.800 321.000 167.400 ;
        RECT 317.400 166.200 321.000 166.800 ;
        RECT 358.200 166.800 361.200 167.400 ;
        RECT 453.600 166.800 456.600 167.400 ;
        RECT 358.200 166.200 361.800 166.800 ;
        RECT 317.400 165.600 320.400 166.200 ;
        RECT 316.800 165.000 320.400 165.600 ;
        RECT 358.800 165.600 361.800 166.200 ;
        RECT 453.600 166.200 459.000 166.800 ;
        RECT 464.400 166.200 471.600 167.400 ;
        RECT 522.000 166.800 525.600 167.400 ;
        RECT 453.600 165.600 460.800 166.200 ;
        RECT 358.800 165.000 362.400 165.600 ;
        RECT 453.600 165.000 462.000 165.600 ;
        RECT 463.800 165.000 471.600 166.200 ;
        RECT 521.400 166.200 525.000 166.800 ;
        RECT 582.600 166.200 585.600 168.000 ;
        RECT 521.400 165.600 524.400 166.200 ;
        RECT 183.600 163.800 186.000 164.400 ;
        RECT 316.200 163.800 319.800 165.000 ;
        RECT 359.400 164.400 363.000 165.000 ;
        RECT 454.800 164.400 471.600 165.000 ;
        RECT 520.800 165.000 524.400 165.600 ;
        RECT 582.000 165.600 585.600 166.200 ;
        RECT 648.600 167.400 654.000 168.000 ;
        RECT 648.600 166.200 654.600 167.400 ;
        RECT 656.400 166.800 660.000 168.000 ;
        RECT 582.000 165.000 585.000 165.600 ;
        RECT 520.800 164.400 523.800 165.000 ;
        RECT 359.400 163.800 363.600 164.400 ;
        RECT 456.600 163.800 466.800 164.400 ;
        RECT 468.000 163.800 471.600 164.400 ;
        RECT 520.200 163.800 523.800 164.400 ;
        RECT 581.400 163.800 585.000 165.000 ;
        RECT 648.600 164.400 655.200 166.200 ;
        RECT 656.400 164.400 660.600 166.800 ;
        RECT 183.600 159.000 186.600 163.800 ;
        RECT 315.600 163.200 320.400 163.800 ;
        RECT 360.000 163.200 364.200 163.800 ;
        RECT 459.000 163.200 466.800 163.800 ;
        RECT 468.600 163.200 472.200 163.800 ;
        RECT 519.600 163.200 523.200 163.800 ;
        RECT 581.400 163.200 584.400 163.800 ;
        RECT 648.600 163.200 660.600 164.400 ;
        RECT 315.000 162.600 321.000 163.200 ;
        RECT 360.600 162.600 364.800 163.200 ;
        RECT 460.200 162.600 466.800 163.200 ;
        RECT 469.200 162.600 472.800 163.200 ;
        RECT 519.600 162.600 522.600 163.200 ;
        RECT 315.000 162.000 321.600 162.600 ;
        RECT 361.200 162.000 365.400 162.600 ;
        RECT 461.400 162.000 466.800 162.600 ;
        RECT 314.400 161.400 322.200 162.000 ;
        RECT 361.800 161.400 366.600 162.000 ;
        RECT 462.000 161.400 466.800 162.000 ;
        RECT 469.800 162.000 472.800 162.600 ;
        RECT 519.000 162.000 522.600 162.600 ;
        RECT 580.800 162.000 584.400 163.200 ;
        RECT 649.200 162.000 660.000 163.200 ;
        RECT 469.800 161.400 473.400 162.000 ;
        RECT 313.800 160.200 317.400 161.400 ;
        RECT 318.600 160.800 322.800 161.400 ;
        RECT 362.400 160.800 367.200 161.400 ;
        RECT 463.200 160.800 467.400 161.400 ;
        RECT 319.200 160.200 323.400 160.800 ;
        RECT 363.000 160.200 368.400 160.800 ;
        RECT 463.800 160.200 467.400 160.800 ;
        RECT 470.400 160.800 473.400 161.400 ;
        RECT 518.400 161.400 522.000 162.000 ;
        RECT 580.800 161.400 583.800 162.000 ;
        RECT 649.800 161.400 659.400 162.000 ;
        RECT 518.400 160.800 521.400 161.400 ;
        RECT 470.400 160.200 474.000 160.800 ;
        RECT 517.800 160.200 521.400 160.800 ;
        RECT 580.200 160.800 583.800 161.400 ;
        RECT 650.400 160.800 659.400 161.400 ;
        RECT 313.200 159.600 316.800 160.200 ;
        RECT 319.800 159.600 324.000 160.200 ;
        RECT 363.600 159.600 369.600 160.200 ;
        RECT 184.200 158.400 186.600 159.000 ;
        RECT 312.600 158.400 316.200 159.600 ;
        RECT 320.400 159.000 324.600 159.600 ;
        RECT 364.800 159.000 370.800 159.600 ;
        RECT 464.400 159.000 468.000 160.200 ;
        RECT 471.000 159.000 474.000 160.200 ;
        RECT 517.200 159.600 520.800 160.200 ;
        RECT 580.200 159.600 583.200 160.800 ;
        RECT 651.000 160.200 658.800 160.800 ;
        RECT 651.600 159.600 658.200 160.200 ;
        RECT 321.000 158.400 325.200 159.000 ;
        RECT 365.400 158.400 372.600 159.000 ;
        RECT 465.000 158.400 468.600 159.000 ;
        RECT 184.200 154.200 187.200 158.400 ;
        RECT 312.000 157.800 315.600 158.400 ;
        RECT 321.600 157.800 325.800 158.400 ;
        RECT 366.600 157.800 374.400 158.400 ;
        RECT 465.600 157.800 468.600 158.400 ;
        RECT 311.400 157.200 315.000 157.800 ;
        RECT 322.200 157.200 326.400 157.800 ;
        RECT 367.800 157.200 376.800 157.800 ;
        RECT 465.600 157.200 469.200 157.800 ;
        RECT 471.600 157.200 474.600 159.000 ;
        RECT 516.600 158.400 520.200 159.600 ;
        RECT 579.600 159.000 583.200 159.600 ;
        RECT 646.800 159.000 650.400 159.600 ;
        RECT 652.800 159.000 657.000 159.600 ;
        RECT 579.600 158.400 582.600 159.000 ;
        RECT 516.000 157.800 519.600 158.400 ;
        RECT 579.000 157.800 582.600 158.400 ;
        RECT 645.600 158.400 651.000 159.000 ;
        RECT 645.600 157.800 652.200 158.400 ;
        RECT 515.400 157.200 519.000 157.800 ;
        RECT 310.800 156.600 314.400 157.200 ;
        RECT 322.800 156.600 327.600 157.200 ;
        RECT 369.000 156.600 379.200 157.200 ;
        RECT 438.000 156.600 440.400 157.200 ;
        RECT 456.000 156.600 458.400 157.200 ;
        RECT 465.600 156.600 469.800 157.200 ;
        RECT 310.200 156.000 314.400 156.600 ;
        RECT 323.400 156.000 328.200 156.600 ;
        RECT 370.800 156.000 381.600 156.600 ;
        RECT 438.000 156.000 441.600 156.600 ;
        RECT 454.800 156.000 459.600 156.600 ;
        RECT 466.200 156.000 470.400 156.600 ;
        RECT 310.200 155.400 313.800 156.000 ;
        RECT 324.000 155.400 328.800 156.000 ;
        RECT 372.000 155.400 384.600 156.000 ;
        RECT 438.000 155.400 442.200 156.000 ;
        RECT 454.200 155.400 460.200 156.000 ;
        RECT 309.600 154.800 313.200 155.400 ;
        RECT 325.200 154.800 329.400 155.400 ;
        RECT 374.400 154.800 388.200 155.400 ;
        RECT 438.600 154.800 442.800 155.400 ;
        RECT 454.200 154.800 460.800 155.400 ;
        RECT 466.200 154.800 471.000 156.000 ;
        RECT 472.200 154.800 475.200 157.200 ;
        RECT 514.800 156.600 518.400 157.200 ;
        RECT 579.000 156.600 582.000 157.800 ;
        RECT 645.600 156.600 652.800 157.800 ;
        RECT 514.200 156.000 518.400 156.600 ;
        RECT 578.400 156.000 582.000 156.600 ;
        RECT 646.200 156.000 653.400 156.600 ;
        RECT 513.600 155.400 517.800 156.000 ;
        RECT 513.600 154.800 517.200 155.400 ;
        RECT 578.400 154.800 581.400 156.000 ;
        RECT 648.000 155.400 653.400 156.000 ;
        RECT 309.000 154.200 312.600 154.800 ;
        RECT 325.800 154.200 330.000 154.800 ;
        RECT 376.200 154.200 393.000 154.800 ;
        RECT 439.200 154.200 444.000 154.800 ;
        RECT 454.200 154.200 461.400 154.800 ;
        RECT 466.200 154.200 475.200 154.800 ;
        RECT 513.000 154.200 516.600 154.800 ;
        RECT 184.800 153.600 187.200 154.200 ;
        RECT 308.400 153.600 312.000 154.200 ;
        RECT 326.400 153.600 330.600 154.200 ;
        RECT 378.600 153.600 397.200 154.200 ;
        RECT 439.800 153.600 444.600 154.200 ;
        RECT 184.800 150.000 187.800 153.600 ;
        RECT 307.800 153.000 311.400 153.600 ;
        RECT 327.000 153.000 331.200 153.600 ;
        RECT 381.600 153.000 399.000 153.600 ;
        RECT 441.000 153.000 444.600 153.600 ;
        RECT 307.200 152.400 311.400 153.000 ;
        RECT 327.600 152.400 332.400 153.000 ;
        RECT 385.200 152.400 400.800 153.000 ;
        RECT 441.600 152.400 445.200 153.000 ;
        RECT 306.600 151.800 310.800 152.400 ;
        RECT 328.200 151.800 333.000 152.400 ;
        RECT 388.800 151.800 402.600 152.400 ;
        RECT 442.200 151.800 445.800 152.400 ;
        RECT 306.000 151.200 310.200 151.800 ;
        RECT 328.800 151.200 333.600 151.800 ;
        RECT 393.600 151.200 404.400 151.800 ;
        RECT 305.400 150.600 309.600 151.200 ;
        RECT 330.000 150.600 334.200 151.200 ;
        RECT 396.600 150.600 405.600 151.200 ;
        RECT 442.800 150.600 446.400 151.800 ;
        RECT 453.600 150.600 456.600 154.200 ;
        RECT 457.800 153.600 462.000 154.200 ;
        RECT 458.400 153.000 462.600 153.600 ;
        RECT 459.000 152.400 462.600 153.000 ;
        RECT 459.600 151.800 463.200 152.400 ;
        RECT 460.200 151.200 463.200 151.800 ;
        RECT 466.200 151.200 475.800 154.200 ;
        RECT 512.400 153.600 516.000 154.200 ;
        RECT 577.800 153.600 580.800 154.800 ;
        RECT 648.600 154.200 653.400 155.400 ;
        RECT 645.600 153.600 653.400 154.200 ;
        RECT 511.800 153.000 515.400 153.600 ;
        RECT 511.200 152.400 515.400 153.000 ;
        RECT 577.200 153.000 580.800 153.600 ;
        RECT 644.400 153.000 653.400 153.600 ;
        RECT 577.200 152.400 580.200 153.000 ;
        RECT 510.600 151.800 514.800 152.400 ;
        RECT 576.600 151.800 580.200 152.400 ;
        RECT 643.800 152.400 652.800 153.000 ;
        RECT 643.800 151.800 652.200 152.400 ;
        RECT 510.000 151.200 514.200 151.800 ;
        RECT 460.200 150.600 463.800 151.200 ;
        RECT 304.200 150.000 309.000 150.600 ;
        RECT 330.600 150.000 335.400 150.600 ;
        RECT 398.400 150.000 408.000 150.600 ;
        RECT 443.400 150.000 447.000 150.600 ;
        RECT 185.400 149.400 187.800 150.000 ;
        RECT 303.600 149.400 308.400 150.000 ;
        RECT 331.200 149.400 336.000 150.000 ;
        RECT 400.800 149.400 409.800 150.000 ;
        RECT 444.000 149.400 447.600 150.000 ;
        RECT 185.400 145.800 188.400 149.400 ;
        RECT 303.000 148.800 307.800 149.400 ;
        RECT 331.800 148.800 336.600 149.400 ;
        RECT 402.000 148.800 411.000 149.400 ;
        RECT 444.600 148.800 447.600 149.400 ;
        RECT 454.200 148.800 457.200 150.600 ;
        RECT 460.800 150.000 463.800 150.600 ;
        RECT 460.800 149.400 464.400 150.000 ;
        RECT 302.400 148.200 306.600 148.800 ;
        RECT 332.400 148.200 337.200 148.800 ;
        RECT 402.000 148.200 412.800 148.800 ;
        RECT 444.600 148.200 448.200 148.800 ;
        RECT 454.200 148.200 457.800 148.800 ;
        RECT 461.400 148.200 464.400 149.400 ;
        RECT 466.200 148.200 469.200 151.200 ;
        RECT 470.400 150.000 475.800 151.200 ;
        RECT 509.400 150.600 513.600 151.200 ;
        RECT 576.600 150.600 579.600 151.800 ;
        RECT 643.800 151.200 651.600 151.800 ;
        RECT 643.800 150.600 651.000 151.200 ;
        RECT 508.800 150.000 513.000 150.600 ;
        RECT 471.000 148.800 475.800 150.000 ;
        RECT 508.200 149.400 512.400 150.000 ;
        RECT 576.000 149.400 579.000 150.600 ;
        RECT 644.400 150.000 651.000 150.600 ;
        RECT 645.000 149.400 651.000 150.000 ;
        RECT 507.600 148.800 511.800 149.400 ;
        RECT 575.400 148.800 579.000 149.400 ;
        RECT 471.000 148.200 475.200 148.800 ;
        RECT 507.000 148.200 511.200 148.800 ;
        RECT 575.400 148.200 578.400 148.800 ;
        RECT 641.400 148.200 643.800 148.800 ;
        RECT 646.200 148.200 651.000 149.400 ;
        RECT 301.200 147.600 306.600 148.200 ;
        RECT 333.600 147.600 338.400 148.200 ;
        RECT 402.600 147.600 414.600 148.200 ;
        RECT 445.200 147.600 448.200 148.200 ;
        RECT 300.600 147.000 306.600 147.600 ;
        RECT 334.200 147.000 339.000 147.600 ;
        RECT 403.200 147.000 415.800 147.600 ;
        RECT 445.200 147.000 448.800 147.600 ;
        RECT 299.400 146.400 306.600 147.000 ;
        RECT 334.800 146.400 339.600 147.000 ;
        RECT 404.400 146.400 417.600 147.000 ;
        RECT 445.800 146.400 448.800 147.000 ;
        RECT 454.800 147.000 457.800 148.200 ;
        RECT 462.000 147.000 469.200 148.200 ;
        RECT 454.800 146.400 458.400 147.000 ;
        RECT 462.000 146.400 468.600 147.000 ;
        RECT 471.600 146.400 475.200 148.200 ;
        RECT 505.800 147.600 510.600 148.200 ;
        RECT 574.800 147.600 578.400 148.200 ;
        RECT 505.200 147.000 510.000 147.600 ;
        RECT 574.800 147.000 577.800 147.600 ;
        RECT 504.600 146.400 509.400 147.000 ;
        RECT 574.200 146.400 577.800 147.000 ;
        RECT 640.800 146.400 650.400 148.200 ;
        RECT 298.800 145.800 306.600 146.400 ;
        RECT 336.000 145.800 340.800 146.400 ;
        RECT 405.000 145.800 418.800 146.400 ;
        RECT 438.000 145.800 439.200 146.400 ;
        RECT 445.800 145.800 449.400 146.400 ;
        RECT 186.000 145.200 188.400 145.800 ;
        RECT 186.000 142.200 189.000 145.200 ;
        RECT 297.600 144.600 306.000 145.800 ;
        RECT 336.600 145.200 341.400 145.800 ;
        RECT 405.600 145.200 419.400 145.800 ;
        RECT 436.200 145.200 441.000 145.800 ;
        RECT 446.400 145.200 449.400 145.800 ;
        RECT 455.400 145.800 458.400 146.400 ;
        RECT 462.600 145.800 468.600 146.400 ;
        RECT 472.200 145.800 474.600 146.400 ;
        RECT 504.000 145.800 508.200 146.400 ;
        RECT 455.400 145.200 459.000 145.800 ;
        RECT 337.200 144.600 342.000 145.200 ;
        RECT 406.800 144.600 412.800 145.200 ;
        RECT 414.000 144.600 420.000 145.200 ;
        RECT 435.600 144.600 441.600 145.200 ;
        RECT 446.400 144.600 450.000 145.200 ;
        RECT 297.000 144.000 301.200 144.600 ;
        RECT 297.000 143.400 300.000 144.000 ;
        RECT 303.000 142.800 306.000 144.600 ;
        RECT 337.800 144.000 343.200 144.600 ;
        RECT 407.400 144.000 412.800 144.600 ;
        RECT 415.200 144.000 420.600 144.600 ;
        RECT 435.000 144.000 442.200 144.600 ;
        RECT 339.000 143.400 343.800 144.000 ;
        RECT 408.600 143.400 413.400 144.000 ;
        RECT 416.400 143.400 420.600 144.000 ;
        RECT 434.400 143.400 442.800 144.000 ;
        RECT 447.000 143.400 450.000 144.600 ;
        RECT 456.000 144.600 459.000 145.200 ;
        RECT 462.600 145.200 468.000 145.800 ;
        RECT 472.800 145.200 474.000 145.800 ;
        RECT 503.400 145.200 507.600 145.800 ;
        RECT 574.200 145.200 577.200 146.400 ;
        RECT 641.400 145.800 649.800 146.400 ;
        RECT 641.400 145.200 649.200 145.800 ;
        RECT 456.000 144.000 459.600 144.600 ;
        RECT 456.600 143.400 459.600 144.000 ;
        RECT 462.600 144.000 467.400 145.200 ;
        RECT 502.200 144.600 507.000 145.200 ;
        RECT 501.600 144.000 506.400 144.600 ;
        RECT 573.600 144.000 576.600 145.200 ;
        RECT 642.600 144.600 648.600 145.200 ;
        RECT 643.200 144.000 648.000 144.600 ;
        RECT 462.600 143.400 466.800 144.000 ;
        RECT 501.000 143.400 505.800 144.000 ;
        RECT 573.000 143.400 576.600 144.000 ;
        RECT 339.600 142.800 345.000 143.400 ;
        RECT 409.200 142.800 414.600 143.400 ;
        RECT 186.600 141.600 189.000 142.200 ;
        RECT 186.600 138.600 189.600 141.600 ;
        RECT 302.400 141.000 305.400 142.800 ;
        RECT 340.800 142.200 345.600 142.800 ;
        RECT 410.400 142.200 415.200 142.800 ;
        RECT 417.600 142.200 421.200 143.400 ;
        RECT 434.400 142.800 443.400 143.400 ;
        RECT 433.800 142.200 437.400 142.800 ;
        RECT 341.400 141.600 346.800 142.200 ;
        RECT 411.000 141.600 415.800 142.200 ;
        RECT 418.200 141.600 421.800 142.200 ;
        RECT 342.000 141.000 347.400 141.600 ;
        RECT 411.600 141.000 417.000 141.600 ;
        RECT 418.800 141.000 421.800 141.600 ;
        RECT 301.800 140.400 305.400 141.000 ;
        RECT 343.200 140.400 348.600 141.000 ;
        RECT 412.800 140.400 417.600 141.000 ;
        RECT 418.800 140.400 422.400 141.000 ;
        RECT 301.800 138.600 304.800 140.400 ;
        RECT 343.800 139.800 349.200 140.400 ;
        RECT 413.400 139.800 423.000 140.400 ;
        RECT 345.000 139.200 350.400 139.800 ;
        RECT 414.600 139.200 423.000 139.800 ;
        RECT 345.600 138.600 351.600 139.200 ;
        RECT 415.200 138.600 423.600 139.200 ;
        RECT 187.200 135.000 190.200 138.600 ;
        RECT 301.200 136.800 304.200 138.600 ;
        RECT 346.800 138.000 352.200 138.600 ;
        RECT 415.800 138.000 424.200 138.600 ;
        RECT 433.800 138.000 436.800 142.200 ;
        RECT 440.400 141.600 444.000 142.800 ;
        RECT 447.600 141.600 450.600 143.400 ;
        RECT 456.600 142.800 460.200 143.400 ;
        RECT 457.200 142.200 460.800 142.800 ;
        RECT 462.600 142.200 466.200 143.400 ;
        RECT 499.800 142.800 504.600 143.400 ;
        RECT 573.000 142.800 576.000 143.400 ;
        RECT 639.000 142.800 643.200 143.400 ;
        RECT 499.200 142.200 504.000 142.800 ;
        RECT 572.400 142.200 576.000 142.800 ;
        RECT 638.400 142.200 643.800 142.800 ;
        RECT 457.200 141.600 461.400 142.200 ;
        RECT 441.000 141.000 444.000 141.600 ;
        RECT 448.200 141.000 452.400 141.600 ;
        RECT 457.800 141.000 461.400 141.600 ;
        RECT 441.600 139.200 444.600 141.000 ;
        RECT 448.200 140.400 453.600 141.000 ;
        RECT 457.800 140.400 462.000 141.000 ;
        RECT 448.200 139.800 462.000 140.400 ;
        RECT 463.200 139.800 465.600 142.200 ;
        RECT 498.000 141.600 503.400 142.200 ;
        RECT 572.400 141.600 575.400 142.200 ;
        RECT 637.800 141.600 644.400 142.200 ;
        RECT 497.400 141.000 502.200 141.600 ;
        RECT 571.800 141.000 575.400 141.600 ;
        RECT 637.200 141.000 645.000 141.600 ;
        RECT 496.200 140.400 501.600 141.000 ;
        RECT 571.800 140.400 574.800 141.000 ;
        RECT 621.600 140.400 622.200 141.000 ;
        RECT 636.600 140.400 645.000 141.000 ;
        RECT 495.600 139.800 501.000 140.400 ;
        RECT 571.200 139.800 574.800 140.400 ;
        RECT 620.400 139.800 623.400 140.400 ;
        RECT 448.200 139.200 465.600 139.800 ;
        RECT 494.400 139.200 499.800 139.800 ;
        RECT 571.200 139.200 574.200 139.800 ;
        RECT 348.000 137.400 353.400 138.000 ;
        RECT 416.400 137.400 424.200 138.000 ;
        RECT 348.600 136.800 354.600 137.400 ;
        RECT 417.600 136.800 424.800 137.400 ;
        RECT 434.400 136.800 437.400 138.000 ;
        RECT 442.200 136.800 445.200 139.200 ;
        RECT 448.800 138.000 465.600 139.200 ;
        RECT 493.800 138.600 499.200 139.200 ;
        RECT 570.600 138.600 574.200 139.200 ;
        RECT 619.800 139.200 624.600 139.800 ;
        RECT 636.000 139.200 645.600 140.400 ;
        RECT 619.800 138.600 625.800 139.200 ;
        RECT 492.600 138.000 498.000 138.600 ;
        RECT 570.600 138.000 573.600 138.600 ;
        RECT 448.800 136.800 451.800 138.000 ;
        RECT 453.600 137.400 458.400 138.000 ;
        RECT 300.600 135.000 303.600 136.800 ;
        RECT 349.800 136.200 355.200 136.800 ;
        RECT 418.200 136.200 425.400 136.800 ;
        RECT 434.400 136.200 438.000 136.800 ;
        RECT 350.400 135.600 356.400 136.200 ;
        RECT 418.800 135.600 426.000 136.200 ;
        RECT 435.000 135.600 438.000 136.200 ;
        RECT 442.800 136.200 445.200 136.800 ;
        RECT 448.200 136.200 451.800 136.800 ;
        RECT 460.200 136.200 465.600 138.000 ;
        RECT 491.400 137.400 497.400 138.000 ;
        RECT 570.000 137.400 573.600 138.000 ;
        RECT 620.400 138.000 627.000 138.600 ;
        RECT 635.400 138.000 640.200 139.200 ;
        RECT 641.400 138.000 645.600 139.200 ;
        RECT 620.400 137.400 627.600 138.000 ;
        RECT 490.800 136.800 496.200 137.400 ;
        RECT 570.000 136.800 573.000 137.400 ;
        RECT 621.000 136.800 629.400 137.400 ;
        RECT 489.600 136.200 495.000 136.800 ;
        RECT 569.400 136.200 573.000 136.800 ;
        RECT 622.200 136.200 630.000 136.800 ;
        RECT 636.000 136.200 645.600 138.000 ;
        RECT 351.600 135.000 357.600 135.600 ;
        RECT 419.400 135.000 426.600 135.600 ;
        RECT 435.000 135.000 438.600 135.600 ;
        RECT 187.800 132.000 190.800 135.000 ;
        RECT 263.400 134.400 264.000 135.000 ;
        RECT 262.800 133.800 264.600 134.400 ;
        RECT 262.800 132.600 265.200 133.800 ;
        RECT 300.000 133.200 303.000 135.000 ;
        RECT 352.800 134.400 358.800 135.000 ;
        RECT 420.000 134.400 427.200 135.000 ;
        RECT 435.600 134.400 438.600 135.000 ;
        RECT 442.800 134.400 445.800 136.200 ;
        RECT 448.200 135.600 451.200 136.200 ;
        RECT 447.600 135.000 451.200 135.600 ;
        RECT 447.000 134.400 450.600 135.000 ;
        RECT 460.800 134.400 465.600 136.200 ;
        RECT 488.400 135.600 494.400 136.200 ;
        RECT 569.400 135.600 572.400 136.200 ;
        RECT 619.200 135.600 621.000 136.200 ;
        RECT 622.800 135.600 631.800 136.200 ;
        RECT 636.600 135.600 645.000 136.200 ;
        RECT 487.200 135.000 493.200 135.600 ;
        RECT 568.800 135.000 572.400 135.600 ;
        RECT 618.000 135.000 621.600 135.600 ;
        RECT 624.000 135.000 632.400 135.600 ;
        RECT 636.600 135.000 644.400 135.600 ;
        RECT 486.000 134.400 492.000 135.000 ;
        RECT 568.800 134.400 571.800 135.000 ;
        RECT 354.000 133.800 360.000 134.400 ;
        RECT 420.600 133.800 427.800 134.400 ;
        RECT 435.600 133.800 439.200 134.400 ;
        RECT 354.600 133.200 361.200 133.800 ;
        RECT 421.800 133.200 429.000 133.800 ;
        RECT 436.200 133.200 439.800 133.800 ;
        RECT 442.800 133.200 450.000 134.400 ;
        RECT 188.400 129.000 191.400 132.000 ;
        RECT 262.800 131.400 265.800 132.600 ;
        RECT 299.400 131.400 302.400 133.200 ;
        RECT 355.800 132.600 362.400 133.200 ;
        RECT 422.400 132.600 430.800 133.200 ;
        RECT 436.200 132.600 440.400 133.200 ;
        RECT 357.000 132.000 363.600 132.600 ;
        RECT 423.000 132.000 440.400 132.600 ;
        RECT 442.800 132.600 449.400 133.200 ;
        RECT 461.400 132.600 465.600 134.400 ;
        RECT 484.800 133.800 491.400 134.400 ;
        RECT 568.200 133.800 571.800 134.400 ;
        RECT 483.600 133.200 490.200 133.800 ;
        RECT 568.200 133.200 571.200 133.800 ;
        RECT 617.400 133.200 621.600 135.000 ;
        RECT 625.200 134.400 634.200 135.000 ;
        RECT 637.200 134.400 644.400 135.000 ;
        RECT 626.400 133.800 634.800 134.400 ;
        RECT 638.400 133.800 643.200 134.400 ;
        RECT 627.000 133.200 636.600 133.800 ;
        RECT 639.000 133.200 642.600 133.800 ;
        RECT 482.400 132.600 489.000 133.200 ;
        RECT 567.600 132.600 571.200 133.200 ;
        RECT 616.800 132.600 621.600 133.200 ;
        RECT 628.200 132.600 637.200 133.200 ;
        RECT 442.800 132.000 448.800 132.600 ;
        RECT 462.000 132.000 465.600 132.600 ;
        RECT 481.200 132.000 487.800 132.600 ;
        RECT 567.000 132.000 570.600 132.600 ;
        RECT 358.200 131.400 364.800 132.000 ;
        RECT 423.600 131.400 441.000 132.000 ;
        RECT 442.800 131.400 447.600 132.000 ;
        RECT 462.000 131.400 465.000 132.000 ;
        RECT 479.400 131.400 486.600 132.000 ;
        RECT 567.000 131.400 570.000 132.000 ;
        RECT 263.400 130.200 266.400 131.400 ;
        RECT 298.800 130.200 301.800 131.400 ;
        RECT 359.400 130.800 366.000 131.400 ;
        RECT 424.200 130.800 441.600 131.400 ;
        RECT 442.800 130.800 447.000 131.400 ;
        RECT 462.600 130.800 465.000 131.400 ;
        RECT 478.200 130.800 485.400 131.400 ;
        RECT 566.400 130.800 570.000 131.400 ;
        RECT 616.800 131.400 621.000 132.600 ;
        RECT 629.400 132.000 639.000 132.600 ;
        RECT 630.600 131.400 639.600 132.000 ;
        RECT 616.800 130.800 621.600 131.400 ;
        RECT 631.800 130.800 640.800 131.400 ;
        RECT 360.600 130.200 367.200 130.800 ;
        RECT 424.800 130.200 445.800 130.800 ;
        RECT 477.000 130.200 484.200 130.800 ;
        RECT 566.400 130.200 569.400 130.800 ;
        RECT 616.800 130.200 622.200 130.800 ;
        RECT 633.000 130.200 640.800 130.800 ;
        RECT 264.000 129.600 267.000 130.200 ;
        RECT 298.200 129.600 301.800 130.200 ;
        RECT 361.800 129.600 369.000 130.200 ;
        RECT 425.400 129.600 436.800 130.200 ;
        RECT 438.600 129.600 445.800 130.200 ;
        RECT 475.200 129.600 483.000 130.200 ;
        RECT 565.800 129.600 569.400 130.200 ;
        RECT 617.400 129.600 622.800 130.200 ;
        RECT 634.200 129.600 641.400 130.200 ;
        RECT 264.000 129.000 267.600 129.600 ;
        RECT 189.000 126.000 192.000 129.000 ;
        RECT 264.600 128.400 267.600 129.000 ;
        RECT 298.200 128.400 301.200 129.600 ;
        RECT 363.000 129.000 370.200 129.600 ;
        RECT 426.000 129.000 430.200 129.600 ;
        RECT 364.200 128.400 371.400 129.000 ;
        RECT 426.600 128.400 430.200 129.000 ;
        RECT 439.200 128.400 445.800 129.600 ;
        RECT 474.000 129.000 481.200 129.600 ;
        RECT 565.800 129.000 568.800 129.600 ;
        RECT 617.400 129.000 623.400 129.600 ;
        RECT 629.400 129.000 631.200 129.600 ;
        RECT 636.000 129.000 641.400 129.600 ;
        RECT 472.200 128.400 480.000 129.000 ;
        RECT 565.200 128.400 568.800 129.000 ;
        RECT 618.000 128.400 624.600 129.000 ;
        RECT 264.600 127.200 268.200 128.400 ;
        RECT 297.600 127.200 300.600 128.400 ;
        RECT 365.400 127.800 373.200 128.400 ;
        RECT 367.200 127.200 375.000 127.800 ;
        RECT 427.200 127.200 430.800 128.400 ;
        RECT 439.800 127.200 445.800 128.400 ;
        RECT 470.400 127.800 478.800 128.400 ;
        RECT 468.600 127.200 477.000 127.800 ;
        RECT 564.600 127.200 568.200 128.400 ;
        RECT 618.600 127.800 625.200 128.400 ;
        RECT 628.200 127.800 631.800 129.000 ;
        RECT 636.600 128.400 641.400 129.000 ;
        RECT 638.400 127.800 640.800 128.400 ;
        RECT 619.200 127.200 631.800 127.800 ;
        RECT 265.200 126.600 268.800 127.200 ;
        RECT 265.800 126.000 268.800 126.600 ;
        RECT 297.000 126.600 300.600 127.200 ;
        RECT 368.400 126.600 376.200 127.200 ;
        RECT 427.800 126.600 431.400 127.200 ;
        RECT 439.800 126.600 445.200 127.200 ;
        RECT 467.400 126.600 475.800 127.200 ;
        RECT 564.000 126.600 567.600 127.200 ;
        RECT 619.800 126.600 631.800 127.200 ;
        RECT 189.600 123.600 192.600 126.000 ;
        RECT 265.800 125.400 269.400 126.000 ;
        RECT 297.000 125.400 300.000 126.600 ;
        RECT 369.600 126.000 378.000 126.600 ;
        RECT 428.400 126.000 431.400 126.600 ;
        RECT 371.400 125.400 379.800 126.000 ;
        RECT 266.400 124.800 269.400 125.400 ;
        RECT 247.800 124.200 249.600 124.800 ;
        RECT 266.400 124.200 270.000 124.800 ;
        RECT 296.400 124.200 299.400 125.400 ;
        RECT 372.600 124.800 381.600 125.400 ;
        RECT 428.400 124.800 432.000 126.000 ;
        RECT 374.400 124.200 384.000 124.800 ;
        RECT 429.000 124.200 432.000 124.800 ;
        RECT 440.400 125.400 445.200 126.600 ;
        RECT 465.600 126.000 474.000 126.600 ;
        RECT 564.000 126.000 567.000 126.600 ;
        RECT 620.400 126.000 631.800 126.600 ;
        RECT 463.200 125.400 472.800 126.000 ;
        RECT 563.400 125.400 567.000 126.000 ;
        RECT 621.600 125.400 631.800 126.000 ;
        RECT 440.400 124.200 444.600 125.400 ;
        RECT 461.400 124.800 471.000 125.400 ;
        RECT 459.000 124.200 469.200 124.800 ;
        RECT 562.800 124.200 566.400 125.400 ;
        RECT 622.200 124.800 632.400 125.400 ;
        RECT 623.400 124.200 633.600 124.800 ;
        RECT 190.200 120.600 193.200 123.600 ;
        RECT 247.200 120.600 250.200 124.200 ;
        RECT 267.000 123.000 270.600 124.200 ;
        RECT 295.800 123.600 299.400 124.200 ;
        RECT 376.200 123.600 385.800 124.200 ;
        RECT 295.800 123.000 298.800 123.600 ;
        RECT 378.000 123.000 388.200 123.600 ;
        RECT 267.600 121.800 271.200 123.000 ;
        RECT 295.200 122.400 298.800 123.000 ;
        RECT 379.800 122.400 391.200 123.000 ;
        RECT 429.000 122.400 432.600 124.200 ;
        RECT 441.000 123.600 444.600 124.200 ;
        RECT 456.600 123.600 467.400 124.200 ;
        RECT 562.200 123.600 565.800 124.200 ;
        RECT 624.000 123.600 634.800 124.200 ;
        RECT 441.600 123.000 444.000 123.600 ;
        RECT 453.600 123.000 465.600 123.600 ;
        RECT 562.200 123.000 565.200 123.600 ;
        RECT 441.600 122.400 443.400 123.000 ;
        RECT 450.600 122.400 463.200 123.000 ;
        RECT 561.600 122.400 565.200 123.000 ;
        RECT 624.600 123.000 635.400 123.600 ;
        RECT 268.200 121.200 271.800 121.800 ;
        RECT 295.200 121.200 298.200 122.400 ;
        RECT 381.600 121.800 393.600 122.400 ;
        RECT 384.000 121.200 396.600 121.800 ;
        RECT 429.600 121.200 432.600 122.400 ;
        RECT 447.600 121.800 461.400 122.400 ;
        RECT 561.000 121.800 564.600 122.400 ;
        RECT 624.600 121.800 636.000 123.000 ;
        RECT 444.000 121.200 459.000 121.800 ;
        RECT 561.000 121.200 564.000 121.800 ;
        RECT 625.200 121.200 636.000 121.800 ;
        RECT 268.200 120.600 272.400 121.200 ;
        RECT 190.800 118.200 193.800 120.600 ;
        RECT 247.800 118.200 250.800 120.600 ;
        RECT 268.800 120.000 272.400 120.600 ;
        RECT 294.600 120.000 297.600 121.200 ;
        RECT 385.800 120.600 400.800 121.200 ;
        RECT 388.200 120.000 405.000 120.600 ;
        RECT 430.200 120.000 433.200 121.200 ;
        RECT 440.400 120.600 456.600 121.200 ;
        RECT 560.400 120.600 564.000 121.200 ;
        RECT 625.800 120.600 627.600 121.200 ;
        RECT 631.200 120.600 636.000 121.200 ;
        RECT 435.000 120.000 453.600 120.600 ;
        RECT 269.400 118.800 273.000 120.000 ;
        RECT 294.000 118.800 297.000 120.000 ;
        RECT 391.200 119.400 412.800 120.000 ;
        RECT 427.800 119.400 450.600 120.000 ;
        RECT 559.800 119.400 563.400 120.600 ;
        RECT 622.200 120.000 624.000 120.600 ;
        RECT 633.000 120.000 635.400 120.600 ;
        RECT 621.600 119.400 624.600 120.000 ;
        RECT 393.600 118.800 447.600 119.400 ;
        RECT 559.200 118.800 562.800 119.400 ;
        RECT 621.000 118.800 625.200 119.400 ;
        RECT 270.000 118.200 273.600 118.800 ;
        RECT 293.400 118.200 296.400 118.800 ;
        RECT 397.200 118.200 444.000 118.800 ;
        RECT 191.400 115.800 194.400 118.200 ;
        RECT 248.400 117.000 251.400 118.200 ;
        RECT 270.600 117.000 274.200 118.200 ;
        RECT 292.800 117.600 296.400 118.200 ;
        RECT 400.800 117.600 439.800 118.200 ;
        RECT 558.600 117.600 562.200 118.800 ;
        RECT 620.400 118.200 625.200 118.800 ;
        RECT 619.800 117.600 625.200 118.200 ;
        RECT 292.800 117.000 295.800 117.600 ;
        RECT 405.600 117.000 434.400 117.600 ;
        RECT 558.000 117.000 561.600 117.600 ;
        RECT 619.800 117.000 624.600 117.600 ;
        RECT 248.400 116.400 252.000 117.000 ;
        RECT 192.000 113.400 195.000 115.800 ;
        RECT 249.000 115.200 252.000 116.400 ;
        RECT 271.200 116.400 274.800 117.000 ;
        RECT 292.200 116.400 295.800 117.000 ;
        RECT 414.000 116.400 426.000 117.000 ;
        RECT 557.400 116.400 561.000 117.000 ;
        RECT 271.200 115.200 275.400 116.400 ;
        RECT 292.200 115.800 295.200 116.400 ;
        RECT 291.600 115.200 295.200 115.800 ;
        RECT 556.800 115.200 560.400 116.400 ;
        RECT 249.000 114.600 252.600 115.200 ;
        RECT 249.600 114.000 252.600 114.600 ;
        RECT 271.200 114.600 276.000 115.200 ;
        RECT 291.600 114.600 294.600 115.200 ;
        RECT 556.200 114.600 559.800 115.200 ;
        RECT 271.200 114.000 276.600 114.600 ;
        RECT 291.000 114.000 294.600 114.600 ;
        RECT 555.600 114.000 559.200 114.600 ;
        RECT 249.600 113.400 253.200 114.000 ;
        RECT 192.600 111.000 195.600 113.400 ;
        RECT 250.200 112.800 253.200 113.400 ;
        RECT 271.200 112.800 277.200 114.000 ;
        RECT 290.400 113.400 294.000 114.000 ;
        RECT 555.000 113.400 559.200 114.000 ;
        RECT 619.800 114.000 624.000 117.000 ;
        RECT 619.800 113.400 624.600 114.000 ;
        RECT 290.400 112.800 293.400 113.400 ;
        RECT 555.000 112.800 558.600 113.400 ;
        RECT 619.800 112.800 625.800 113.400 ;
        RECT 229.800 112.200 231.000 112.800 ;
        RECT 250.200 112.200 253.800 112.800 ;
        RECT 229.200 111.600 231.600 112.200 ;
        RECT 250.800 111.600 253.800 112.200 ;
        RECT 271.200 112.200 277.800 112.800 ;
        RECT 289.800 112.200 293.400 112.800 ;
        RECT 554.400 112.200 558.000 112.800 ;
        RECT 620.400 112.200 627.600 112.800 ;
        RECT 271.200 111.600 278.400 112.200 ;
        RECT 289.200 111.600 292.800 112.200 ;
        RECT 553.800 111.600 557.400 112.200 ;
        RECT 620.400 111.600 628.800 112.200 ;
        RECT 193.200 109.200 196.200 111.000 ;
        RECT 229.200 110.400 232.200 111.600 ;
        RECT 250.800 111.000 254.400 111.600 ;
        RECT 251.400 110.400 254.400 111.000 ;
        RECT 271.800 111.000 279.000 111.600 ;
        RECT 271.800 110.400 279.600 111.000 ;
        RECT 288.600 110.400 292.200 111.600 ;
        RECT 553.200 111.000 557.400 111.600 ;
        RECT 616.800 111.000 619.200 111.600 ;
        RECT 621.000 111.000 628.800 111.600 ;
        RECT 553.200 110.400 556.800 111.000 ;
        RECT 616.200 110.400 619.200 111.000 ;
        RECT 621.600 110.400 628.800 111.000 ;
        RECT 193.800 107.400 196.800 109.200 ;
        RECT 229.800 108.600 232.800 110.400 ;
        RECT 251.400 109.800 255.000 110.400 ;
        RECT 252.000 109.200 255.000 109.800 ;
        RECT 252.000 108.600 255.600 109.200 ;
        RECT 230.400 107.400 233.400 108.600 ;
        RECT 252.600 108.000 256.200 108.600 ;
        RECT 253.200 107.400 256.200 108.000 ;
        RECT 193.800 106.800 197.400 107.400 ;
        RECT 194.400 105.600 197.400 106.800 ;
        RECT 231.000 106.200 234.000 107.400 ;
        RECT 253.200 106.800 256.800 107.400 ;
        RECT 253.800 106.200 257.400 106.800 ;
        RECT 231.000 105.600 234.600 106.200 ;
        RECT 194.400 105.000 198.000 105.600 ;
        RECT 195.000 104.400 198.000 105.000 ;
        RECT 231.600 105.000 234.600 105.600 ;
        RECT 254.400 105.600 258.000 106.200 ;
        RECT 231.600 104.400 235.200 105.000 ;
        RECT 254.400 104.400 258.600 105.600 ;
        RECT 195.000 103.200 198.600 104.400 ;
        RECT 232.200 103.200 235.800 104.400 ;
        RECT 254.400 103.800 259.200 104.400 ;
        RECT 254.400 103.200 259.800 103.800 ;
        RECT 195.600 102.000 198.600 103.200 ;
        RECT 232.800 102.000 236.400 103.200 ;
        RECT 254.400 102.600 260.400 103.200 ;
        RECT 254.400 102.000 261.600 102.600 ;
        RECT 271.800 102.000 274.800 110.400 ;
        RECT 276.000 109.800 280.200 110.400 ;
        RECT 288.000 109.800 291.600 110.400 ;
        RECT 552.600 109.800 556.200 110.400 ;
        RECT 276.600 109.200 280.800 109.800 ;
        RECT 287.400 109.200 291.000 109.800 ;
        RECT 552.000 109.200 555.600 109.800 ;
        RECT 277.200 108.600 281.400 109.200 ;
        RECT 286.800 108.600 290.400 109.200 ;
        RECT 551.400 108.600 555.000 109.200 ;
        RECT 615.000 108.600 619.200 110.400 ;
        RECT 622.200 109.800 628.800 110.400 ;
        RECT 623.400 109.200 628.800 109.800 ;
        RECT 625.200 108.600 627.600 109.200 ;
        RECT 277.800 108.000 282.000 108.600 ;
        RECT 286.200 108.000 290.400 108.600 ;
        RECT 550.800 108.000 555.000 108.600 ;
        RECT 278.400 107.400 282.600 108.000 ;
        RECT 285.600 107.400 289.800 108.000 ;
        RECT 550.200 107.400 554.400 108.000 ;
        RECT 614.400 107.400 618.600 108.600 ;
        RECT 279.000 106.800 283.200 107.400 ;
        RECT 284.400 106.800 289.200 107.400 ;
        RECT 549.600 106.800 553.800 107.400 ;
        RECT 279.600 106.200 288.600 106.800 ;
        RECT 549.600 106.200 553.200 106.800 ;
        RECT 613.800 106.200 618.000 107.400 ;
        RECT 280.200 105.600 288.000 106.200 ;
        RECT 549.000 105.600 552.600 106.200 ;
        RECT 280.800 105.000 287.400 105.600 ;
        RECT 548.400 105.000 552.000 105.600 ;
        RECT 613.800 105.000 618.600 106.200 ;
        RECT 281.400 104.400 286.800 105.000 ;
        RECT 547.800 104.400 551.400 105.000 ;
        RECT 282.000 103.800 285.600 104.400 ;
        RECT 547.200 103.800 551.400 104.400 ;
        RECT 614.400 104.400 619.200 105.000 ;
        RECT 614.400 103.800 620.400 104.400 ;
        RECT 282.600 103.200 284.400 103.800 ;
        RECT 546.600 103.200 550.800 103.800 ;
        RECT 615.000 103.200 622.200 103.800 ;
        RECT 546.000 102.600 550.200 103.200 ;
        RECT 615.000 102.600 623.400 103.200 ;
        RECT 545.400 102.000 549.600 102.600 ;
        RECT 615.600 102.000 623.400 102.600 ;
        RECT 195.600 100.800 199.200 102.000 ;
        RECT 196.200 100.200 199.200 100.800 ;
        RECT 232.200 100.800 237.000 102.000 ;
        RECT 253.800 101.400 262.200 102.000 ;
        RECT 253.800 100.800 262.800 101.400 ;
        RECT 232.200 100.200 237.600 100.800 ;
        RECT 196.200 99.000 199.800 100.200 ;
        RECT 232.200 99.000 238.200 100.200 ;
        RECT 196.800 98.400 199.800 99.000 ;
        RECT 231.600 98.400 238.800 99.000 ;
        RECT 253.800 98.400 256.800 100.800 ;
        RECT 258.600 100.200 264.000 100.800 ;
        RECT 259.200 99.600 265.200 100.200 ;
        RECT 259.800 99.000 267.600 99.600 ;
        RECT 271.200 99.000 274.800 102.000 ;
        RECT 544.800 101.400 549.000 102.000 ;
        RECT 616.200 101.400 624.000 102.000 ;
        RECT 544.200 100.800 548.400 101.400 ;
        RECT 616.800 100.800 623.400 101.400 ;
        RECT 543.600 100.200 547.800 100.800 ;
        RECT 618.000 100.200 623.400 100.800 ;
        RECT 543.000 99.600 547.200 100.200 ;
        RECT 619.800 99.600 622.800 100.200 ;
        RECT 542.400 99.000 546.600 99.600 ;
        RECT 260.400 98.400 274.200 99.000 ;
        RECT 541.800 98.400 546.000 99.000 ;
        RECT 618.000 98.400 619.800 99.000 ;
        RECT 196.800 97.200 200.400 98.400 ;
        RECT 197.400 96.600 200.400 97.200 ;
        RECT 231.600 96.600 234.600 98.400 ;
        RECT 235.800 97.200 239.400 98.400 ;
        RECT 236.400 96.600 240.000 97.200 ;
        RECT 197.400 96.000 201.000 96.600 ;
        RECT 198.000 95.400 201.000 96.000 ;
        RECT 198.000 94.200 201.600 95.400 ;
        RECT 231.000 94.800 234.000 96.600 ;
        RECT 237.000 96.000 240.600 96.600 ;
        RECT 237.000 95.400 241.200 96.000 ;
        RECT 253.200 95.400 256.200 98.400 ;
        RECT 261.600 97.800 274.200 98.400 ;
        RECT 540.600 97.800 545.400 98.400 ;
        RECT 615.600 97.800 621.000 98.400 ;
        RECT 262.200 97.200 274.200 97.800 ;
        RECT 540.000 97.200 544.800 97.800 ;
        RECT 610.200 97.200 621.000 97.800 ;
        RECT 263.400 96.600 273.600 97.200 ;
        RECT 539.400 96.600 544.200 97.200 ;
        RECT 609.600 96.600 621.000 97.200 ;
        RECT 264.000 96.000 273.000 96.600 ;
        RECT 538.800 96.000 543.000 96.600 ;
        RECT 609.000 96.000 621.000 96.600 ;
        RECT 265.200 95.400 271.800 96.000 ;
        RECT 538.200 95.400 542.400 96.000 ;
        RECT 609.000 95.400 620.400 96.000 ;
        RECT 237.600 94.800 241.200 95.400 ;
        RECT 198.600 93.600 201.600 94.200 ;
        RECT 198.600 92.400 202.200 93.600 ;
        RECT 230.400 93.000 233.400 94.800 ;
        RECT 238.200 94.200 241.800 94.800 ;
        RECT 238.800 93.600 242.400 94.200 ;
        RECT 238.800 93.000 243.000 93.600 ;
        RECT 199.200 91.200 202.800 92.400 ;
        RECT 229.800 91.200 232.800 93.000 ;
        RECT 239.400 92.400 243.600 93.000 ;
        RECT 252.600 92.400 255.600 95.400 ;
        RECT 265.800 94.800 271.800 95.400 ;
        RECT 537.600 94.800 541.800 95.400 ;
        RECT 608.400 94.800 620.400 95.400 ;
        RECT 267.000 94.200 272.400 94.800 ;
        RECT 537.000 94.200 541.200 94.800 ;
        RECT 268.200 93.600 273.600 94.200 ;
        RECT 536.400 93.600 540.600 94.200 ;
        RECT 608.400 93.600 619.200 94.800 ;
        RECT 268.800 93.000 274.800 93.600 ;
        RECT 535.800 93.000 540.000 93.600 ;
        RECT 607.800 93.000 619.200 93.600 ;
        RECT 270.000 92.400 275.400 93.000 ;
        RECT 535.200 92.400 539.400 93.000 ;
        RECT 240.000 91.800 244.200 92.400 ;
        RECT 240.600 91.200 244.200 91.800 ;
        RECT 199.800 90.000 203.400 91.200 ;
        RECT 229.200 90.000 232.200 91.200 ;
        RECT 241.200 90.600 244.800 91.200 ;
        RECT 241.800 90.000 245.400 90.600 ;
        RECT 200.400 89.400 203.400 90.000 ;
        RECT 228.600 89.400 232.200 90.000 ;
        RECT 242.400 89.400 246.000 90.000 ;
        RECT 252.000 89.400 255.000 92.400 ;
        RECT 271.200 91.800 276.600 92.400 ;
        RECT 534.600 91.800 538.800 92.400 ;
        RECT 603.000 91.800 606.000 92.400 ;
        RECT 271.800 91.200 277.800 91.800 ;
        RECT 534.000 91.200 538.200 91.800 ;
        RECT 602.400 91.200 606.000 91.800 ;
        RECT 273.000 90.600 279.000 91.200 ;
        RECT 533.400 90.600 537.600 91.200 ;
        RECT 274.200 90.000 279.600 90.600 ;
        RECT 532.800 90.000 537.000 90.600 ;
        RECT 274.800 89.400 280.800 90.000 ;
        RECT 531.600 89.400 536.400 90.000 ;
        RECT 601.800 89.400 606.000 91.200 ;
        RECT 607.800 90.600 612.000 93.000 ;
        RECT 614.400 92.400 619.200 93.000 ;
        RECT 200.400 88.800 204.000 89.400 ;
        RECT 201.000 88.200 204.000 88.800 ;
        RECT 228.600 88.200 231.600 89.400 ;
        RECT 243.000 88.800 246.600 89.400 ;
        RECT 243.000 88.200 247.800 88.800 ;
        RECT 201.000 87.600 204.600 88.200 ;
        RECT 201.600 87.000 204.600 87.600 ;
        RECT 228.000 87.600 231.600 88.200 ;
        RECT 243.600 87.600 248.400 88.200 ;
        RECT 228.000 87.000 231.000 87.600 ;
        RECT 244.800 87.000 249.000 87.600 ;
        RECT 201.600 86.400 205.200 87.000 ;
        RECT 227.400 86.400 231.000 87.000 ;
        RECT 245.400 86.400 249.600 87.000 ;
        RECT 251.400 86.400 254.400 89.400 ;
        RECT 276.000 88.800 282.000 89.400 ;
        RECT 531.000 88.800 535.800 89.400 ;
        RECT 601.200 88.800 606.000 89.400 ;
        RECT 608.400 90.000 612.000 90.600 ;
        RECT 608.400 89.400 612.600 90.000 ;
        RECT 615.000 89.400 619.200 92.400 ;
        RECT 608.400 88.800 613.200 89.400 ;
        RECT 614.400 88.800 619.200 89.400 ;
        RECT 277.200 88.200 283.200 88.800 ;
        RECT 530.400 88.200 535.200 88.800 ;
        RECT 567.000 88.200 572.400 88.800 ;
        RECT 598.800 88.200 599.400 88.800 ;
        RECT 601.200 88.200 605.400 88.800 ;
        RECT 608.400 88.200 619.200 88.800 ;
        RECT 278.400 87.600 284.400 88.200 ;
        RECT 529.800 87.600 534.000 88.200 ;
        RECT 565.800 87.600 573.600 88.200 ;
        RECT 597.600 87.600 605.400 88.200 ;
        RECT 609.000 87.600 619.200 88.200 ;
        RECT 279.000 87.000 285.000 87.600 ;
        RECT 529.200 87.000 533.400 87.600 ;
        RECT 564.600 87.000 574.800 87.600 ;
        RECT 280.200 86.400 286.200 87.000 ;
        RECT 528.000 86.400 532.800 87.000 ;
        RECT 564.000 86.400 575.400 87.000 ;
        RECT 202.200 85.200 205.800 86.400 ;
        RECT 227.400 85.200 230.400 86.400 ;
        RECT 246.000 85.800 250.200 86.400 ;
        RECT 251.400 85.800 253.800 86.400 ;
        RECT 281.400 85.800 287.400 86.400 ;
        RECT 527.400 85.800 532.200 86.400 ;
        RECT 563.400 85.800 575.400 86.400 ;
        RECT 597.000 85.800 604.800 87.600 ;
        RECT 609.000 87.000 618.600 87.600 ;
        RECT 609.600 86.400 618.000 87.000 ;
        RECT 610.200 85.800 617.400 86.400 ;
        RECT 246.600 85.200 253.800 85.800 ;
        RECT 282.600 85.200 288.600 85.800 ;
        RECT 526.800 85.200 531.600 85.800 ;
        RECT 562.800 85.200 576.000 85.800 ;
        RECT 597.600 85.200 606.600 85.800 ;
        RECT 610.800 85.200 616.800 85.800 ;
        RECT 202.800 84.000 206.400 85.200 ;
        RECT 226.800 84.000 229.800 85.200 ;
        RECT 247.200 84.600 253.800 85.200 ;
        RECT 283.800 84.600 289.800 85.200 ;
        RECT 526.200 84.600 531.000 85.200 ;
        RECT 562.200 84.600 576.600 85.200 ;
        RECT 598.200 84.600 607.800 85.200 ;
        RECT 612.000 84.600 616.200 85.200 ;
        RECT 248.400 84.000 253.800 84.600 ;
        RECT 284.400 84.000 291.000 84.600 ;
        RECT 525.000 84.000 529.800 84.600 ;
        RECT 561.600 84.000 567.600 84.600 ;
        RECT 571.800 84.000 576.600 84.600 ;
        RECT 598.800 84.000 609.000 84.600 ;
        RECT 203.400 82.800 207.000 84.000 ;
        RECT 226.200 83.400 229.800 84.000 ;
        RECT 249.000 83.400 253.800 84.000 ;
        RECT 285.600 83.400 292.200 84.000 ;
        RECT 524.400 83.400 529.200 84.000 ;
        RECT 561.600 83.400 566.400 84.000 ;
        RECT 572.400 83.400 577.200 84.000 ;
        RECT 598.800 83.400 610.200 84.000 ;
        RECT 226.200 82.800 229.200 83.400 ;
        RECT 250.800 82.800 253.800 83.400 ;
        RECT 286.800 82.800 293.400 83.400 ;
        RECT 523.800 82.800 528.600 83.400 ;
        RECT 550.800 82.800 555.600 83.400 ;
        RECT 204.000 82.200 207.600 82.800 ;
        RECT 204.600 81.600 207.600 82.200 ;
        RECT 225.600 82.200 229.200 82.800 ;
        RECT 251.400 82.200 253.200 82.800 ;
        RECT 288.000 82.200 294.600 82.800 ;
        RECT 522.600 82.200 528.000 82.800 ;
        RECT 548.400 82.200 558.000 82.800 ;
        RECT 561.000 82.200 565.800 83.400 ;
        RECT 573.000 82.200 577.800 83.400 ;
        RECT 598.800 82.800 611.400 83.400 ;
        RECT 598.800 82.200 613.200 82.800 ;
        RECT 225.600 81.600 228.600 82.200 ;
        RECT 289.200 81.600 295.800 82.200 ;
        RECT 522.000 81.600 526.800 82.200 ;
        RECT 547.800 81.600 558.600 82.200 ;
        RECT 560.400 81.600 565.200 82.200 ;
        RECT 204.600 81.000 208.200 81.600 ;
        RECT 225.000 81.000 228.600 81.600 ;
        RECT 290.400 81.000 297.000 81.600 ;
        RECT 521.400 81.000 526.200 81.600 ;
        RECT 546.600 81.000 564.600 81.600 ;
        RECT 205.200 80.400 208.800 81.000 ;
        RECT 225.000 80.400 228.000 81.000 ;
        RECT 291.600 80.400 298.200 81.000 ;
        RECT 520.200 80.400 525.600 81.000 ;
        RECT 205.800 79.800 208.800 80.400 ;
        RECT 224.400 79.800 228.000 80.400 ;
        RECT 292.800 79.800 299.400 80.400 ;
        RECT 519.600 79.800 524.400 80.400 ;
        RECT 546.000 79.800 564.600 81.000 ;
        RECT 205.800 79.200 209.400 79.800 ;
        RECT 224.400 79.200 227.400 79.800 ;
        RECT 294.000 79.200 300.600 79.800 ;
        RECT 518.400 79.200 523.800 79.800 ;
        RECT 545.400 79.200 552.600 79.800 ;
        RECT 554.400 79.200 564.600 79.800 ;
        RECT 206.400 78.600 209.400 79.200 ;
        RECT 223.800 78.600 227.400 79.200 ;
        RECT 295.200 78.600 301.800 79.200 ;
        RECT 517.800 78.600 522.600 79.200 ;
        RECT 544.800 78.600 550.800 79.200 ;
        RECT 555.600 78.600 564.600 79.200 ;
        RECT 206.400 78.000 210.000 78.600 ;
        RECT 223.800 78.000 226.800 78.600 ;
        RECT 296.400 78.000 303.600 78.600 ;
        RECT 516.600 78.000 522.000 78.600 ;
        RECT 544.200 78.000 549.600 78.600 ;
        RECT 556.800 78.000 564.600 78.600 ;
        RECT 207.000 77.400 210.600 78.000 ;
        RECT 223.200 77.400 226.800 78.000 ;
        RECT 297.600 77.400 304.800 78.000 ;
        RECT 516.000 77.400 521.400 78.000 ;
        RECT 544.200 77.400 549.000 78.000 ;
        RECT 558.000 77.400 564.600 78.000 ;
        RECT 207.600 76.200 211.200 77.400 ;
        RECT 223.200 76.800 226.200 77.400 ;
        RECT 298.800 76.800 306.000 77.400 ;
        RECT 514.800 76.800 520.200 77.400 ;
        RECT 543.600 76.800 548.400 77.400 ;
        RECT 558.600 76.800 564.600 77.400 ;
        RECT 573.600 76.800 577.800 82.200 ;
        RECT 598.200 81.600 603.000 82.200 ;
        RECT 604.200 81.600 613.800 82.200 ;
        RECT 598.200 81.000 602.400 81.600 ;
        RECT 605.400 81.000 614.400 81.600 ;
        RECT 598.800 80.400 601.800 81.000 ;
        RECT 607.200 80.400 614.400 81.000 ;
        RECT 599.400 79.800 601.200 80.400 ;
        RECT 608.400 79.800 614.400 80.400 ;
        RECT 609.600 79.200 614.400 79.800 ;
        RECT 603.000 78.600 606.000 79.200 ;
        RECT 610.800 78.600 613.800 79.200 ;
        RECT 602.400 78.000 607.200 78.600 ;
        RECT 592.800 77.400 594.600 78.000 ;
        RECT 601.800 77.400 607.800 78.000 ;
        RECT 592.200 76.800 595.200 77.400 ;
        RECT 601.200 76.800 607.800 77.400 ;
        RECT 222.600 76.200 226.200 76.800 ;
        RECT 300.000 76.200 307.200 76.800 ;
        RECT 514.200 76.200 519.600 76.800 ;
        RECT 543.600 76.200 547.800 76.800 ;
        RECT 208.200 75.600 211.800 76.200 ;
        RECT 222.000 75.600 225.600 76.200 ;
        RECT 301.800 75.600 309.000 76.200 ;
        RECT 513.000 75.600 518.400 76.200 ;
        RECT 208.800 75.000 212.400 75.600 ;
        RECT 209.400 74.400 213.000 75.000 ;
        RECT 221.400 74.400 225.000 75.600 ;
        RECT 303.000 75.000 310.200 75.600 ;
        RECT 511.800 75.000 517.800 75.600 ;
        RECT 543.000 75.000 547.800 76.200 ;
        RECT 559.200 75.600 564.600 76.800 ;
        RECT 573.000 76.200 579.000 76.800 ;
        RECT 591.600 76.200 595.200 76.800 ;
        RECT 573.000 75.600 581.400 76.200 ;
        RECT 559.800 75.000 564.600 75.600 ;
        RECT 572.400 75.000 583.200 75.600 ;
        RECT 304.200 74.400 311.400 75.000 ;
        RECT 511.200 74.400 516.600 75.000 ;
        RECT 209.400 73.800 213.600 74.400 ;
        RECT 220.800 73.800 224.400 74.400 ;
        RECT 305.400 73.800 313.200 74.400 ;
        RECT 510.000 73.800 515.400 74.400 ;
        RECT 543.000 73.800 547.200 75.000 ;
        RECT 559.800 73.800 565.200 75.000 ;
        RECT 572.400 74.400 583.800 75.000 ;
        RECT 571.800 73.800 585.000 74.400 ;
        RECT 210.000 73.200 214.200 73.800 ;
        RECT 220.200 73.200 223.800 73.800 ;
        RECT 307.200 73.200 314.400 73.800 ;
        RECT 508.800 73.200 514.800 73.800 ;
        RECT 210.600 72.600 215.400 73.200 ;
        RECT 219.600 72.600 223.800 73.200 ;
        RECT 308.400 72.600 316.200 73.200 ;
        RECT 507.600 72.600 513.600 73.200 ;
        RECT 211.200 72.000 216.000 72.600 ;
        RECT 219.000 72.000 223.200 72.600 ;
        RECT 309.600 72.000 317.400 72.600 ;
        RECT 507.000 72.000 512.400 72.600 ;
        RECT 211.800 71.400 216.600 72.000 ;
        RECT 218.400 71.400 222.600 72.000 ;
        RECT 311.400 71.400 319.200 72.000 ;
        RECT 505.800 71.400 511.800 72.000 ;
        RECT 212.400 70.800 222.000 71.400 ;
        RECT 312.600 70.800 320.400 71.400 ;
        RECT 504.600 70.800 510.600 71.400 ;
        RECT 213.000 70.200 221.400 70.800 ;
        RECT 314.400 70.200 322.200 70.800 ;
        RECT 503.400 70.200 509.400 70.800 ;
        RECT 213.600 69.600 220.800 70.200 ;
        RECT 315.600 69.600 324.000 70.200 ;
        RECT 502.200 69.600 508.200 70.200 ;
        RECT 542.400 69.600 546.600 73.800 ;
        RECT 560.400 72.000 565.200 73.800 ;
        RECT 571.200 73.200 585.000 73.800 ;
        RECT 571.200 72.600 585.600 73.200 ;
        RECT 570.600 72.000 577.200 72.600 ;
        RECT 579.000 72.000 586.200 72.600 ;
        RECT 591.000 72.000 595.200 76.200 ;
        RECT 600.600 76.200 607.800 76.800 ;
        RECT 600.600 75.600 608.400 76.200 ;
        RECT 600.000 75.000 608.400 75.600 ;
        RECT 599.400 74.400 608.400 75.000 ;
        RECT 598.800 73.800 608.400 74.400 ;
        RECT 598.200 73.200 608.400 73.800 ;
        RECT 597.600 72.600 603.000 73.200 ;
        RECT 597.000 72.000 602.400 72.600 ;
        RECT 561.000 70.200 564.600 72.000 ;
        RECT 570.000 71.400 576.600 72.000 ;
        RECT 580.800 71.400 586.800 72.000 ;
        RECT 569.400 70.800 575.400 71.400 ;
        RECT 569.400 70.200 574.800 70.800 ;
        RECT 582.000 70.200 586.800 71.400 ;
        RECT 591.000 71.400 602.400 72.000 ;
        RECT 591.000 70.800 601.800 71.400 ;
        RECT 591.600 70.200 601.200 70.800 ;
        RECT 604.200 70.200 608.400 73.200 ;
        RECT 561.600 69.600 564.000 70.200 ;
        RECT 569.400 69.600 574.200 70.200 ;
        RECT 582.600 69.600 587.400 70.200 ;
        RECT 591.600 69.600 600.600 70.200 ;
        RECT 214.200 69.000 219.600 69.600 ;
        RECT 317.400 69.000 325.800 69.600 ;
        RECT 501.000 69.000 507.000 69.600 ;
        RECT 214.800 68.400 219.000 69.000 ;
        RECT 318.600 68.400 327.000 69.000 ;
        RECT 499.200 68.400 506.400 69.000 ;
        RECT 543.000 68.400 547.200 69.600 ;
        RECT 561.600 69.000 563.400 69.600 ;
        RECT 569.400 69.000 573.600 69.600 ;
        RECT 570.600 68.400 571.800 69.000 ;
        RECT 216.000 67.800 218.400 68.400 ;
        RECT 320.400 67.800 328.800 68.400 ;
        RECT 498.000 67.800 505.200 68.400 ;
        RECT 322.200 67.200 330.600 67.800 ;
        RECT 496.800 67.200 504.000 67.800 ;
        RECT 543.000 67.200 547.800 68.400 ;
        RECT 323.400 66.600 332.400 67.200 ;
        RECT 495.600 66.600 502.800 67.200 ;
        RECT 543.600 66.600 547.800 67.200 ;
        RECT 565.200 66.600 568.800 67.200 ;
        RECT 325.200 66.000 334.200 66.600 ;
        RECT 493.800 66.000 501.000 66.600 ;
        RECT 543.600 66.000 548.400 66.600 ;
        RECT 564.600 66.000 569.400 66.600 ;
        RECT 327.000 65.400 336.600 66.000 ;
        RECT 492.600 65.400 499.800 66.000 ;
        RECT 544.200 65.400 549.000 66.000 ;
        RECT 564.000 65.400 569.400 66.000 ;
        RECT 583.200 65.400 587.400 69.600 ;
        RECT 592.200 69.000 599.400 69.600 ;
        RECT 603.600 69.000 607.800 70.200 ;
        RECT 592.800 68.400 598.800 69.000 ;
        RECT 603.000 68.400 607.800 69.000 ;
        RECT 593.400 67.800 597.600 68.400 ;
        RECT 603.000 67.800 607.200 68.400 ;
        RECT 602.400 67.200 607.200 67.800 ;
        RECT 601.800 66.600 607.200 67.200 ;
        RECT 601.200 66.000 606.600 66.600 ;
        RECT 600.600 65.400 606.000 66.000 ;
        RECT 612.000 65.400 613.200 66.000 ;
        RECT 328.800 64.800 338.400 65.400 ;
        RECT 490.800 64.800 498.600 65.400 ;
        RECT 544.800 64.800 549.600 65.400 ;
        RECT 564.000 64.800 570.000 65.400 ;
        RECT 582.600 64.800 586.800 65.400 ;
        RECT 600.000 64.800 605.400 65.400 ;
        RECT 330.600 64.200 340.200 64.800 ;
        RECT 489.000 64.200 497.400 64.800 ;
        RECT 544.800 64.200 550.800 64.800 ;
        RECT 332.400 63.600 342.600 64.200 ;
        RECT 487.200 63.600 495.600 64.200 ;
        RECT 545.400 63.600 551.400 64.200 ;
        RECT 334.200 63.000 344.400 63.600 ;
        RECT 485.400 63.000 494.400 63.600 ;
        RECT 546.000 63.000 560.400 63.600 ;
        RECT 563.400 63.000 570.000 64.800 ;
        RECT 582.000 63.600 586.800 64.800 ;
        RECT 600.600 64.200 604.800 64.800 ;
        RECT 611.400 64.200 613.200 65.400 ;
        RECT 600.600 63.600 604.200 64.200 ;
        RECT 610.800 63.600 613.200 64.200 ;
        RECT 573.000 63.000 576.000 63.600 ;
        RECT 580.800 63.000 586.200 63.600 ;
        RECT 610.200 63.000 613.200 63.600 ;
        RECT 336.000 62.400 346.800 63.000 ;
        RECT 483.600 62.400 492.600 63.000 ;
        RECT 546.600 62.400 561.000 63.000 ;
        RECT 338.400 61.800 349.200 62.400 ;
        RECT 481.800 61.800 491.400 62.400 ;
        RECT 547.200 61.800 561.000 62.400 ;
        RECT 340.200 61.200 351.600 61.800 ;
        RECT 479.400 61.200 491.400 61.800 ;
        RECT 547.800 61.200 561.000 61.800 ;
        RECT 564.000 62.400 570.000 63.000 ;
        RECT 572.400 62.400 586.200 63.000 ;
        RECT 609.600 62.400 613.200 63.000 ;
        RECT 564.000 61.200 569.400 62.400 ;
        RECT 572.400 61.800 585.600 62.400 ;
        RECT 609.000 61.800 612.600 62.400 ;
        RECT 572.400 61.200 585.000 61.800 ;
        RECT 608.400 61.200 612.000 61.800 ;
        RECT 342.000 60.600 354.000 61.200 ;
        RECT 477.600 60.600 491.400 61.200 ;
        RECT 548.400 60.600 561.000 61.200 ;
        RECT 565.200 60.600 568.800 61.200 ;
        RECT 572.400 60.600 584.400 61.200 ;
        RECT 607.800 60.600 612.000 61.200 ;
        RECT 344.400 60.000 356.400 60.600 ;
        RECT 474.600 60.000 493.200 60.600 ;
        RECT 549.600 60.000 559.800 60.600 ;
        RECT 573.000 60.000 584.400 60.600 ;
        RECT 607.200 60.000 612.000 60.600 ;
        RECT 346.800 59.400 359.400 60.000 ;
        RECT 472.200 59.400 484.200 60.000 ;
        RECT 487.200 59.400 495.600 60.000 ;
        RECT 550.800 59.400 559.200 60.000 ;
        RECT 573.600 59.400 584.400 60.000 ;
        RECT 606.000 59.400 611.400 60.000 ;
        RECT 349.200 58.800 362.400 59.400 ;
        RECT 469.200 58.800 481.800 59.400 ;
        RECT 488.400 58.800 499.800 59.400 ;
        RECT 552.600 58.800 558.600 59.400 ;
        RECT 574.800 58.800 585.600 59.400 ;
        RECT 605.400 58.800 610.800 59.400 ;
        RECT 351.600 58.200 365.400 58.800 ;
        RECT 465.600 58.200 480.000 58.800 ;
        RECT 489.600 58.200 505.800 58.800 ;
        RECT 552.600 58.200 558.000 58.800 ;
        RECT 576.000 58.200 586.800 58.800 ;
        RECT 604.800 58.200 610.800 58.800 ;
        RECT 354.000 57.600 368.400 58.200 ;
        RECT 462.600 57.600 477.600 58.200 ;
        RECT 490.800 57.600 517.800 58.200 ;
        RECT 356.400 57.000 372.000 57.600 ;
        RECT 458.400 57.000 475.200 57.600 ;
        RECT 493.200 57.000 525.000 57.600 ;
        RECT 552.600 57.000 557.400 58.200 ;
        RECT 576.600 57.600 588.000 58.200 ;
        RECT 603.600 57.600 610.200 58.200 ;
        RECT 577.200 57.000 589.800 57.600 ;
        RECT 602.400 57.000 609.600 57.600 ;
        RECT 359.400 56.400 376.200 57.000 ;
        RECT 454.800 56.400 472.200 57.000 ;
        RECT 495.600 56.400 528.600 57.000 ;
        RECT 552.000 56.400 556.800 57.000 ;
        RECT 577.800 56.400 591.600 57.000 ;
        RECT 601.800 56.400 609.000 57.000 ;
        RECT 362.400 55.800 380.400 56.400 ;
        RECT 450.000 55.800 469.200 56.400 ;
        RECT 500.400 55.800 531.000 56.400 ;
        RECT 552.000 55.800 556.200 56.400 ;
        RECT 365.400 55.200 385.200 55.800 ;
        RECT 444.600 55.200 465.600 55.800 ;
        RECT 506.400 55.200 532.800 55.800 ;
        RECT 551.400 55.200 556.200 55.800 ;
        RECT 566.400 55.200 569.400 56.400 ;
        RECT 578.400 55.800 608.400 56.400 ;
        RECT 579.000 55.200 607.200 55.800 ;
        RECT 368.400 54.600 391.200 55.200 ;
        RECT 438.000 54.600 462.000 55.200 ;
        RECT 519.600 54.600 534.000 55.200 ;
        RECT 372.000 54.000 399.600 54.600 ;
        RECT 430.200 54.000 458.400 54.600 ;
        RECT 525.600 54.000 534.600 54.600 ;
        RECT 551.400 54.000 555.600 55.200 ;
        RECT 376.200 53.400 454.200 54.000 ;
        RECT 528.600 53.400 535.200 54.000 ;
        RECT 380.400 52.800 449.400 53.400 ;
        RECT 530.400 52.800 535.200 53.400 ;
        RECT 550.800 53.400 555.600 54.000 ;
        RECT 565.800 53.400 570.000 55.200 ;
        RECT 385.800 52.200 444.600 52.800 ;
        RECT 532.200 52.200 535.800 52.800 ;
        RECT 391.800 51.600 441.600 52.200 ;
        RECT 533.400 51.600 535.800 52.200 ;
        RECT 400.800 51.000 441.600 51.600 ;
        RECT 534.000 51.000 537.000 51.600 ;
        RECT 411.600 49.800 415.200 51.000 ;
        RECT 425.400 50.400 442.200 51.000 ;
        RECT 534.600 50.400 537.600 51.000 ;
        RECT 426.000 49.800 436.200 50.400 ;
        RECT 412.200 48.600 415.800 49.800 ;
        RECT 427.800 49.200 436.200 49.800 ;
        RECT 439.200 49.800 442.800 50.400 ;
        RECT 535.200 49.800 538.200 50.400 ;
        RECT 439.200 49.200 443.400 49.800 ;
        RECT 535.800 49.200 538.800 49.800 ;
        RECT 430.200 48.600 436.800 49.200 ;
        RECT 439.800 48.600 443.400 49.200 ;
        RECT 518.400 48.600 525.000 49.200 ;
        RECT 536.400 48.600 539.400 49.200 ;
        RECT 550.800 48.600 555.000 53.400 ;
        RECT 565.200 51.000 570.000 53.400 ;
        RECT 579.000 51.000 583.200 55.200 ;
        RECT 585.000 54.600 606.600 55.200 ;
        RECT 586.200 54.000 605.400 54.600 ;
        RECT 587.400 53.400 604.800 54.000 ;
        RECT 589.800 52.800 603.600 53.400 ;
        RECT 591.600 52.200 601.200 52.800 ;
        RECT 596.400 51.600 597.600 52.200 ;
        RECT 564.600 49.800 570.600 51.000 ;
        RECT 578.400 50.400 583.200 51.000 ;
        RECT 578.400 49.800 582.600 50.400 ;
        RECT 564.000 49.200 570.600 49.800 ;
        RECT 577.800 49.200 582.600 49.800 ;
        RECT 564.000 48.600 571.800 49.200 ;
        RECT 577.200 48.600 582.600 49.200 ;
        RECT 412.800 48.000 416.400 48.600 ;
        RECT 431.400 48.000 438.600 48.600 ;
        RECT 439.800 48.000 444.000 48.600 ;
        RECT 516.600 48.000 526.200 48.600 ;
        RECT 536.400 48.000 540.000 48.600 ;
        RECT 550.800 48.000 555.600 48.600 ;
        RECT 563.400 48.000 572.400 48.600 ;
        RECT 577.200 48.000 582.000 48.600 ;
        RECT 413.400 46.800 417.000 48.000 ;
        RECT 432.000 47.400 445.200 48.000 ;
        RECT 515.400 47.400 527.400 48.000 ;
        RECT 537.000 47.400 540.000 48.000 ;
        RECT 551.400 47.400 556.200 48.000 ;
        RECT 562.200 47.400 581.400 48.000 ;
        RECT 433.200 46.800 445.800 47.400 ;
        RECT 514.200 46.800 528.600 47.400 ;
        RECT 537.000 46.800 540.600 47.400 ;
        RECT 551.400 46.800 556.800 47.400 ;
        RECT 561.600 46.800 581.400 47.400 ;
        RECT 414.000 46.200 417.600 46.800 ;
        RECT 434.400 46.200 445.800 46.800 ;
        RECT 513.600 46.200 529.200 46.800 ;
        RECT 414.600 45.600 418.200 46.200 ;
        RECT 436.200 45.600 445.200 46.200 ;
        RECT 513.000 45.600 518.400 46.200 ;
        RECT 524.400 45.600 529.800 46.200 ;
        RECT 415.200 45.000 418.800 45.600 ;
        RECT 438.600 45.000 444.600 45.600 ;
        RECT 513.000 45.000 517.200 45.600 ;
        RECT 526.200 45.000 530.400 45.600 ;
        RECT 537.600 45.000 540.600 46.800 ;
        RECT 552.000 46.200 567.000 46.800 ;
        RECT 568.200 46.200 580.800 46.800 ;
        RECT 552.000 45.600 566.400 46.200 ;
        RECT 568.800 45.600 580.200 46.200 ;
        RECT 552.600 45.000 565.800 45.600 ;
        RECT 569.400 45.000 579.600 45.600 ;
        RECT 415.200 44.400 419.400 45.000 ;
        RECT 513.000 44.400 516.000 45.000 ;
        RECT 526.800 44.400 531.000 45.000 ;
        RECT 537.600 44.400 541.200 45.000 ;
        RECT 553.200 44.400 565.200 45.000 ;
        RECT 570.000 44.400 579.000 45.000 ;
        RECT 415.800 43.800 419.400 44.400 ;
        RECT 498.000 43.800 499.200 44.400 ;
        RECT 513.000 43.800 515.400 44.400 ;
        RECT 527.400 43.800 531.600 44.400 ;
        RECT 536.400 43.800 541.800 44.400 ;
        RECT 553.800 43.800 564.600 44.400 ;
        RECT 571.800 43.800 577.200 44.400 ;
        RECT 416.400 43.200 420.000 43.800 ;
        RECT 493.200 43.200 502.800 43.800 ;
        RECT 513.000 43.200 514.800 43.800 ;
        RECT 528.000 43.200 531.600 43.800 ;
        RECT 535.800 43.200 543.000 43.800 ;
        RECT 555.000 43.200 564.000 43.800 ;
        RECT 417.000 42.600 420.600 43.200 ;
        RECT 490.800 42.600 504.600 43.200 ;
        RECT 528.600 42.600 532.200 43.200 ;
        RECT 535.200 42.600 543.600 43.200 ;
        RECT 556.200 42.600 562.800 43.200 ;
        RECT 417.600 42.000 421.200 42.600 ;
        RECT 489.000 42.000 505.800 42.600 ;
        RECT 529.200 42.000 532.200 42.600 ;
        RECT 534.600 42.000 543.600 42.600 ;
        RECT 559.200 42.000 560.400 42.600 ;
        RECT 417.600 41.400 421.800 42.000 ;
        RECT 487.200 41.400 507.000 42.000 ;
        RECT 529.200 41.400 532.800 42.000 ;
        RECT 418.200 40.800 422.400 41.400 ;
        RECT 486.600 40.800 496.800 41.400 ;
        RECT 500.400 40.800 507.600 41.400 ;
        RECT 418.800 40.200 423.000 40.800 ;
        RECT 486.000 40.200 493.200 40.800 ;
        RECT 502.800 40.200 508.800 40.800 ;
        RECT 529.800 40.200 532.800 41.400 ;
        RECT 534.600 41.400 538.200 42.000 ;
        RECT 540.600 41.400 544.200 42.000 ;
        RECT 534.600 40.800 537.600 41.400 ;
        RECT 541.200 40.800 544.200 41.400 ;
        RECT 419.400 39.600 424.200 40.200 ;
        RECT 486.600 39.600 490.800 40.200 ;
        RECT 504.000 39.600 509.400 40.200 ;
        RECT 420.000 39.000 424.800 39.600 ;
        RECT 487.200 39.000 488.400 39.600 ;
        RECT 505.200 39.000 510.000 39.600 ;
        RECT 420.600 38.400 425.400 39.000 ;
        RECT 506.400 38.400 510.600 39.000 ;
        RECT 421.800 37.800 426.000 38.400 ;
        RECT 507.000 37.800 510.600 38.400 ;
        RECT 530.400 37.800 533.400 40.200 ;
        RECT 534.600 37.800 537.000 40.800 ;
        RECT 541.200 40.200 544.800 40.800 ;
        RECT 422.400 37.200 427.200 37.800 ;
        RECT 507.600 37.200 511.200 37.800 ;
        RECT 531.000 37.200 537.000 37.800 ;
        RECT 423.000 36.600 427.800 37.200 ;
        RECT 423.600 36.000 429.000 36.600 ;
        RECT 508.200 36.000 511.800 37.200 ;
        RECT 522.600 36.000 525.600 36.600 ;
        RECT 424.200 35.400 429.600 36.000 ;
        RECT 508.800 35.400 511.800 36.000 ;
        RECT 522.000 35.400 526.200 36.000 ;
        RECT 425.400 34.800 430.800 35.400 ;
        RECT 426.000 34.200 432.000 34.800 ;
        RECT 427.200 33.600 433.800 34.200 ;
        RECT 427.800 33.000 435.600 33.600 ;
        RECT 509.400 33.000 512.400 35.400 ;
        RECT 521.400 34.200 526.800 35.400 ;
        RECT 521.400 33.600 527.400 34.200 ;
        RECT 520.800 33.000 527.400 33.600 ;
        RECT 429.000 32.400 437.400 33.000 ;
        RECT 430.200 31.800 439.800 32.400 ;
        RECT 504.000 31.800 506.400 32.400 ;
        RECT 432.000 31.200 442.200 31.800 ;
        RECT 502.800 31.200 507.600 31.800 ;
        RECT 433.800 30.600 444.600 31.200 ;
        RECT 502.200 30.600 508.200 31.200 ;
        RECT 435.600 30.000 447.600 30.600 ;
        RECT 502.200 30.000 508.800 30.600 ;
        RECT 437.400 29.400 451.200 30.000 ;
        RECT 501.600 29.400 508.800 30.000 ;
        RECT 510.000 29.400 513.000 33.000 ;
        RECT 520.800 32.400 528.000 33.000 ;
        RECT 520.800 30.600 523.800 32.400 ;
        RECT 525.000 30.600 528.000 32.400 ;
        RECT 531.000 31.800 537.600 37.200 ;
        RECT 541.800 34.800 544.800 40.200 ;
        RECT 541.200 33.000 544.200 34.800 ;
        RECT 531.000 31.200 533.400 31.800 ;
        RECT 520.800 30.000 523.200 30.600 ;
        RECT 439.800 28.800 453.600 29.400 ;
        RECT 501.000 28.800 504.600 29.400 ;
        RECT 505.800 28.800 513.000 29.400 ;
        RECT 442.200 28.200 456.000 28.800 ;
        RECT 444.600 27.600 457.800 28.200 ;
        RECT 447.600 27.000 459.600 27.600 ;
        RECT 501.000 27.000 504.000 28.800 ;
        RECT 506.400 27.600 512.400 28.800 ;
        RECT 450.000 26.400 461.400 27.000 ;
        RECT 453.000 25.800 462.600 26.400 ;
        RECT 456.000 25.200 464.400 25.800 ;
        RECT 457.800 24.600 465.600 25.200 ;
        RECT 459.600 24.000 466.800 24.600 ;
        RECT 460.800 23.400 468.600 24.000 ;
        RECT 462.600 22.800 469.800 23.400 ;
        RECT 463.800 22.200 471.000 22.800 ;
        RECT 465.000 21.600 472.200 22.200 ;
        RECT 466.800 21.000 473.400 21.600 ;
        RECT 500.400 21.000 503.400 27.000 ;
        RECT 507.000 25.800 512.400 27.600 ;
        RECT 507.600 23.400 511.800 25.800 ;
        RECT 520.200 23.400 523.200 30.000 ;
        RECT 525.600 30.000 528.000 30.600 ;
        RECT 525.600 25.200 528.600 30.000 ;
        RECT 530.400 27.600 533.400 31.200 ;
        RECT 534.600 28.200 537.600 31.800 ;
        RECT 540.600 32.400 544.200 33.000 ;
        RECT 540.600 31.200 543.600 32.400 ;
        RECT 540.000 30.000 543.000 31.200 ;
        RECT 539.400 29.400 543.000 30.000 ;
        RECT 539.400 28.800 542.400 29.400 ;
        RECT 535.200 27.600 537.600 28.200 ;
        RECT 538.800 28.200 542.400 28.800 ;
        RECT 538.800 27.600 541.800 28.200 ;
        RECT 529.800 25.200 532.800 27.600 ;
        RECT 535.200 27.000 541.800 27.600 ;
        RECT 535.200 25.800 541.200 27.000 ;
        RECT 534.600 25.200 540.600 25.800 ;
        RECT 525.600 24.600 540.600 25.200 ;
        RECT 507.600 21.600 511.200 23.400 ;
        RECT 468.000 20.400 474.600 21.000 ;
        RECT 501.000 20.400 503.400 21.000 ;
        RECT 507.000 20.400 510.600 21.600 ;
        RECT 519.600 20.400 523.200 23.400 ;
        RECT 525.000 23.400 528.000 24.600 ;
        RECT 529.200 23.400 540.000 24.600 ;
        RECT 525.000 22.800 539.400 23.400 ;
        RECT 525.000 22.200 538.800 22.800 ;
        RECT 525.000 21.600 538.200 22.200 ;
        RECT 525.000 21.000 532.800 21.600 ;
        RECT 535.200 21.000 537.600 21.600 ;
        RECT 469.200 19.800 475.800 20.400 ;
        RECT 470.400 19.200 477.000 19.800 ;
        RECT 471.600 18.600 478.200 19.200 ;
        RECT 472.800 18.000 479.400 18.600 ;
        RECT 474.000 17.400 480.600 18.000 ;
        RECT 501.000 17.400 504.000 20.400 ;
        RECT 507.000 19.800 511.200 20.400 ;
        RECT 520.200 19.800 523.200 20.400 ;
        RECT 524.400 20.400 531.000 21.000 ;
        RECT 507.000 19.200 511.800 19.800 ;
        RECT 506.400 18.600 511.800 19.200 ;
        RECT 520.200 18.600 522.600 19.800 ;
        RECT 524.400 19.200 530.400 20.400 ;
        RECT 506.400 18.000 512.400 18.600 ;
        RECT 506.400 17.400 513.000 18.000 ;
        RECT 519.600 17.400 522.600 18.600 ;
        RECT 523.800 18.000 529.800 19.200 ;
        RECT 523.800 17.400 529.200 18.000 ;
        RECT 475.200 16.800 481.800 17.400 ;
        RECT 476.400 16.200 483.600 16.800 ;
        RECT 477.600 15.600 484.800 16.200 ;
        RECT 478.800 15.000 486.000 15.600 ;
        RECT 501.600 15.000 504.600 17.400 ;
        RECT 506.400 16.800 513.600 17.400 ;
        RECT 519.600 16.800 528.600 17.400 ;
        RECT 505.800 15.000 508.800 16.800 ;
        RECT 510.000 16.200 514.800 16.800 ;
        RECT 519.600 16.200 528.000 16.800 ;
        RECT 510.600 15.600 528.000 16.200 ;
        RECT 511.200 15.000 527.400 15.600 ;
        RECT 480.600 14.400 487.200 15.000 ;
        RECT 481.800 13.800 489.000 14.400 ;
        RECT 501.600 13.800 508.200 15.000 ;
        RECT 511.800 14.400 526.200 15.000 ;
        RECT 513.000 13.800 525.600 14.400 ;
        RECT 483.000 13.200 490.800 13.800 ;
        RECT 500.400 13.200 508.200 13.800 ;
        RECT 514.200 13.200 525.000 13.800 ;
        RECT 484.200 12.600 507.600 13.200 ;
        RECT 485.400 12.000 507.600 12.600 ;
        RECT 519.000 12.000 524.400 13.200 ;
        RECT 487.200 11.400 507.600 12.000 ;
        RECT 518.400 11.400 523.800 12.000 ;
        RECT 488.400 10.800 507.000 11.400 ;
        RECT 490.800 10.200 500.400 10.800 ;
        RECT 502.200 10.200 507.000 10.800 ;
        RECT 518.400 10.200 523.200 11.400 ;
        RECT 502.200 8.400 506.400 10.200 ;
        RECT 517.800 9.600 522.600 10.200 ;
        RECT 517.800 9.000 521.400 9.600 ;
        RECT 518.400 8.400 520.800 9.000 ;
        RECT 502.200 7.200 505.800 8.400 ;
        RECT 501.600 6.600 505.200 7.200 ;
        RECT 501.600 6.000 504.600 6.600 ;
        RECT 502.200 5.400 504.600 6.000 ;
        RECT 502.200 4.800 504.000 5.400 ;
  END
END tholin
END LIBRARY

